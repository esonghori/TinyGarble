
module aes_comb ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [1279:0] key;
  output [127:0] out;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683;

  XNOR U1 ( .A(n29497), .B(n29488), .Z(n29495) );
  XNOR U2 ( .A(n28559), .B(n28550), .Z(n28557) );
  XNOR U3 ( .A(n29396), .B(n29386), .Z(n29393) );
  XOR U4 ( .A(n27465), .B(n27472), .Z(n27471) );
  XNOR U5 ( .A(n27353), .B(n27344), .Z(n27351) );
  XOR U6 ( .A(n28915), .B(n28922), .Z(n28921) );
  XOR U7 ( .A(n17269), .B(n15172), .Z(n17268) );
  XOR U8 ( .A(key[840]), .B(n10987), .Z(n10992) );
  XNOR U9 ( .A(n28158), .B(n28148), .Z(n28155) );
  XNOR U10 ( .A(n28691), .B(n28682), .Z(n28689) );
  XNOR U11 ( .A(n27979), .B(n27969), .Z(n27976) );
  XNOR U12 ( .A(n27265), .B(n27256), .Z(n27263) );
  XNOR U13 ( .A(n29287), .B(n29278), .Z(n29285) );
  XNOR U14 ( .A(n27441), .B(n27431), .Z(n27438) );
  XNOR U15 ( .A(n27177), .B(n27167), .Z(n27175) );
  XNOR U16 ( .A(n28506), .B(n28516), .Z(n28521) );
  XOR U17 ( .A(n29420), .B(n29427), .Z(n29426) );
  NOR U18 ( .A(n29498), .B(n29497), .Z(n29494) );
  NOR U19 ( .A(n28872), .B(n28886), .Z(n28877) );
  XNOR U20 ( .A(n29589), .B(n29603), .Z(n29182) );
  XNOR U21 ( .A(n26960), .B(n27334), .Z(n26954) );
  XNOR U22 ( .A(n23309), .B(n21519), .Z(n21511) );
  XOR U23 ( .A(n22940), .B(n22931), .Z(n22742) );
  XNOR U24 ( .A(n21058), .B(n21108), .Z(n20972) );
  XNOR U25 ( .A(n18134), .B(n18124), .Z(n18131) );
  AND U26 ( .A(n19328), .B(n18991), .Z(n19319) );
  XOR U27 ( .A(n18057), .B(n18519), .Z(n17979) );
  XOR U28 ( .A(n17671), .B(n19573), .Z(n17604) );
  NANDN U29 ( .A(n19589), .B(n17674), .Z(n18661) );
  XNOR U30 ( .A(n11997), .B(n11993), .Z(n11981) );
  XNOR U31 ( .A(n9478), .B(n10358), .Z(n10363) );
  XOR U32 ( .A(n14630), .B(n14731), .Z(n14629) );
  ANDN U33 ( .B(n13424), .A(n13447), .Z(n12920) );
  XNOR U34 ( .A(n10968), .B(n9430), .Z(n11890) );
  NANDN U35 ( .A(n9646), .B(n8675), .Z(n8570) );
  XNOR U36 ( .A(n27871), .B(n27862), .Z(n27869) );
  XOR U37 ( .A(n28003), .B(n28010), .Z(n28009) );
  XOR U38 ( .A(n27959), .B(n27828), .Z(n27957) );
  XOR U39 ( .A(n29646), .B(n29653), .Z(n29652) );
  XOR U40 ( .A(n28184), .B(n28191), .Z(n28190) );
  XNOR U41 ( .A(n28371), .B(n28664), .Z(n28666) );
  XNOR U42 ( .A(n28891), .B(n28881), .Z(n28888) );
  XNOR U43 ( .A(n28791), .B(n28782), .Z(n28789) );
  NOR U44 ( .A(n29288), .B(n29287), .Z(n29284) );
  XNOR U45 ( .A(n29161), .B(n29478), .Z(n29214) );
  XNOR U46 ( .A(n27267), .B(n27254), .Z(n26971) );
  NOR U47 ( .A(n27354), .B(n27353), .Z(n27350) );
  XNOR U48 ( .A(n26972), .B(n27246), .Z(n26966) );
  XNOR U49 ( .A(n27179), .B(n27165), .Z(n27011) );
  XOR U50 ( .A(n29175), .B(n29377), .Z(n29174) );
  XNOR U51 ( .A(n28641), .B(n28636), .Z(n28474) );
  XNOR U52 ( .A(n28508), .B(n28533), .Z(n28409) );
  XNOR U53 ( .A(n29201), .B(n29170), .Z(n25550) );
  XOR U54 ( .A(n27107), .B(n27118), .Z(n27000) );
  XOR U55 ( .A(n24638), .B(n25114), .Z(n26297) );
  XOR U56 ( .A(n25925), .B(n25900), .Z(n25936) );
  XNOR U57 ( .A(n25380), .B(n26185), .Z(n26181) );
  ANDN U58 ( .B(n24898), .A(n25122), .Z(n24930) );
  XNOR U59 ( .A(n23885), .B(n24184), .Z(n24101) );
  ANDN U60 ( .B(n24876), .A(n25429), .Z(n24942) );
  XNOR U61 ( .A(n24612), .B(n24611), .Z(n24610) );
  XOR U62 ( .A(n24895), .B(n24913), .Z(n24826) );
  XNOR U63 ( .A(n23896), .B(n24383), .Z(n23918) );
  XOR U64 ( .A(n24052), .B(n24095), .Z(n23840) );
  XNOR U65 ( .A(n22472), .B(n22462), .Z(n22469) );
  XNOR U66 ( .A(n21684), .B(n25815), .Z(n25814) );
  XOR U67 ( .A(n21233), .B(n23032), .Z(n26559) );
  XNOR U68 ( .A(n21511), .B(n24764), .Z(n24755) );
  ANDN U69 ( .B(n21071), .A(n21114), .Z(n21060) );
  ANDN U70 ( .B(n21948), .A(n22116), .Z(n21886) );
  XOR U71 ( .A(n23707), .B(n23702), .Z(n23579) );
  XOR U72 ( .A(n22882), .B(n22888), .Z(n22767) );
  XOR U73 ( .A(n23167), .B(n23178), .Z(n22759) );
  XNOR U74 ( .A(n20892), .B(n20893), .Z(n18617) );
  XNOR U75 ( .A(n20347), .B(n20337), .Z(n20344) );
  XOR U76 ( .A(n22680), .B(n22793), .Z(n22838) );
  XNOR U77 ( .A(key[511]), .B(n18341), .Z(n18337) );
  XNOR U78 ( .A(n20810), .B(n20800), .Z(n20807) );
  XOR U79 ( .A(n18204), .B(n20277), .Z(n20273) );
  XNOR U80 ( .A(n20566), .B(n20780), .Z(n20775) );
  ANDN U81 ( .B(n17984), .A(n17983), .Z(n17981) );
  OR U82 ( .A(n20317), .B(n19892), .Z(n20316) );
  NOR U83 ( .A(n19760), .B(n19906), .Z(n19839) );
  XNOR U84 ( .A(n17937), .B(n17969), .Z(n17858) );
  ANDN U85 ( .B(n19807), .A(n20178), .Z(n19833) );
  XOR U86 ( .A(n21719), .B(n21710), .Z(n20657) );
  XNOR U87 ( .A(n16216), .B(n17263), .Z(n17853) );
  XOR U88 ( .A(n22602), .B(n22593), .Z(n20574) );
  XNOR U89 ( .A(n18791), .B(n18899), .Z(n18898) );
  XNOR U90 ( .A(n18928), .B(n19432), .Z(n18897) );
  XNOR U91 ( .A(n15599), .B(n16391), .Z(n17380) );
  XNOR U92 ( .A(n15463), .B(n15464), .Z(n15462) );
  XOR U93 ( .A(n17681), .B(n17693), .Z(n17598) );
  XOR U94 ( .A(n17715), .B(n17727), .Z(n17588) );
  XOR U95 ( .A(n16999), .B(n17019), .Z(n16722) );
  XNOR U96 ( .A(n12471), .B(n12487), .Z(n14126) );
  XNOR U97 ( .A(n17602), .B(n19562), .Z(n17649) );
  XNOR U98 ( .A(n12384), .B(n12374), .Z(n12381) );
  ANDN U99 ( .B(n12023), .A(n12502), .Z(n12317) );
  NANDN U100 ( .A(n17442), .B(n14643), .Z(n17413) );
  XNOR U101 ( .A(n12799), .B(n12858), .Z(n12760) );
  XNOR U102 ( .A(n12851), .B(n13132), .Z(n12952) );
  AND U103 ( .A(n14665), .B(n14666), .Z(n14662) );
  XOR U104 ( .A(n14617), .B(n14613), .Z(n14547) );
  XNOR U105 ( .A(n17411), .B(n17436), .Z(n14619) );
  XNOR U106 ( .A(n9976), .B(n9966), .Z(n9973) );
  XNOR U107 ( .A(n10881), .B(n10871), .Z(n10878) );
  XNOR U108 ( .A(n10489), .B(n11394), .Z(n9597) );
  XOR U109 ( .A(n12909), .B(n12932), .Z(n12786) );
  XNOR U110 ( .A(n10366), .B(n10948), .Z(n10991) );
  XNOR U111 ( .A(n11752), .B(n11742), .Z(n11749) );
  XNOR U112 ( .A(n11622), .B(n12676), .Z(n12668) );
  XNOR U113 ( .A(key[850]), .B(n9471), .Z(n10327) );
  AND U114 ( .A(n9971), .B(n9935), .Z(n9962) );
  XNOR U115 ( .A(n12871), .B(n12973), .Z(n10214) );
  XNOR U116 ( .A(n10746), .B(n11036), .Z(n11028) );
  XNOR U117 ( .A(n9003), .B(n9173), .Z(n8914) );
  XNOR U118 ( .A(n8677), .B(n9720), .Z(n8688) );
  XOR U119 ( .A(n5951), .B(n5956), .Z(n5970) );
  XNOR U120 ( .A(n3012), .B(n2992), .Z(n4963) );
  XOR U121 ( .A(n4112), .B(n4110), .Z(n4107) );
  XNOR U122 ( .A(n5144), .B(n5134), .Z(n5141) );
  XNOR U123 ( .A(n3603), .B(n3813), .Z(n3865) );
  XOR U124 ( .A(n2687), .B(n3945), .Z(n3941) );
  XNOR U125 ( .A(n4652), .B(n4664), .Z(n4728) );
  XOR U126 ( .A(n3524), .B(n3499), .Z(n3523) );
  XOR U127 ( .A(n542), .B(n533), .Z(n462) );
  XNOR U128 ( .A(n29593), .B(n29108), .Z(n29640) );
  XNOR U129 ( .A(n28074), .B(n28061), .Z(n28069) );
  XOR U130 ( .A(n27863), .B(n27877), .Z(n27874) );
  XOR U131 ( .A(n28683), .B(n28697), .Z(n28694) );
  XNOR U132 ( .A(n28671), .B(n28661), .Z(n28670) );
  XNOR U133 ( .A(n29476), .B(n29466), .Z(n29475) );
  XNOR U134 ( .A(n27101), .B(n27097), .Z(n27100) );
  XNOR U135 ( .A(n29258), .B(n29254), .Z(n29257) );
  XNOR U136 ( .A(n29499), .B(n29486), .Z(n29220) );
  XOR U137 ( .A(n29623), .B(n29614), .Z(n29567) );
  OR U138 ( .A(n27794), .B(n27647), .Z(n27793) );
  NOR U139 ( .A(n27872), .B(n27871), .Z(n27868) );
  NOR U140 ( .A(n28692), .B(n28691), .Z(n28688) );
  XNOR U141 ( .A(n28561), .B(n28548), .Z(n28450) );
  XNOR U142 ( .A(n29289), .B(n29276), .Z(n29190) );
  XOR U143 ( .A(n29147), .B(n29143), .Z(n29135) );
  XNOR U144 ( .A(n27355), .B(n27342), .Z(n26959) );
  XOR U145 ( .A(n27052), .B(n27063), .Z(n26896) );
  XOR U146 ( .A(n27733), .B(n27937), .Z(n27656) );
  AND U147 ( .A(n26971), .B(n26970), .Z(n26968) );
  XOR U148 ( .A(n28793), .B(n28780), .Z(n28481) );
  XOR U149 ( .A(n28445), .B(n28518), .Z(n28452) );
  XNOR U150 ( .A(n27044), .B(n27417), .Z(n27036) );
  AND U151 ( .A(n27011), .B(n27010), .Z(n27008) );
  XOR U152 ( .A(n27134), .B(n27154), .Z(n26953) );
  XNOR U153 ( .A(n27682), .B(n27620), .Z(n26082) );
  XNOR U154 ( .A(n25571), .B(n24466), .Z(n24504) );
  XNOR U155 ( .A(n26365), .B(n26355), .Z(n26362) );
  XNOR U156 ( .A(n29080), .B(n29140), .Z(n25545) );
  XNOR U157 ( .A(n25311), .B(n25301), .Z(n25308) );
  XOR U158 ( .A(n28635), .B(n28631), .Z(n28442) );
  XNOR U159 ( .A(n26160), .B(n26163), .Z(n26186) );
  XNOR U160 ( .A(n26603), .B(n26769), .Z(n26779) );
  XOR U161 ( .A(n25846), .B(n26387), .Z(n25857) );
  XNOR U162 ( .A(n25737), .B(n25871), .Z(n25881) );
  XOR U163 ( .A(n25460), .B(n25451), .Z(n24869) );
  XOR U164 ( .A(n26815), .B(n26806), .Z(n26642) );
  XNOR U165 ( .A(n24601), .B(n24600), .Z(n24599) );
  XOR U166 ( .A(n24944), .B(n25426), .Z(n24762) );
  ANDN U167 ( .B(n25830), .A(n26344), .Z(n25836) );
  XOR U168 ( .A(n25265), .B(n24889), .Z(n25276) );
  ANDN U169 ( .B(n24887), .A(n25291), .Z(n25280) );
  XNOR U170 ( .A(n25634), .B(n25624), .Z(n25631) );
  ANDN U171 ( .B(n23973), .A(n24385), .Z(n23979) );
  XOR U172 ( .A(n25895), .B(n25923), .Z(n25772) );
  XNOR U173 ( .A(n21577), .B(n21567), .Z(n21574) );
  XNOR U174 ( .A(n22142), .B(n22132), .Z(n22139) );
  XNOR U175 ( .A(n24860), .B(n24902), .Z(n21519) );
  XOR U176 ( .A(n23855), .B(n24086), .Z(n21391) );
  XNOR U177 ( .A(n22202), .B(n21241), .Z(n26698) );
  XOR U178 ( .A(n23970), .B(n23987), .Z(n23902) );
  XOR U179 ( .A(n24038), .B(n24066), .Z(n23915) );
  XNOR U180 ( .A(n23343), .B(n23333), .Z(n23340) );
  XNOR U181 ( .A(n26607), .B(n26608), .Z(n26606) );
  XNOR U182 ( .A(n23422), .B(n23414), .Z(n23425) );
  XNOR U183 ( .A(n21033), .B(n21632), .Z(n21042) );
  XNOR U184 ( .A(n21073), .B(n21190), .Z(n21065) );
  XOR U185 ( .A(n23705), .B(n25656), .Z(n25614) );
  ANDN U186 ( .B(n25587), .A(n25586), .Z(n23698) );
  XNOR U187 ( .A(n21337), .B(n21340), .Z(n21366) );
  XNOR U188 ( .A(key[272]), .B(n21541), .Z(n21537) );
  ANDN U189 ( .B(n21902), .A(n22446), .Z(n22440) );
  NANDN U190 ( .A(n22923), .B(n22900), .Z(n22879) );
  NANDN U191 ( .A(n23324), .B(n23170), .Z(n22868) );
  XOR U192 ( .A(n21899), .B(n22424), .Z(n21906) );
  XOR U193 ( .A(n23644), .B(n23638), .Z(n23565) );
  ANDN U194 ( .B(n21926), .A(n21982), .Z(n21893) );
  XOR U195 ( .A(n22897), .B(n22907), .Z(n22765) );
  XNOR U196 ( .A(n18409), .B(n18399), .Z(n18406) );
  XNOR U197 ( .A(n18541), .B(n18531), .Z(n18538) );
  XNOR U198 ( .A(n18267), .B(n18257), .Z(n18264) );
  XNOR U199 ( .A(n19999), .B(n18471), .Z(n18510) );
  XNOR U200 ( .A(n20072), .B(n20062), .Z(n20069) );
  XOR U201 ( .A(n22781), .B(n22834), .Z(n22682) );
  XNOR U202 ( .A(n18648), .B(n18646), .Z(n18642) );
  XOR U203 ( .A(n18242), .B(n18241), .Z(n18240) );
  XNOR U204 ( .A(key[504]), .B(n18385), .Z(n18384) );
  XNOR U205 ( .A(n19430), .B(n20006), .Z(n23606) );
  XNOR U206 ( .A(n19809), .B(n20254), .Z(n19814) );
  NANDN U207 ( .A(n18119), .B(n18095), .Z(n17982) );
  XOR U208 ( .A(n20735), .B(n20727), .Z(n20745) );
  AND U209 ( .A(n18536), .B(n18089), .Z(n18527) );
  XOR U210 ( .A(n19460), .B(n19451), .Z(n18836) );
  XOR U211 ( .A(n19898), .B(n19708), .Z(n19916) );
  XNOR U212 ( .A(n18961), .B(n19315), .Z(n18887) );
  NANDN U213 ( .A(n19309), .B(n18973), .Z(n18963) );
  XNOR U214 ( .A(n20580), .B(n20688), .Z(n20697) );
  NOR U215 ( .A(n19852), .B(n20047), .Z(n19877) );
  XNOR U216 ( .A(n17985), .B(n17991), .Z(n17922) );
  XOR U217 ( .A(n20561), .B(n20776), .Z(n20668) );
  XNOR U218 ( .A(n19888), .B(n20306), .Z(n19802) );
  XNOR U219 ( .A(n17185), .B(n17175), .Z(n17182) );
  XOR U220 ( .A(n17284), .B(n15190), .Z(n16208) );
  XOR U221 ( .A(n16219), .B(n17279), .Z(n15163) );
  XOR U222 ( .A(n16177), .B(n16207), .Z(n15189) );
  XNOR U223 ( .A(n19841), .B(n19903), .Z(n19672) );
  NANDN U224 ( .A(n20790), .B(n20725), .Z(n20638) );
  XOR U225 ( .A(n20629), .B(n22582), .Z(n20623) );
  XOR U226 ( .A(n19804), .B(n19816), .Z(n19787) );
  XNOR U227 ( .A(n19745), .B(n19744), .Z(n15584) );
  XOR U228 ( .A(n20620), .B(n20621), .Z(n20583) );
  XNOR U229 ( .A(n16511), .B(n16957), .Z(n16954) );
  XOR U230 ( .A(n20641), .B(n20791), .Z(n20635) );
  XNOR U231 ( .A(n17566), .B(n17726), .Z(n17736) );
  XOR U232 ( .A(n16120), .B(n16111), .Z(n15791) );
  XNOR U233 ( .A(n17573), .B(n18767), .Z(n18673) );
  XOR U234 ( .A(n15162), .B(n16195), .Z(n17918) );
  XNOR U235 ( .A(n20520), .B(n20523), .Z(n20598) );
  ANDN U236 ( .B(n17684), .A(n17751), .Z(n17710) );
  XNOR U237 ( .A(n16399), .B(n16489), .Z(n16406) );
  XNOR U238 ( .A(n15949), .B(n15865), .Z(n15861) );
  XOR U239 ( .A(n16283), .B(n16274), .Z(n15885) );
  AND U240 ( .A(n15378), .B(n15030), .Z(n15369) );
  NANDN U241 ( .A(n17008), .B(n17002), .Z(n16804) );
  XOR U242 ( .A(n15967), .B(n15957), .Z(n15781) );
  ANDN U243 ( .B(n15936), .A(n15935), .Z(n15802) );
  XOR U244 ( .A(n16843), .B(n16854), .Z(n16660) );
  XOR U245 ( .A(n16816), .B(n16827), .Z(n16666) );
  XNOR U246 ( .A(n14063), .B(n14053), .Z(n14060) );
  XOR U247 ( .A(n12603), .B(n14297), .Z(n12583) );
  XNOR U248 ( .A(n13976), .B(n13537), .Z(n12142) );
  XNOR U249 ( .A(n13150), .B(n13140), .Z(n13147) );
  XNOR U250 ( .A(key[713]), .B(n13127), .Z(n14159) );
  XNOR U251 ( .A(key[665]), .B(n13412), .Z(n14424) );
  XOR U252 ( .A(n13531), .B(n12153), .Z(n14001) );
  XNOR U253 ( .A(n16628), .B(n16631), .Z(n16710) );
  XOR U254 ( .A(n13252), .B(n12625), .Z(n15033) );
  XOR U255 ( .A(key[647]), .B(n12311), .Z(n17577) );
  XOR U256 ( .A(key[727]), .B(n12497), .Z(n15771) );
  XOR U257 ( .A(n14337), .B(n14328), .Z(n13717) );
  AND U258 ( .A(n14198), .B(n14183), .Z(n14189) );
  XOR U259 ( .A(n12385), .B(n12372), .Z(n11903) );
  NANDN U260 ( .A(n14675), .B(n14676), .Z(n14626) );
  ANDN U261 ( .B(n13273), .A(n13279), .Z(n12987) );
  XOR U262 ( .A(n11986), .B(n12003), .Z(n11875) );
  XOR U263 ( .A(n14640), .B(n17421), .Z(n14647) );
  ANDN U264 ( .B(n14645), .A(n17443), .Z(n17441) );
  XNOR U265 ( .A(n9067), .B(n9057), .Z(n9064) );
  ANDN U266 ( .B(n12912), .A(n13002), .Z(n12860) );
  XOR U267 ( .A(n13270), .B(n13289), .Z(n12844) );
  XNOR U268 ( .A(n9200), .B(n9190), .Z(n9197) );
  XNOR U269 ( .A(n14545), .B(n14612), .Z(n9614) );
  XOR U270 ( .A(n10351), .B(n10961), .Z(n10337) );
  XOR U271 ( .A(n9260), .B(n10201), .Z(n11157) );
  XNOR U272 ( .A(n10968), .B(n11816), .Z(n10983) );
  XNOR U273 ( .A(n9841), .B(n10390), .Z(n10382) );
  AND U274 ( .A(n9062), .B(n8974), .Z(n9053) );
  XOR U275 ( .A(key[800]), .B(n11144), .Z(n11142) );
  XNOR U276 ( .A(n10061), .B(n10045), .Z(n11259) );
  XOR U277 ( .A(n12704), .B(n12695), .Z(n11616) );
  XOR U278 ( .A(n9015), .B(n9222), .Z(n9026) );
  XNOR U279 ( .A(n10467), .B(n10470), .Z(n10494) );
  XNOR U280 ( .A(n10882), .B(n10869), .Z(n10802) );
  ANDN U281 ( .B(n10766), .A(n11300), .Z(n10792) );
  XOR U282 ( .A(n10418), .B(n10409), .Z(n9835) );
  ANDN U283 ( .B(n8931), .A(n9491), .Z(n8986) );
  XOR U284 ( .A(n9905), .B(n9922), .Z(n9806) );
  NANDN U285 ( .A(n10083), .B(n9853), .Z(n9883) );
  XOR U286 ( .A(n11064), .B(n11055), .Z(n10740) );
  XNOR U287 ( .A(n11753), .B(n11740), .Z(n11641) );
  XOR U288 ( .A(n8860), .B(n9480), .Z(n8832) );
  XNOR U289 ( .A(n10569), .B(n10559), .Z(n10566) );
  XOR U290 ( .A(n6106), .B(n6139), .Z(n9846) );
  XNOR U291 ( .A(n6152), .B(n8225), .Z(n7058) );
  XNOR U292 ( .A(n8874), .B(n8949), .Z(n6580) );
  XNOR U293 ( .A(n11523), .B(n11504), .Z(n6276) );
  XNOR U294 ( .A(n6202), .B(n6192), .Z(n6199) );
  XNOR U295 ( .A(n7721), .B(n8016), .Z(n7998) );
  XNOR U296 ( .A(n6442), .B(n10751), .Z(n10750) );
  XNOR U297 ( .A(n10648), .B(n10631), .Z(n6416) );
  XOR U298 ( .A(n11493), .B(n11487), .Z(n11498) );
  XOR U299 ( .A(n10540), .B(n10591), .Z(n10549) );
  XOR U300 ( .A(n6158), .B(n6224), .Z(n6178) );
  ANDN U301 ( .B(n7811), .A(n8267), .Z(n7800) );
  XOR U302 ( .A(n8725), .B(n8776), .Z(n8734) );
  ANDN U303 ( .B(n8715), .A(n8739), .Z(n8611) );
  XOR U304 ( .A(n6394), .B(n6388), .Z(n6399) );
  NANDN U305 ( .A(n6183), .B(n6161), .Z(n5916) );
  ANDN U306 ( .B(n6900), .A(n7241), .Z(n6926) );
  XOR U307 ( .A(n7394), .B(n7385), .Z(n6771) );
  XNOR U308 ( .A(n4958), .B(n2993), .Z(n3006) );
  XOR U309 ( .A(n8494), .B(n8495), .Z(n8657) );
  XNOR U310 ( .A(n5006), .B(n4996), .Z(n5003) );
  XOR U311 ( .A(n3654), .B(n3554), .Z(n3676) );
  XNOR U312 ( .A(n6731), .B(n6730), .Z(n4084) );
  XNOR U313 ( .A(n2907), .B(n2897), .Z(n2904) );
  XNOR U314 ( .A(n2582), .B(n2572), .Z(n2579) );
  XNOR U315 ( .A(n3002), .B(n2981), .Z(n4268) );
  NANDN U316 ( .A(n3967), .B(n3633), .Z(n3638) );
  XOR U317 ( .A(n5145), .B(n5136), .Z(n4814) );
  ANDN U318 ( .B(n4732), .A(n5247), .Z(n4783) );
  AND U319 ( .A(n3833), .B(n3613), .Z(n3824) );
  ANDN U320 ( .B(n2459), .A(n3027), .Z(n2848) );
  XOR U321 ( .A(n1705), .B(n3497), .Z(n3489) );
  XNOR U322 ( .A(n849), .B(n850), .Z(n848) );
  XNOR U323 ( .A(n591), .B(n594), .Z(n617) );
  XOR U324 ( .A(key[1204]), .B(n420), .Z(n419) );
  XNOR U325 ( .A(n4548), .B(n4538), .Z(n4545) );
  XOR U326 ( .A(n895), .B(n890), .Z(n441) );
  XOR U327 ( .A(n1932), .B(n1927), .Z(n1916) );
  XOR U328 ( .A(n1732), .B(n1727), .Z(n1715) );
  XOR U329 ( .A(n1529), .B(n1524), .Z(n1513) );
  XOR U330 ( .A(n1307), .B(n1302), .Z(n1291) );
  XOR U331 ( .A(n1102), .B(n1097), .Z(n1086) );
  XOR U332 ( .A(n876), .B(n871), .Z(n860) );
  XOR U333 ( .A(n464), .B(n459), .Z(n446) );
  XOR U334 ( .A(n253), .B(n248), .Z(n237) );
  XOR U335 ( .A(n38), .B(n33), .Z(n22) );
  XOR U336 ( .A(n4288), .B(n4283), .Z(n3387) );
  XOR U337 ( .A(n3207), .B(n3202), .Z(n3191) );
  XOR U338 ( .A(n2187), .B(n2182), .Z(n2171) );
  XNOR U339 ( .A(n27794), .B(n27646), .Z(n28177) );
  XNOR U340 ( .A(n27947), .B(n27713), .Z(n27997) );
  XNOR U341 ( .A(n29179), .B(n29098), .Z(n29414) );
  XNOR U342 ( .A(n29622), .B(n29612), .Z(n29619) );
  XOR U343 ( .A(n29489), .B(n29503), .Z(n29500) );
  XOR U344 ( .A(n27257), .B(n27271), .Z(n27268) );
  XNOR U345 ( .A(n28639), .B(n28400), .Z(n28909) );
  XOR U346 ( .A(n28551), .B(n28565), .Z(n28562) );
  XNOR U347 ( .A(n27423), .B(n26944), .Z(n27459) );
  XOR U348 ( .A(n29279), .B(n29293), .Z(n29290) );
  XOR U349 ( .A(n27345), .B(n27359), .Z(n27356) );
  XOR U350 ( .A(n27168), .B(n27183), .Z(n27180) );
  XNOR U351 ( .A(n28121), .B(n28119), .Z(n28107) );
  XNOR U352 ( .A(n27852), .B(n27837), .Z(n27850) );
  XNOR U353 ( .A(n27075), .B(n27071), .Z(n27074) );
  XNOR U354 ( .A(n28531), .B(n28526), .Z(n28530) );
  XOR U355 ( .A(n28783), .B(n28797), .Z(n28794) );
  XNOR U356 ( .A(n28772), .B(n28761), .Z(n28770) );
  XNOR U357 ( .A(n27173), .B(n27162), .Z(n27164) );
  XOR U358 ( .A(n28159), .B(n28150), .Z(n27675) );
  XOR U359 ( .A(n28068), .B(n28059), .Z(n27663) );
  XOR U360 ( .A(n27873), .B(n27860), .Z(n27637) );
  XNOR U361 ( .A(n28693), .B(n28680), .Z(n28492) );
  XOR U362 ( .A(n27980), .B(n27971), .Z(n27707) );
  NOR U363 ( .A(n27266), .B(n27265), .Z(n27262) );
  NOR U364 ( .A(n28560), .B(n28559), .Z(n28556) );
  XOR U365 ( .A(n27442), .B(n27433), .Z(n26997) );
  XOR U366 ( .A(n29397), .B(n29388), .Z(n29092) );
  AND U367 ( .A(n29220), .B(n29219), .Z(n29216) );
  XOR U368 ( .A(n29351), .B(n29574), .Z(n29172) );
  XNOR U369 ( .A(n27613), .B(n27611), .Z(n27670) );
  NOR U370 ( .A(n27178), .B(n27177), .Z(n27174) );
  XOR U371 ( .A(n29185), .B(n29245), .Z(n29193) );
  XOR U372 ( .A(n29157), .B(n29153), .Z(n29082) );
  XOR U373 ( .A(n28426), .B(n28422), .Z(n28354) );
  XOR U374 ( .A(n28892), .B(n28883), .Z(n28629) );
  NOR U375 ( .A(n28792), .B(n28791), .Z(n28788) );
  XOR U376 ( .A(n27078), .B(n27089), .Z(n27032) );
  AND U377 ( .A(n26959), .B(n26958), .Z(n26956) );
  XNOR U378 ( .A(n26881), .B(n26966), .Z(n26309) );
  AND U379 ( .A(n29190), .B(n29268), .Z(n29266) );
  XOR U380 ( .A(n25221), .B(n25220), .Z(n24202) );
  XNOR U381 ( .A(n27531), .B(n27521), .Z(n27528) );
  XNOR U382 ( .A(n26992), .B(n27003), .Z(n26905) );
  XNOR U383 ( .A(n24129), .B(n24119), .Z(n24126) );
  XNOR U384 ( .A(n26239), .B(n26229), .Z(n26236) );
  XNOR U385 ( .A(n29182), .B(n29102), .Z(n24488) );
  XNOR U386 ( .A(n25985), .B(n25975), .Z(n25982) );
  XNOR U387 ( .A(n27629), .B(n27628), .Z(n25212) );
  XNOR U388 ( .A(n25142), .B(n25132), .Z(n25139) );
  XNOR U389 ( .A(n24875), .B(n25433), .Z(n25425) );
  XNOR U390 ( .A(n24405), .B(n24395), .Z(n24402) );
  XOR U391 ( .A(n24504), .B(n24503), .Z(n24502) );
  XOR U392 ( .A(n24915), .B(n24900), .Z(n24926) );
  XNOR U393 ( .A(n25509), .B(n25512), .Z(n25539) );
  XNOR U394 ( .A(key[239]), .B(n24353), .Z(n26175) );
  XNOR U395 ( .A(n26663), .B(n28227), .Z(n28237) );
  XNOR U396 ( .A(n23880), .B(n24014), .Z(n24023) );
  XNOR U397 ( .A(n24541), .B(n24531), .Z(n24538) );
  XOR U398 ( .A(n26290), .B(n26283), .Z(n26295) );
  XOR U399 ( .A(n25947), .B(n26007), .Z(n25965) );
  XOR U400 ( .A(n24644), .B(n24626), .Z(n26336) );
  XOR U401 ( .A(n28996), .B(n28987), .Z(n26673) );
  XNOR U402 ( .A(n24803), .B(n24968), .Z(n24977) );
  XOR U403 ( .A(n23989), .B(n23975), .Z(n24000) );
  XOR U404 ( .A(n26154), .B(n26163), .Z(n26173) );
  XOR U405 ( .A(n24068), .B(n24043), .Z(n24079) );
  XOR U406 ( .A(n25013), .B(n25004), .Z(n24838) );
  XNOR U407 ( .A(n24235), .B(n24234), .Z(n24233) );
  XOR U408 ( .A(n24090), .B(n23885), .Z(n24108) );
  ANDN U409 ( .B(n26731), .A(n27510), .Z(n26726) );
  XOR U410 ( .A(n28273), .B(n28263), .Z(n26656) );
  NANDN U411 ( .A(n24098), .B(n23953), .Z(n24050) );
  ANDN U412 ( .B(n25898), .A(n26218), .Z(n25940) );
  XOR U413 ( .A(n26111), .B(n26102), .Z(n25766) );
  NANDN U414 ( .A(n25955), .B(n25811), .Z(n25906) );
  XOR U415 ( .A(n24264), .B(n24255), .Z(n23909) );
  XOR U416 ( .A(n24884), .B(n25263), .Z(n24831) );
  XNOR U417 ( .A(n26501), .B(n26491), .Z(n26498) );
  XNOR U418 ( .A(n24773), .B(n25417), .Z(n22569) );
  XNOR U419 ( .A(n23414), .B(n22082), .Z(n21654) );
  XNOR U420 ( .A(n21135), .B(n21125), .Z(n21132) );
  ANDN U421 ( .B(n24041), .A(n24521), .Z(n24083) );
  XNOR U422 ( .A(n25753), .B(n26342), .Z(n25775) );
  XOR U423 ( .A(n25827), .B(n25844), .Z(n25759) );
  XNOR U424 ( .A(n24937), .B(n24891), .Z(n23309) );
  XNOR U425 ( .A(n23777), .B(n23767), .Z(n23774) );
  XNOR U426 ( .A(n24698), .B(n24688), .Z(n24695) );
  XNOR U427 ( .A(n23920), .B(n23919), .Z(n21388) );
  XNOR U428 ( .A(n22302), .B(n22291), .Z(n22299) );
  XNOR U429 ( .A(n23158), .B(n22385), .Z(n21357) );
  XOR U430 ( .A(key[276]), .B(n21527), .Z(n21523) );
  XNOR U431 ( .A(n20969), .B(n21428), .Z(n21410) );
  XNOR U432 ( .A(n21495), .B(n21502), .Z(n21503) );
  XNOR U433 ( .A(n26581), .B(n26704), .Z(n23022) );
  XNOR U434 ( .A(n22008), .B(n21998), .Z(n22005) );
  XOR U435 ( .A(n23689), .B(n26523), .Z(n26481) );
  XNOR U436 ( .A(n22989), .B(n22992), .Z(n23016) );
  XOR U437 ( .A(n21513), .B(n22575), .Z(n23318) );
  XNOR U438 ( .A(n23875), .B(n22376), .Z(n23128) );
  NANDN U439 ( .A(n23693), .B(n23694), .Z(n23667) );
  XOR U440 ( .A(n23613), .B(n23718), .Z(n23747) );
  XNOR U441 ( .A(key[368]), .B(n21358), .Z(n24058) );
  XOR U442 ( .A(n23627), .B(n23648), .Z(n24668) );
  XNOR U443 ( .A(key[288]), .B(n21664), .Z(n25915) );
  XOR U444 ( .A(n21057), .B(n21073), .Z(n21083) );
  XOR U445 ( .A(n21241), .B(n21242), .Z(n21240) );
  XNOR U446 ( .A(n20989), .B(n21260), .Z(n21252) );
  XOR U447 ( .A(n21446), .B(n21436), .Z(n20963) );
  XNOR U448 ( .A(n22669), .B(n22906), .Z(n22914) );
  XOR U449 ( .A(n21023), .B(n21033), .Z(n21049) );
  ANDN U450 ( .B(n21031), .A(n21556), .Z(n21026) );
  XOR U451 ( .A(n23180), .B(n23172), .Z(n23190) );
  XNOR U452 ( .A(n22707), .B(n22857), .Z(n22852) );
  XNOR U453 ( .A(n23216), .B(n23207), .Z(n22717) );
  NOR U454 ( .A(n23752), .B(n23756), .Z(n23617) );
  ANDN U455 ( .B(n24673), .A(n24677), .Z(n23631) );
  NANDN U456 ( .A(n22261), .B(n21920), .Z(n22249) );
  XOR U457 ( .A(n25574), .B(n25605), .Z(n23581) );
  XNOR U458 ( .A(n21889), .B(n21885), .Z(n21802) );
  XNOR U459 ( .A(n22443), .B(n22439), .Z(n21861) );
  XOR U460 ( .A(n21024), .B(n21550), .Z(n20973) );
  XOR U461 ( .A(n21288), .B(n21279), .Z(n20982) );
  NANDN U462 ( .A(n21256), .B(n21090), .Z(n21100) );
  ANDN U463 ( .B(n22870), .A(n22869), .Z(n22867) );
  XOR U464 ( .A(n23068), .B(n23058), .Z(n22701) );
  XNOR U465 ( .A(n19038), .B(n19028), .Z(n19035) );
  XNOR U466 ( .A(n19198), .B(n19188), .Z(n19195) );
  XNOR U467 ( .A(n23603), .B(n23602), .Z(n18493) );
  XOR U468 ( .A(n21808), .B(n21809), .Z(n21872) );
  XNOR U469 ( .A(key[384]), .B(n18518), .Z(n18514) );
  XOR U470 ( .A(n18339), .B(n20439), .Z(n19531) );
  XNOR U471 ( .A(key[424]), .B(n18658), .Z(n18657) );
  XNOR U472 ( .A(n19937), .B(n19927), .Z(n19934) );
  XNOR U473 ( .A(n20972), .B(n20937), .Z(n18645) );
  XNOR U474 ( .A(n22746), .B(n22747), .Z(n22745) );
  XNOR U475 ( .A(n22692), .B(n22763), .Z(n20296) );
  XNOR U476 ( .A(n20199), .B(n20189), .Z(n20196) );
  XNOR U477 ( .A(key[464]), .B(n18243), .Z(n18239) );
  XOR U478 ( .A(key[500]), .B(n20410), .Z(n20421) );
  XOR U479 ( .A(n18479), .B(n20017), .Z(n20012) );
  XOR U480 ( .A(n18513), .B(n19998), .Z(n19994) );
  XNOR U481 ( .A(n22658), .B(n20258), .Z(n20287) );
  ANDN U482 ( .B(n18922), .A(n19172), .Z(n19147) );
  XOR U483 ( .A(n19863), .B(n19855), .Z(n19874) );
  XOR U484 ( .A(n18236), .B(n20259), .Z(n20255) );
  XOR U485 ( .A(n19334), .B(n19325), .Z(n18844) );
  XNOR U486 ( .A(n21771), .B(n21852), .Z(n21791) );
  XNOR U487 ( .A(n23486), .B(n23477), .Z(n20609) );
  ANDN U488 ( .B(n18002), .A(n18394), .Z(n17928) );
  XOR U489 ( .A(n18066), .B(n18077), .Z(n17976) );
  XOR U490 ( .A(n18092), .B(n18103), .Z(n17921) );
  NANDN U491 ( .A(n18247), .B(n18030), .Z(n17940) );
  XOR U492 ( .A(n20348), .B(n20335), .Z(n19800) );
  XNOR U493 ( .A(n18887), .B(n18886), .Z(n18775) );
  XOR U494 ( .A(n19818), .B(n19809), .Z(n19829) );
  XOR U495 ( .A(n18801), .B(n18796), .Z(n18773) );
  XOR U496 ( .A(n17999), .B(n18011), .Z(n17972) );
  AND U497 ( .A(n18055), .B(n18056), .Z(n18053) );
  NOR U498 ( .A(n18959), .B(n18958), .Z(n18955) );
  XNOR U499 ( .A(n17922), .B(n17836), .Z(n17264) );
  XNOR U500 ( .A(n17943), .B(n18248), .Z(n17937) );
  XNOR U501 ( .A(n19801), .B(n19802), .Z(n19723) );
  XNOR U502 ( .A(n18712), .B(n18702), .Z(n18709) );
  NANDN U503 ( .A(n22581), .B(n20681), .Z(n20626) );
  XNOR U504 ( .A(n19880), .B(n19876), .Z(n19764) );
  XNOR U505 ( .A(n15248), .B(n15238), .Z(n15245) );
  XNOR U506 ( .A(n18903), .B(n18902), .Z(n15467) );
  XNOR U507 ( .A(n15076), .B(n15066), .Z(n15073) );
  XOR U508 ( .A(n16032), .B(n17101), .Z(n15307) );
  XNOR U509 ( .A(n20762), .B(n20768), .Z(n20652) );
  XNOR U510 ( .A(n17041), .B(n17031), .Z(n17038) );
  XNOR U511 ( .A(n16434), .B(n16424), .Z(n16431) );
  XNOR U512 ( .A(n17556), .B(n17692), .Z(n17702) );
  XNOR U513 ( .A(n17826), .B(n17829), .Z(n17906) );
  XOR U514 ( .A(n19672), .B(n19671), .Z(n19667) );
  XNOR U515 ( .A(n19605), .B(n19595), .Z(n19602) );
  XOR U516 ( .A(n20722), .B(n20733), .Z(n20675) );
  XOR U517 ( .A(n20678), .B(n20689), .Z(n20671) );
  XNOR U518 ( .A(n19683), .B(n19786), .Z(n16382) );
  XNOR U519 ( .A(n15346), .B(n16064), .Z(n17132) );
  XNOR U520 ( .A(n16336), .B(n16340), .Z(n16335) );
  XNOR U521 ( .A(n15523), .B(n15513), .Z(n15520) );
  XNOR U522 ( .A(n16692), .B(n16853), .Z(n16862) );
  XNOR U523 ( .A(n16706), .B(n16826), .Z(n16835) );
  XOR U524 ( .A(n18682), .B(n17573), .Z(n18691) );
  XOR U525 ( .A(n19575), .B(n17676), .Z(n19584) );
  XOR U526 ( .A(n15056), .B(n15098), .Z(n15071) );
  XOR U527 ( .A(n15457), .B(n16530), .Z(n18994) );
  XOR U528 ( .A(n14959), .B(n14969), .Z(n14985) );
  XOR U529 ( .A(n17777), .B(n17768), .Z(n17595) );
  XOR U530 ( .A(n15911), .B(n16399), .Z(n16413) );
  XNOR U531 ( .A(n16172), .B(n16200), .Z(n15844) );
  XOR U532 ( .A(n15207), .B(n15270), .Z(n15218) );
  ANDN U533 ( .B(n15012), .A(n15359), .Z(n15007) );
  XOR U534 ( .A(n15384), .B(n15375), .Z(n14869) );
  NANDN U535 ( .A(n16883), .B(n16846), .Z(n16729) );
  XOR U536 ( .A(n16899), .B(n16890), .Z(n16685) );
  NANDN U537 ( .A(n17293), .B(n16819), .Z(n16741) );
  XOR U538 ( .A(n17309), .B(n17300), .Z(n16699) );
  XOR U539 ( .A(n20514), .B(n20523), .Z(n20543) );
  XOR U540 ( .A(n20471), .B(n20462), .Z(n17585) );
  XOR U541 ( .A(n17143), .B(n17163), .Z(n16708) );
  XOR U542 ( .A(n15793), .B(n15788), .Z(n15745) );
  ANDN U543 ( .B(n17718), .A(n20445), .Z(n17744) );
  XNOR U544 ( .A(n15886), .B(n15881), .Z(n15757) );
  ANDN U545 ( .B(n14967), .A(n15498), .Z(n14962) );
  XOR U546 ( .A(n15783), .B(n15778), .Z(n15750) );
  XOR U547 ( .A(key[687]), .B(n12612), .Z(n14860) );
  XNOR U548 ( .A(n14749), .B(n14739), .Z(n14746) );
  XNOR U549 ( .A(n17524), .B(n18669), .Z(n12309) );
  XOR U550 ( .A(n12268), .B(n13408), .Z(n14406) );
  XNOR U551 ( .A(n17609), .B(n17549), .Z(n14393) );
  XNOR U552 ( .A(n17462), .B(n17452), .Z(n17459) );
  XNOR U553 ( .A(n15668), .B(n15657), .Z(n15665) );
  XNOR U554 ( .A(n13900), .B(n13890), .Z(n13897) );
  XNOR U555 ( .A(n11860), .B(n11963), .Z(n11973) );
  XNOR U556 ( .A(n13312), .B(n13301), .Z(n13309) );
  XNOR U557 ( .A(n16722), .B(n16723), .Z(n16774) );
  XNOR U558 ( .A(n11842), .B(n12332), .Z(n12327) );
  XNOR U559 ( .A(n15730), .B(n15887), .Z(n12495) );
  XNOR U560 ( .A(n15799), .B(n15798), .Z(n13103) );
  XNOR U561 ( .A(n12254), .B(n12278), .Z(n12262) );
  XOR U562 ( .A(n12068), .B(n12059), .Z(n11884) );
  XOR U563 ( .A(key[642]), .B(n13382), .Z(n17520) );
  XOR U564 ( .A(key[767]), .B(n12170), .Z(n16653) );
  XNOR U565 ( .A(n13021), .B(n13011), .Z(n13018) );
  XOR U566 ( .A(n12935), .B(n12914), .Z(n12949) );
  XNOR U567 ( .A(n12834), .B(n13430), .Z(n13438) );
  XNOR U568 ( .A(n14588), .B(n16551), .Z(n16547) );
  XOR U569 ( .A(n13463), .B(n13454), .Z(n12876) );
  XOR U570 ( .A(n12528), .B(n12519), .Z(n11915) );
  XOR U571 ( .A(n13702), .B(n13869), .Z(n13757) );
  AND U572 ( .A(n14744), .B(n14729), .Z(n14735) );
  XOR U573 ( .A(n14611), .B(n15648), .Z(n15663) );
  XNOR U574 ( .A(n12202), .B(n12193), .Z(n11874) );
  XOR U575 ( .A(n17423), .B(n14646), .Z(n17434) );
  XOR U576 ( .A(n13291), .B(n13275), .Z(n13307) );
  NANDN U577 ( .A(n14703), .B(n14704), .Z(n14698) );
  XOR U578 ( .A(n16579), .B(n16570), .Z(n14689) );
  NOR U579 ( .A(n14317), .B(n14316), .Z(n14313) );
  ANDN U580 ( .B(n13852), .A(n13851), .Z(n13834) );
  XOR U581 ( .A(n14204), .B(n14195), .Z(n13841) );
  XOR U582 ( .A(n13151), .B(n13138), .Z(n12850) );
  XOR U583 ( .A(n11897), .B(n12352), .Z(n11904) );
  XNOR U584 ( .A(n14004), .B(n14043), .Z(n13747) );
  XOR U585 ( .A(n12900), .B(n12958), .Z(n12792) );
  XOR U586 ( .A(n10198), .B(n11120), .Z(n9290) );
  XNOR U587 ( .A(n11321), .B(n11311), .Z(n11318) );
  XOR U588 ( .A(n11260), .B(n10051), .Z(n10037) );
  XNOR U589 ( .A(n14523), .B(n14619), .Z(n9612) );
  XNOR U590 ( .A(n9370), .B(n9360), .Z(n9367) );
  XNOR U591 ( .A(n10270), .B(n10260), .Z(n10267) );
  XNOR U592 ( .A(n12857), .B(n12915), .Z(n9259) );
  XNOR U593 ( .A(n10104), .B(n10094), .Z(n10101) );
  XNOR U594 ( .A(key[769]), .B(n9170), .Z(n10067) );
  XOR U595 ( .A(n10189), .B(n11133), .Z(n9286) );
  XNOR U596 ( .A(n11537), .B(n11684), .Z(n11696) );
  XOR U597 ( .A(key[842]), .B(n10369), .Z(n10967) );
  XNOR U598 ( .A(key[881]), .B(n9614), .Z(n11412) );
  XOR U599 ( .A(key[887]), .B(n10504), .Z(n11398) );
  XNOR U600 ( .A(n8930), .B(n9495), .Z(n9487) );
  XOR U601 ( .A(n9321), .B(n9392), .Z(n9341) );
  XOR U602 ( .A(n10221), .B(n10292), .Z(n10241) );
  XNOR U603 ( .A(n9468), .B(n10372), .Z(n10371) );
  XNOR U604 ( .A(n10731), .B(n11012), .Z(n11002) );
  XOR U605 ( .A(n14459), .B(n14450), .Z(n11569) );
  ANDN U606 ( .B(n11623), .A(n12672), .Z(n11716) );
  XOR U607 ( .A(n11186), .B(n11177), .Z(n10724) );
  XOR U608 ( .A(n11548), .B(n12661), .Z(n11506) );
  XOR U609 ( .A(n13600), .B(n13591), .Z(n11600) );
  XOR U610 ( .A(n11636), .B(n11654), .Z(n11582) );
  XOR U611 ( .A(n9523), .B(n9514), .Z(n8924) );
  XOR U612 ( .A(n8938), .B(n8961), .Z(n8896) );
  NANDN U613 ( .A(n9179), .B(n8999), .Z(n9005) );
  XOR U614 ( .A(n8996), .B(n9013), .Z(n8881) );
  AND U615 ( .A(n9044), .B(n8943), .Z(n9042) );
  XOR U616 ( .A(n9875), .B(n10126), .Z(n9895) );
  XNOR U617 ( .A(n10214), .B(n9287), .Z(n10213) );
  XOR U618 ( .A(n8385), .B(n8368), .Z(n11513) );
  ANDN U619 ( .B(n9842), .A(n10386), .Z(n9940) );
  AND U620 ( .A(n9953), .B(n9910), .Z(n9951) );
  XNOR U621 ( .A(n10687), .B(n11298), .Z(n10713) );
  XNOR U622 ( .A(n6590), .B(n7966), .Z(n7341) );
  ANDN U623 ( .B(n10747), .A(n11032), .Z(n10834) );
  XOR U624 ( .A(n10673), .B(n11021), .Z(n10633) );
  XOR U625 ( .A(n10797), .B(n10815), .Z(n10704) );
  XNOR U626 ( .A(n11518), .B(n11516), .Z(n11564) );
  XNOR U627 ( .A(n8288), .B(n8278), .Z(n8285) );
  XNOR U628 ( .A(n8754), .B(n8744), .Z(n8751) );
  XNOR U629 ( .A(n7880), .B(n7870), .Z(n7877) );
  XNOR U630 ( .A(n8375), .B(n7186), .Z(n6293) );
  XOR U631 ( .A(n9770), .B(n10375), .Z(n9742) );
  XNOR U632 ( .A(n9665), .B(n9655), .Z(n9662) );
  XNOR U633 ( .A(n8215), .B(n6134), .Z(n7050) );
  XNOR U634 ( .A(n11442), .B(n11432), .Z(n11439) );
  XNOR U635 ( .A(n6483), .B(n6473), .Z(n6480) );
  XNOR U636 ( .A(n7262), .B(n7252), .Z(n7259) );
  XOR U637 ( .A(n6588), .B(n6545), .Z(n7357) );
  XOR U638 ( .A(key[1019]), .B(n8255), .Z(n9902) );
  XNOR U639 ( .A(n7634), .B(n7780), .Z(n7769) );
  XNOR U640 ( .A(n6808), .B(n6939), .Z(n6958) );
  XNOR U641 ( .A(n6045), .B(n6035), .Z(n6042) );
  XNOR U642 ( .A(n6343), .B(n6333), .Z(n6340) );
  XNOR U643 ( .A(n6825), .B(n7094), .Z(n7084) );
  XNOR U644 ( .A(n7475), .B(n8094), .Z(n10854) );
  XOR U645 ( .A(n8033), .B(n8024), .Z(n7714) );
  ANDN U646 ( .B(n7703), .A(n7849), .Z(n7728) );
  XOR U647 ( .A(n6911), .B(n7284), .Z(n6922) );
  ANDN U648 ( .B(n10530), .A(n10554), .Z(n8699) );
  XOR U649 ( .A(n8681), .B(n8677), .Z(n8695) );
  XOR U650 ( .A(n8155), .B(n8146), .Z(n7671) );
  NANDN U651 ( .A(n8129), .B(n7753), .Z(n7773) );
  XOR U652 ( .A(n6975), .B(n6965), .Z(n6800) );
  XOR U653 ( .A(n5977), .B(n5982), .Z(n5996) );
  XOR U654 ( .A(n7129), .B(n7120), .Z(n6818) );
  XOR U655 ( .A(n8643), .B(n11464), .Z(n8653) );
  ANDN U656 ( .B(n8626), .A(n11423), .Z(n8559) );
  XOR U657 ( .A(n6006), .B(n6011), .Z(n6024) );
  XOR U658 ( .A(n10527), .B(n10538), .Z(n8604) );
  XOR U659 ( .A(n7793), .B(n7809), .Z(n7621) );
  XOR U660 ( .A(key[1113]), .B(n4111), .Z(n4110) );
  NANDN U661 ( .A(n6029), .B(n6009), .Z(n5905) );
  NANDN U662 ( .A(n6327), .B(n5954), .Z(n5868) );
  XOR U663 ( .A(n8552), .B(n8553), .Z(n8710) );
  XOR U664 ( .A(n5811), .B(n6169), .Z(n5943) );
  XNOR U665 ( .A(n5925), .B(n5809), .Z(n5783) );
  XNOR U666 ( .A(n6863), .B(n6870), .Z(n6855) );
  XNOR U667 ( .A(n7540), .B(n7530), .Z(n7537) );
  XNOR U668 ( .A(n2718), .B(n2708), .Z(n2715) );
  XNOR U669 ( .A(n7636), .B(n7635), .Z(n2790) );
  XNOR U670 ( .A(n4621), .B(n4972), .Z(n5051) );
  XNOR U671 ( .A(n8579), .B(n8470), .Z(n4236) );
  XNOR U672 ( .A(n3705), .B(n3695), .Z(n3702) );
  XNOR U673 ( .A(n4006), .B(n3996), .Z(n4003) );
  XNOR U674 ( .A(n4228), .B(n4255), .Z(n4240) );
  XOR U675 ( .A(n5801), .B(n5800), .Z(n5798) );
  ANDN U676 ( .B(n5192), .A(n5110), .Z(n5178) );
  XNOR U677 ( .A(n5880), .B(n5879), .Z(n5804) );
  XNOR U678 ( .A(n5865), .B(n5935), .Z(n5794) );
  XNOR U679 ( .A(n6644), .B(n6634), .Z(n6641) );
  XNOR U680 ( .A(n5491), .B(n5629), .Z(n5638) );
  XNOR U681 ( .A(n6860), .B(n6813), .Z(n3158) );
  XNOR U682 ( .A(n3053), .B(n3043), .Z(n3050) );
  XOR U683 ( .A(n3955), .B(n3548), .Z(n3977) );
  XNOR U684 ( .A(n4632), .B(n4754), .Z(n4769) );
  XNOR U685 ( .A(n4642), .B(n4780), .Z(n4795) );
  XNOR U686 ( .A(n5501), .B(n5662), .Z(n5671) );
  XNOR U687 ( .A(n3624), .B(n4142), .Z(n4132) );
  XOR U688 ( .A(key[1076]), .B(n3796), .Z(n3795) );
  XOR U689 ( .A(n5713), .B(n5704), .Z(n5521) );
  XOR U690 ( .A(n3892), .B(n3890), .Z(n3900) );
  XOR U691 ( .A(n2908), .B(n2895), .Z(n2381) );
  ANDN U692 ( .B(n2512), .A(n2556), .Z(n2538) );
  ANDN U693 ( .B(n5612), .A(n7509), .Z(n6593) );
  ANDN U694 ( .B(n2468), .A(n2692), .Z(n2483) );
  XOR U695 ( .A(n4867), .B(n4858), .Z(n4679) );
  ANDN U696 ( .B(n4742), .A(n4841), .Z(n4757) );
  XOR U697 ( .A(n5007), .B(n4998), .Z(n4622) );
  XOR U698 ( .A(n5273), .B(n5264), .Z(n4669) );
  XOR U699 ( .A(n8414), .B(n8405), .Z(n5531) );
  XOR U700 ( .A(n4176), .B(n4167), .Z(n4125) );
  NANDN U701 ( .A(n3666), .B(n3585), .Z(n3590) );
  XNOR U702 ( .A(n4808), .B(n5122), .Z(n4807) );
  ANDN U703 ( .B(n5576), .A(n6613), .Z(n5584) );
  NANDN U704 ( .A(n8388), .B(n5654), .Z(n5680) );
  XOR U705 ( .A(n3839), .B(n3830), .Z(n3542) );
  XNOR U706 ( .A(n2429), .B(n2472), .Z(n2341) );
  XOR U707 ( .A(n1057), .B(n4447), .Z(n412) );
  XOR U708 ( .A(n2399), .B(n2400), .Z(n2453) );
  XOR U709 ( .A(n2509), .B(n2521), .Z(n2411) );
  XNOR U710 ( .A(n5398), .B(n5388), .Z(n5395) );
  XOR U711 ( .A(n1945), .B(n1506), .Z(n1960) );
  XNOR U712 ( .A(n2035), .B(n2025), .Z(n2032) );
  XOR U713 ( .A(n1985), .B(n1975), .Z(n2000) );
  XNOR U714 ( .A(n1810), .B(n1800), .Z(n1807) );
  XNOR U715 ( .A(n1607), .B(n1597), .Z(n1604) );
  XNOR U716 ( .A(n1384), .B(n1374), .Z(n1381) );
  XOR U717 ( .A(n1334), .B(n1324), .Z(n1349) );
  XNOR U718 ( .A(n1182), .B(n1172), .Z(n1179) );
  XOR U719 ( .A(n1132), .B(n1119), .Z(n1147) );
  XNOR U720 ( .A(n4802), .B(n4711), .Z(n1288) );
  XNOR U721 ( .A(n970), .B(n960), .Z(n967) );
  XNOR U722 ( .A(n804), .B(n828), .Z(n814) );
  XNOR U723 ( .A(n681), .B(n717), .Z(n711) );
  XNOR U724 ( .A(n330), .B(n320), .Z(n327) );
  XOR U725 ( .A(n280), .B(n270), .Z(n295) );
  XNOR U726 ( .A(n118), .B(n108), .Z(n115) );
  XOR U727 ( .A(n68), .B(n55), .Z(n83) );
  XOR U728 ( .A(n3527), .B(n3502), .Z(n3526) );
  ANDN U729 ( .B(n4596), .A(n4493), .Z(n4582) );
  XNOR U730 ( .A(n4691), .B(n4637), .Z(n1266) );
  XNOR U731 ( .A(n4366), .B(n4356), .Z(n4363) );
  XNOR U732 ( .A(n3285), .B(n3275), .Z(n3282) );
  XNOR U733 ( .A(n2265), .B(n2255), .Z(n2262) );
  NANDN U734 ( .A(n5377), .B(n1504), .Z(n1964) );
  NANDN U735 ( .A(n3396), .B(n3166), .Z(n2160) );
  XOR U736 ( .A(n3416), .B(n3407), .Z(n2149) );
  NANDN U737 ( .A(n2014), .B(n1973), .Z(n2004) );
  NANDN U738 ( .A(n1789), .B(n1747), .Z(n1778) );
  NANDN U739 ( .A(n1586), .B(n1544), .Z(n1575) );
  NANDN U740 ( .A(n1363), .B(n1322), .Z(n1353) );
  NANDN U741 ( .A(n1161), .B(n1117), .Z(n1151) );
  NANDN U742 ( .A(n949), .B(n907), .Z(n938) );
  XOR U743 ( .A(n752), .B(n743), .Z(n675) );
  NANDN U744 ( .A(n309), .B(n268), .Z(n299) );
  NANDN U745 ( .A(n97), .B(n53), .Z(n87) );
  NANDN U746 ( .A(n4345), .B(n4303), .Z(n4334) );
  NANDN U747 ( .A(n3264), .B(n3222), .Z(n3253) );
  NANDN U748 ( .A(n2244), .B(n2202), .Z(n2233) );
  XOR U749 ( .A(n665), .B(n1500), .Z(n440) );
  XOR U750 ( .A(n1921), .B(n1969), .Z(n1915) );
  XOR U751 ( .A(n1720), .B(n1743), .Z(n1714) );
  XOR U752 ( .A(n1518), .B(n1540), .Z(n1512) );
  XOR U753 ( .A(n1296), .B(n1318), .Z(n1290) );
  XOR U754 ( .A(n1091), .B(n1113), .Z(n1085) );
  XOR U755 ( .A(n865), .B(n903), .Z(n859) );
  XOR U756 ( .A(n585), .B(n594), .Z(n603) );
  XNOR U757 ( .A(n487), .B(n475), .Z(n445) );
  XOR U758 ( .A(n242), .B(n264), .Z(n236) );
  XOR U759 ( .A(n27), .B(n49), .Z(n21) );
  XOR U760 ( .A(n4473), .B(n4480), .Z(n10) );
  XOR U761 ( .A(n3392), .B(n4299), .Z(n3386) );
  XOR U762 ( .A(n3196), .B(n3218), .Z(n3190) );
  XOR U763 ( .A(n2176), .B(n2198), .Z(n2170) );
  XOR U764 ( .A(n1), .B(n2), .Z(out[9]) );
  XNOR U765 ( .A(n3), .B(n4), .Z(n2) );
  XOR U766 ( .A(key[1161]), .B(n5), .Z(n1) );
  XOR U767 ( .A(n6), .B(n7), .Z(out[99]) );
  XNOR U768 ( .A(n8), .B(n9), .Z(n7) );
  XOR U769 ( .A(n10), .B(n11), .Z(n6) );
  XNOR U770 ( .A(key[1251]), .B(n12), .Z(n11) );
  XNOR U771 ( .A(key[1250]), .B(n13), .Z(out[98]) );
  XOR U772 ( .A(n14), .B(n15), .Z(out[97]) );
  XNOR U773 ( .A(n8), .B(n16), .Z(n15) );
  XNOR U774 ( .A(key[1249]), .B(n12), .Z(n14) );
  XOR U775 ( .A(n17), .B(n18), .Z(out[96]) );
  XNOR U776 ( .A(key[1248]), .B(n19), .Z(n18) );
  XOR U777 ( .A(n20), .B(n21), .Z(out[95]) );
  XOR U778 ( .A(n22), .B(n23), .Z(n20) );
  XNOR U779 ( .A(key[1247]), .B(n24), .Z(n23) );
  XNOR U780 ( .A(n25), .B(n26), .Z(out[94]) );
  XNOR U781 ( .A(key[1246]), .B(n27), .Z(n26) );
  XOR U782 ( .A(n28), .B(n29), .Z(out[93]) );
  XNOR U783 ( .A(n30), .B(n31), .Z(n29) );
  XOR U784 ( .A(n22), .B(n32), .Z(n31) );
  XNOR U785 ( .A(n34), .B(n35), .Z(n33) );
  NANDN U786 ( .A(n36), .B(n37), .Z(n35) );
  XOR U787 ( .A(n39), .B(n40), .Z(n28) );
  XOR U788 ( .A(key[1245]), .B(n41), .Z(n40) );
  ANDN U789 ( .B(n42), .A(n43), .Z(n39) );
  XNOR U790 ( .A(n44), .B(n45), .Z(out[92]) );
  XNOR U791 ( .A(key[1244]), .B(n46), .Z(n45) );
  XOR U792 ( .A(n47), .B(n48), .Z(out[91]) );
  XNOR U793 ( .A(n49), .B(n25), .Z(n48) );
  XNOR U794 ( .A(n50), .B(n51), .Z(n25) );
  XNOR U795 ( .A(n52), .B(n41), .Z(n51) );
  ANDN U796 ( .B(n53), .A(n54), .Z(n41) );
  NOR U797 ( .A(n55), .B(n56), .Z(n52) );
  XNOR U798 ( .A(n57), .B(n58), .Z(n47) );
  XOR U799 ( .A(key[1243]), .B(n59), .Z(n58) );
  XOR U800 ( .A(key[1242]), .B(n44), .Z(out[90]) );
  XNOR U801 ( .A(n24), .B(n60), .Z(n44) );
  IV U802 ( .A(n59), .Z(n24) );
  XNOR U803 ( .A(n61), .B(n62), .Z(out[8]) );
  XNOR U804 ( .A(key[1160]), .B(n63), .Z(n62) );
  XOR U805 ( .A(n64), .B(n21), .Z(out[89]) );
  XNOR U806 ( .A(n50), .B(n65), .Z(n49) );
  XNOR U807 ( .A(n66), .B(n67), .Z(n65) );
  NANDN U808 ( .A(n68), .B(n37), .Z(n67) );
  XNOR U809 ( .A(n32), .B(n69), .Z(n50) );
  XNOR U810 ( .A(n70), .B(n71), .Z(n69) );
  NANDN U811 ( .A(n72), .B(n73), .Z(n71) );
  XOR U812 ( .A(n60), .B(n57), .Z(n27) );
  XNOR U813 ( .A(n32), .B(n74), .Z(n57) );
  XNOR U814 ( .A(n66), .B(n75), .Z(n74) );
  NANDN U815 ( .A(n76), .B(n77), .Z(n75) );
  OR U816 ( .A(n78), .B(n79), .Z(n66) );
  XOR U817 ( .A(n80), .B(n70), .Z(n32) );
  NANDN U818 ( .A(n81), .B(n82), .Z(n70) );
  ANDN U819 ( .B(n83), .A(n84), .Z(n80) );
  XOR U820 ( .A(key[1241]), .B(n59), .Z(n64) );
  XOR U821 ( .A(n85), .B(n86), .Z(n59) );
  XNOR U822 ( .A(n87), .B(n88), .Z(n86) );
  NANDN U823 ( .A(n89), .B(n42), .Z(n88) );
  XNOR U824 ( .A(n30), .B(n90), .Z(out[88]) );
  XOR U825 ( .A(key[1240]), .B(n60), .Z(n90) );
  XNOR U826 ( .A(n85), .B(n91), .Z(n60) );
  XOR U827 ( .A(n92), .B(n34), .Z(n91) );
  OR U828 ( .A(n93), .B(n78), .Z(n34) );
  XNOR U829 ( .A(n37), .B(n77), .Z(n78) );
  ANDN U830 ( .B(n77), .A(n94), .Z(n92) );
  IV U831 ( .A(n46), .Z(n30) );
  XOR U832 ( .A(n38), .B(n95), .Z(n46) );
  XOR U833 ( .A(n96), .B(n87), .Z(n95) );
  XNOR U834 ( .A(n56), .B(n42), .Z(n53) );
  NOR U835 ( .A(n98), .B(n56), .Z(n96) );
  XNOR U836 ( .A(n85), .B(n99), .Z(n38) );
  XNOR U837 ( .A(n100), .B(n101), .Z(n99) );
  NANDN U838 ( .A(n72), .B(n102), .Z(n101) );
  XOR U839 ( .A(n103), .B(n100), .Z(n85) );
  OR U840 ( .A(n81), .B(n104), .Z(n100) );
  XOR U841 ( .A(n105), .B(n72), .Z(n81) );
  XNOR U842 ( .A(n77), .B(n42), .Z(n72) );
  XOR U843 ( .A(n106), .B(n107), .Z(n42) );
  NANDN U844 ( .A(n108), .B(n109), .Z(n107) );
  XOR U845 ( .A(n110), .B(n111), .Z(n77) );
  NANDN U846 ( .A(n108), .B(n112), .Z(n111) );
  ANDN U847 ( .B(n105), .A(n113), .Z(n103) );
  IV U848 ( .A(n84), .Z(n105) );
  XOR U849 ( .A(n56), .B(n37), .Z(n84) );
  XNOR U850 ( .A(n114), .B(n110), .Z(n37) );
  NANDN U851 ( .A(n115), .B(n116), .Z(n110) );
  XOR U852 ( .A(n112), .B(n117), .Z(n116) );
  ANDN U853 ( .B(n117), .A(n118), .Z(n114) );
  XOR U854 ( .A(n119), .B(n106), .Z(n56) );
  NANDN U855 ( .A(n115), .B(n120), .Z(n106) );
  XOR U856 ( .A(n121), .B(n109), .Z(n120) );
  XNOR U857 ( .A(n122), .B(n123), .Z(n108) );
  XOR U858 ( .A(n124), .B(n125), .Z(n123) );
  XNOR U859 ( .A(n126), .B(n127), .Z(n122) );
  XNOR U860 ( .A(n128), .B(n129), .Z(n127) );
  ANDN U861 ( .B(n121), .A(n125), .Z(n128) );
  ANDN U862 ( .B(n121), .A(n118), .Z(n119) );
  XNOR U863 ( .A(n124), .B(n130), .Z(n118) );
  XOR U864 ( .A(n131), .B(n129), .Z(n130) );
  NAND U865 ( .A(n132), .B(n133), .Z(n129) );
  XNOR U866 ( .A(n126), .B(n109), .Z(n133) );
  IV U867 ( .A(n121), .Z(n126) );
  XNOR U868 ( .A(n112), .B(n125), .Z(n132) );
  IV U869 ( .A(n117), .Z(n125) );
  XOR U870 ( .A(n134), .B(n135), .Z(n117) );
  XNOR U871 ( .A(n136), .B(n137), .Z(n135) );
  XNOR U872 ( .A(n138), .B(n139), .Z(n134) );
  NOR U873 ( .A(n55), .B(n98), .Z(n138) );
  AND U874 ( .A(n109), .B(n112), .Z(n131) );
  XNOR U875 ( .A(n109), .B(n112), .Z(n124) );
  XNOR U876 ( .A(n140), .B(n141), .Z(n112) );
  XNOR U877 ( .A(n142), .B(n137), .Z(n141) );
  XOR U878 ( .A(n143), .B(n144), .Z(n140) );
  XNOR U879 ( .A(n145), .B(n139), .Z(n144) );
  OR U880 ( .A(n54), .B(n97), .Z(n139) );
  XNOR U881 ( .A(n98), .B(n89), .Z(n97) );
  XNOR U882 ( .A(n55), .B(n43), .Z(n54) );
  ANDN U883 ( .B(n146), .A(n89), .Z(n145) );
  XNOR U884 ( .A(n147), .B(n148), .Z(n109) );
  XNOR U885 ( .A(n137), .B(n149), .Z(n148) );
  XOR U886 ( .A(n68), .B(n143), .Z(n149) );
  XNOR U887 ( .A(n98), .B(n150), .Z(n137) );
  XOR U888 ( .A(n36), .B(n151), .Z(n147) );
  XNOR U889 ( .A(n152), .B(n153), .Z(n151) );
  ANDN U890 ( .B(n154), .A(n94), .Z(n152) );
  XNOR U891 ( .A(n155), .B(n156), .Z(n121) );
  XNOR U892 ( .A(n142), .B(n157), .Z(n156) );
  XNOR U893 ( .A(n76), .B(n136), .Z(n157) );
  XOR U894 ( .A(n143), .B(n158), .Z(n136) );
  XNOR U895 ( .A(n159), .B(n160), .Z(n158) );
  NAND U896 ( .A(n102), .B(n73), .Z(n160) );
  XNOR U897 ( .A(n161), .B(n159), .Z(n143) );
  NANDN U898 ( .A(n104), .B(n82), .Z(n159) );
  XOR U899 ( .A(n83), .B(n73), .Z(n82) );
  XNOR U900 ( .A(n154), .B(n43), .Z(n73) );
  XOR U901 ( .A(n113), .B(n102), .Z(n104) );
  XNOR U902 ( .A(n94), .B(n162), .Z(n102) );
  ANDN U903 ( .B(n83), .A(n113), .Z(n161) );
  XNOR U904 ( .A(n36), .B(n98), .Z(n113) );
  XOR U905 ( .A(n163), .B(n164), .Z(n98) );
  XNOR U906 ( .A(n165), .B(n166), .Z(n164) );
  XOR U907 ( .A(n162), .B(n146), .Z(n142) );
  IV U908 ( .A(n43), .Z(n146) );
  XOR U909 ( .A(n167), .B(n168), .Z(n43) );
  XNOR U910 ( .A(n169), .B(n166), .Z(n168) );
  IV U911 ( .A(n89), .Z(n162) );
  XOR U912 ( .A(n166), .B(n170), .Z(n89) );
  XNOR U913 ( .A(n171), .B(n172), .Z(n155) );
  XNOR U914 ( .A(n173), .B(n153), .Z(n172) );
  OR U915 ( .A(n79), .B(n93), .Z(n153) );
  XNOR U916 ( .A(n36), .B(n94), .Z(n93) );
  IV U917 ( .A(n171), .Z(n94) );
  XOR U918 ( .A(n68), .B(n154), .Z(n79) );
  IV U919 ( .A(n76), .Z(n154) );
  XOR U920 ( .A(n150), .B(n174), .Z(n76) );
  XNOR U921 ( .A(n169), .B(n163), .Z(n174) );
  XOR U922 ( .A(n175), .B(n176), .Z(n163) );
  XOR U923 ( .A(n177), .B(n178), .Z(n176) );
  XNOR U924 ( .A(n179), .B(n180), .Z(n175) );
  XNOR U925 ( .A(key[1242]), .B(n181), .Z(n180) );
  IV U926 ( .A(n55), .Z(n150) );
  XOR U927 ( .A(n167), .B(n182), .Z(n55) );
  XOR U928 ( .A(n166), .B(n183), .Z(n182) );
  NOR U929 ( .A(n68), .B(n36), .Z(n173) );
  XOR U930 ( .A(n167), .B(n184), .Z(n68) );
  XOR U931 ( .A(n166), .B(n185), .Z(n184) );
  XOR U932 ( .A(n186), .B(n187), .Z(n166) );
  XOR U933 ( .A(n188), .B(n189), .Z(n187) );
  XOR U934 ( .A(n36), .B(n190), .Z(n186) );
  XNOR U935 ( .A(key[1246]), .B(n191), .Z(n190) );
  IV U936 ( .A(n170), .Z(n167) );
  XOR U937 ( .A(n192), .B(n193), .Z(n170) );
  XOR U938 ( .A(n194), .B(n195), .Z(n193) );
  XNOR U939 ( .A(n196), .B(n197), .Z(n192) );
  XNOR U940 ( .A(key[1245]), .B(n198), .Z(n197) );
  XOR U941 ( .A(n199), .B(n200), .Z(n171) );
  XNOR U942 ( .A(n185), .B(n183), .Z(n200) );
  XNOR U943 ( .A(n201), .B(n202), .Z(n183) );
  XNOR U944 ( .A(n203), .B(n204), .Z(n202) );
  XOR U945 ( .A(key[1247]), .B(n205), .Z(n201) );
  XNOR U946 ( .A(n206), .B(n207), .Z(n185) );
  XOR U947 ( .A(n208), .B(n209), .Z(n207) );
  XNOR U948 ( .A(n210), .B(n211), .Z(n206) );
  XNOR U949 ( .A(key[1244]), .B(n212), .Z(n211) );
  XNOR U950 ( .A(n36), .B(n165), .Z(n199) );
  XOR U951 ( .A(n213), .B(n214), .Z(n165) );
  XNOR U952 ( .A(n215), .B(n216), .Z(n214) );
  XOR U953 ( .A(n169), .B(n217), .Z(n216) );
  XOR U954 ( .A(n218), .B(n219), .Z(n169) );
  XNOR U955 ( .A(n220), .B(n221), .Z(n219) );
  XOR U956 ( .A(n222), .B(n223), .Z(n218) );
  XNOR U957 ( .A(key[1241]), .B(n224), .Z(n223) );
  XNOR U958 ( .A(n225), .B(n226), .Z(n213) );
  XNOR U959 ( .A(key[1243]), .B(n227), .Z(n226) );
  XNOR U960 ( .A(n228), .B(n229), .Z(n36) );
  XOR U961 ( .A(n230), .B(n231), .Z(n229) );
  XOR U962 ( .A(n232), .B(n233), .Z(n228) );
  XNOR U963 ( .A(key[1240]), .B(n234), .Z(n233) );
  XOR U964 ( .A(n235), .B(n236), .Z(out[87]) );
  XOR U965 ( .A(n237), .B(n238), .Z(n235) );
  XNOR U966 ( .A(key[1239]), .B(n239), .Z(n238) );
  XNOR U967 ( .A(n240), .B(n241), .Z(out[86]) );
  XNOR U968 ( .A(key[1238]), .B(n242), .Z(n241) );
  XOR U969 ( .A(n243), .B(n244), .Z(out[85]) );
  XNOR U970 ( .A(n245), .B(n246), .Z(n244) );
  XOR U971 ( .A(n237), .B(n247), .Z(n246) );
  XNOR U972 ( .A(n249), .B(n250), .Z(n248) );
  NANDN U973 ( .A(n251), .B(n252), .Z(n250) );
  XOR U974 ( .A(n254), .B(n255), .Z(n243) );
  XOR U975 ( .A(key[1237]), .B(n256), .Z(n255) );
  ANDN U976 ( .B(n257), .A(n258), .Z(n254) );
  XNOR U977 ( .A(n259), .B(n260), .Z(out[84]) );
  XNOR U978 ( .A(key[1236]), .B(n261), .Z(n260) );
  XOR U979 ( .A(n262), .B(n263), .Z(out[83]) );
  XNOR U980 ( .A(n264), .B(n240), .Z(n263) );
  XNOR U981 ( .A(n265), .B(n266), .Z(n240) );
  XNOR U982 ( .A(n267), .B(n256), .Z(n266) );
  ANDN U983 ( .B(n268), .A(n269), .Z(n256) );
  NOR U984 ( .A(n270), .B(n271), .Z(n267) );
  XNOR U985 ( .A(n272), .B(n273), .Z(n262) );
  XOR U986 ( .A(key[1235]), .B(n274), .Z(n273) );
  XOR U987 ( .A(key[1234]), .B(n259), .Z(out[82]) );
  XNOR U988 ( .A(n239), .B(n275), .Z(n259) );
  IV U989 ( .A(n274), .Z(n239) );
  XOR U990 ( .A(n276), .B(n236), .Z(out[81]) );
  XNOR U991 ( .A(n265), .B(n277), .Z(n264) );
  XNOR U992 ( .A(n278), .B(n279), .Z(n277) );
  NANDN U993 ( .A(n280), .B(n252), .Z(n279) );
  XNOR U994 ( .A(n247), .B(n281), .Z(n265) );
  XNOR U995 ( .A(n282), .B(n283), .Z(n281) );
  NANDN U996 ( .A(n284), .B(n285), .Z(n283) );
  XOR U997 ( .A(n275), .B(n272), .Z(n242) );
  XNOR U998 ( .A(n247), .B(n286), .Z(n272) );
  XNOR U999 ( .A(n278), .B(n287), .Z(n286) );
  NANDN U1000 ( .A(n288), .B(n289), .Z(n287) );
  OR U1001 ( .A(n290), .B(n291), .Z(n278) );
  XOR U1002 ( .A(n292), .B(n282), .Z(n247) );
  NANDN U1003 ( .A(n293), .B(n294), .Z(n282) );
  ANDN U1004 ( .B(n295), .A(n296), .Z(n292) );
  XOR U1005 ( .A(key[1233]), .B(n274), .Z(n276) );
  XOR U1006 ( .A(n297), .B(n298), .Z(n274) );
  XNOR U1007 ( .A(n299), .B(n300), .Z(n298) );
  NANDN U1008 ( .A(n301), .B(n257), .Z(n300) );
  XNOR U1009 ( .A(n245), .B(n302), .Z(out[80]) );
  XOR U1010 ( .A(key[1232]), .B(n275), .Z(n302) );
  XNOR U1011 ( .A(n297), .B(n303), .Z(n275) );
  XOR U1012 ( .A(n304), .B(n249), .Z(n303) );
  OR U1013 ( .A(n305), .B(n290), .Z(n249) );
  XNOR U1014 ( .A(n252), .B(n289), .Z(n290) );
  ANDN U1015 ( .B(n289), .A(n306), .Z(n304) );
  IV U1016 ( .A(n261), .Z(n245) );
  XOR U1017 ( .A(n253), .B(n307), .Z(n261) );
  XOR U1018 ( .A(n308), .B(n299), .Z(n307) );
  XNOR U1019 ( .A(n271), .B(n257), .Z(n268) );
  NOR U1020 ( .A(n310), .B(n271), .Z(n308) );
  XNOR U1021 ( .A(n297), .B(n311), .Z(n253) );
  XNOR U1022 ( .A(n312), .B(n313), .Z(n311) );
  NANDN U1023 ( .A(n284), .B(n314), .Z(n313) );
  XOR U1024 ( .A(n315), .B(n312), .Z(n297) );
  OR U1025 ( .A(n293), .B(n316), .Z(n312) );
  XOR U1026 ( .A(n317), .B(n284), .Z(n293) );
  XNOR U1027 ( .A(n289), .B(n257), .Z(n284) );
  XOR U1028 ( .A(n318), .B(n319), .Z(n257) );
  NANDN U1029 ( .A(n320), .B(n321), .Z(n319) );
  XOR U1030 ( .A(n322), .B(n323), .Z(n289) );
  NANDN U1031 ( .A(n320), .B(n324), .Z(n323) );
  ANDN U1032 ( .B(n317), .A(n325), .Z(n315) );
  IV U1033 ( .A(n296), .Z(n317) );
  XOR U1034 ( .A(n271), .B(n252), .Z(n296) );
  XNOR U1035 ( .A(n326), .B(n322), .Z(n252) );
  NANDN U1036 ( .A(n327), .B(n328), .Z(n322) );
  XOR U1037 ( .A(n324), .B(n329), .Z(n328) );
  ANDN U1038 ( .B(n329), .A(n330), .Z(n326) );
  XOR U1039 ( .A(n331), .B(n318), .Z(n271) );
  NANDN U1040 ( .A(n327), .B(n332), .Z(n318) );
  XOR U1041 ( .A(n333), .B(n321), .Z(n332) );
  XNOR U1042 ( .A(n334), .B(n335), .Z(n320) );
  XOR U1043 ( .A(n336), .B(n337), .Z(n335) );
  XNOR U1044 ( .A(n338), .B(n339), .Z(n334) );
  XNOR U1045 ( .A(n340), .B(n341), .Z(n339) );
  ANDN U1046 ( .B(n333), .A(n337), .Z(n340) );
  ANDN U1047 ( .B(n333), .A(n330), .Z(n331) );
  XNOR U1048 ( .A(n336), .B(n342), .Z(n330) );
  XOR U1049 ( .A(n343), .B(n341), .Z(n342) );
  NAND U1050 ( .A(n344), .B(n345), .Z(n341) );
  XNOR U1051 ( .A(n338), .B(n321), .Z(n345) );
  IV U1052 ( .A(n333), .Z(n338) );
  XNOR U1053 ( .A(n324), .B(n337), .Z(n344) );
  IV U1054 ( .A(n329), .Z(n337) );
  XOR U1055 ( .A(n346), .B(n347), .Z(n329) );
  XNOR U1056 ( .A(n348), .B(n349), .Z(n347) );
  XNOR U1057 ( .A(n350), .B(n351), .Z(n346) );
  NOR U1058 ( .A(n270), .B(n310), .Z(n350) );
  AND U1059 ( .A(n321), .B(n324), .Z(n343) );
  XNOR U1060 ( .A(n321), .B(n324), .Z(n336) );
  XNOR U1061 ( .A(n352), .B(n353), .Z(n324) );
  XNOR U1062 ( .A(n354), .B(n349), .Z(n353) );
  XOR U1063 ( .A(n355), .B(n356), .Z(n352) );
  XNOR U1064 ( .A(n357), .B(n351), .Z(n356) );
  OR U1065 ( .A(n269), .B(n309), .Z(n351) );
  XNOR U1066 ( .A(n310), .B(n301), .Z(n309) );
  XNOR U1067 ( .A(n270), .B(n258), .Z(n269) );
  ANDN U1068 ( .B(n358), .A(n301), .Z(n357) );
  XNOR U1069 ( .A(n359), .B(n360), .Z(n321) );
  XNOR U1070 ( .A(n349), .B(n361), .Z(n360) );
  XOR U1071 ( .A(n280), .B(n355), .Z(n361) );
  XNOR U1072 ( .A(n310), .B(n362), .Z(n349) );
  XOR U1073 ( .A(n251), .B(n363), .Z(n359) );
  XNOR U1074 ( .A(n364), .B(n365), .Z(n363) );
  ANDN U1075 ( .B(n366), .A(n306), .Z(n364) );
  XNOR U1076 ( .A(n367), .B(n368), .Z(n333) );
  XNOR U1077 ( .A(n354), .B(n369), .Z(n368) );
  XNOR U1078 ( .A(n288), .B(n348), .Z(n369) );
  XOR U1079 ( .A(n355), .B(n370), .Z(n348) );
  XNOR U1080 ( .A(n371), .B(n372), .Z(n370) );
  NAND U1081 ( .A(n314), .B(n285), .Z(n372) );
  XNOR U1082 ( .A(n373), .B(n371), .Z(n355) );
  NANDN U1083 ( .A(n316), .B(n294), .Z(n371) );
  XOR U1084 ( .A(n295), .B(n285), .Z(n294) );
  XNOR U1085 ( .A(n366), .B(n258), .Z(n285) );
  XOR U1086 ( .A(n325), .B(n314), .Z(n316) );
  XNOR U1087 ( .A(n306), .B(n374), .Z(n314) );
  ANDN U1088 ( .B(n295), .A(n325), .Z(n373) );
  XNOR U1089 ( .A(n251), .B(n310), .Z(n325) );
  XOR U1090 ( .A(n375), .B(n376), .Z(n310) );
  XNOR U1091 ( .A(n377), .B(n378), .Z(n376) );
  XOR U1092 ( .A(n374), .B(n358), .Z(n354) );
  IV U1093 ( .A(n258), .Z(n358) );
  XOR U1094 ( .A(n379), .B(n380), .Z(n258) );
  XNOR U1095 ( .A(n381), .B(n378), .Z(n380) );
  IV U1096 ( .A(n301), .Z(n374) );
  XOR U1097 ( .A(n378), .B(n382), .Z(n301) );
  XNOR U1098 ( .A(n383), .B(n384), .Z(n367) );
  XNOR U1099 ( .A(n385), .B(n365), .Z(n384) );
  OR U1100 ( .A(n291), .B(n305), .Z(n365) );
  XNOR U1101 ( .A(n251), .B(n306), .Z(n305) );
  IV U1102 ( .A(n383), .Z(n306) );
  XOR U1103 ( .A(n280), .B(n366), .Z(n291) );
  IV U1104 ( .A(n288), .Z(n366) );
  XOR U1105 ( .A(n362), .B(n386), .Z(n288) );
  XNOR U1106 ( .A(n381), .B(n375), .Z(n386) );
  XOR U1107 ( .A(n387), .B(n388), .Z(n375) );
  XNOR U1108 ( .A(n389), .B(n390), .Z(n388) );
  XNOR U1109 ( .A(key[1202]), .B(n391), .Z(n387) );
  IV U1110 ( .A(n270), .Z(n362) );
  XOR U1111 ( .A(n379), .B(n392), .Z(n270) );
  XOR U1112 ( .A(n378), .B(n393), .Z(n392) );
  NOR U1113 ( .A(n280), .B(n251), .Z(n385) );
  XOR U1114 ( .A(n379), .B(n394), .Z(n280) );
  XOR U1115 ( .A(n378), .B(n395), .Z(n394) );
  XOR U1116 ( .A(n396), .B(n397), .Z(n378) );
  XOR U1117 ( .A(n398), .B(n399), .Z(n397) );
  XNOR U1118 ( .A(n400), .B(n401), .Z(n396) );
  XOR U1119 ( .A(key[1206]), .B(n251), .Z(n401) );
  IV U1120 ( .A(n382), .Z(n379) );
  XOR U1121 ( .A(n402), .B(n403), .Z(n382) );
  XNOR U1122 ( .A(n404), .B(n405), .Z(n403) );
  XNOR U1123 ( .A(key[1205]), .B(n406), .Z(n402) );
  XOR U1124 ( .A(n407), .B(n408), .Z(n383) );
  XNOR U1125 ( .A(n395), .B(n393), .Z(n408) );
  XNOR U1126 ( .A(n409), .B(n410), .Z(n393) );
  XNOR U1127 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U1128 ( .A(key[1207]), .B(n413), .Z(n409) );
  XNOR U1129 ( .A(n414), .B(n415), .Z(n395) );
  XNOR U1130 ( .A(n416), .B(n417), .Z(n415) );
  XNOR U1131 ( .A(n418), .B(n419), .Z(n414) );
  XNOR U1132 ( .A(n251), .B(n377), .Z(n407) );
  XOR U1133 ( .A(n421), .B(n422), .Z(n377) );
  XNOR U1134 ( .A(n423), .B(n424), .Z(n422) );
  XNOR U1135 ( .A(n381), .B(n425), .Z(n424) );
  XOR U1136 ( .A(n426), .B(n427), .Z(n381) );
  XOR U1137 ( .A(n428), .B(n429), .Z(n427) );
  XOR U1138 ( .A(key[1201]), .B(n430), .Z(n426) );
  XNOR U1139 ( .A(n431), .B(n432), .Z(n421) );
  XNOR U1140 ( .A(key[1203]), .B(n433), .Z(n432) );
  XNOR U1141 ( .A(n434), .B(n435), .Z(n251) );
  XOR U1142 ( .A(n436), .B(n437), .Z(n435) );
  XNOR U1143 ( .A(key[1200]), .B(n438), .Z(n434) );
  XOR U1144 ( .A(n439), .B(n440), .Z(out[7]) );
  XOR U1145 ( .A(n441), .B(n442), .Z(n439) );
  XNOR U1146 ( .A(key[1159]), .B(n443), .Z(n442) );
  XOR U1147 ( .A(n444), .B(n445), .Z(out[79]) );
  XOR U1148 ( .A(n446), .B(n447), .Z(n444) );
  XNOR U1149 ( .A(key[1231]), .B(n448), .Z(n447) );
  XOR U1150 ( .A(n449), .B(n450), .Z(out[78]) );
  XNOR U1151 ( .A(n451), .B(n452), .Z(n450) );
  XNOR U1152 ( .A(key[1230]), .B(n453), .Z(n449) );
  XOR U1153 ( .A(n454), .B(n455), .Z(out[77]) );
  XNOR U1154 ( .A(n456), .B(n457), .Z(n455) );
  XOR U1155 ( .A(n446), .B(n458), .Z(n457) );
  XNOR U1156 ( .A(n460), .B(n461), .Z(n459) );
  OR U1157 ( .A(n462), .B(n463), .Z(n461) );
  XOR U1158 ( .A(n465), .B(n466), .Z(n454) );
  XOR U1159 ( .A(key[1229]), .B(n467), .Z(n466) );
  ANDN U1160 ( .B(n468), .A(n469), .Z(n465) );
  XNOR U1161 ( .A(n470), .B(n471), .Z(out[76]) );
  XNOR U1162 ( .A(key[1228]), .B(n472), .Z(n471) );
  XOR U1163 ( .A(n473), .B(n474), .Z(out[75]) );
  XNOR U1164 ( .A(n475), .B(n452), .Z(n474) );
  XNOR U1165 ( .A(n476), .B(n477), .Z(n452) );
  XNOR U1166 ( .A(n478), .B(n467), .Z(n477) );
  NOR U1167 ( .A(n479), .B(n480), .Z(n467) );
  NOR U1168 ( .A(n481), .B(n482), .Z(n478) );
  XOR U1169 ( .A(n483), .B(n484), .Z(n473) );
  XOR U1170 ( .A(key[1227]), .B(n485), .Z(n484) );
  XOR U1171 ( .A(key[1226]), .B(n470), .Z(out[74]) );
  XNOR U1172 ( .A(n448), .B(n453), .Z(n470) );
  IV U1173 ( .A(n485), .Z(n448) );
  XOR U1174 ( .A(n486), .B(n445), .Z(out[73]) );
  XNOR U1175 ( .A(n476), .B(n488), .Z(n475) );
  XOR U1176 ( .A(n489), .B(n490), .Z(n488) );
  NOR U1177 ( .A(n491), .B(n462), .Z(n489) );
  XNOR U1178 ( .A(n458), .B(n492), .Z(n476) );
  XNOR U1179 ( .A(n493), .B(n494), .Z(n492) );
  NAND U1180 ( .A(n495), .B(n496), .Z(n494) );
  XOR U1181 ( .A(n453), .B(n483), .Z(n487) );
  IV U1182 ( .A(n451), .Z(n483) );
  XNOR U1183 ( .A(n458), .B(n497), .Z(n451) );
  XNOR U1184 ( .A(n490), .B(n498), .Z(n497) );
  NANDN U1185 ( .A(n499), .B(n500), .Z(n498) );
  OR U1186 ( .A(n501), .B(n502), .Z(n490) );
  XOR U1187 ( .A(n503), .B(n493), .Z(n458) );
  NANDN U1188 ( .A(n504), .B(n505), .Z(n493) );
  AND U1189 ( .A(n506), .B(n507), .Z(n503) );
  XOR U1190 ( .A(key[1225]), .B(n485), .Z(n486) );
  XOR U1191 ( .A(n508), .B(n509), .Z(n485) );
  XNOR U1192 ( .A(n510), .B(n511), .Z(n509) );
  NANDN U1193 ( .A(n469), .B(n512), .Z(n511) );
  XNOR U1194 ( .A(n456), .B(n513), .Z(out[72]) );
  XOR U1195 ( .A(key[1224]), .B(n453), .Z(n513) );
  XNOR U1196 ( .A(n508), .B(n514), .Z(n453) );
  XOR U1197 ( .A(n515), .B(n460), .Z(n514) );
  OR U1198 ( .A(n516), .B(n501), .Z(n460) );
  XNOR U1199 ( .A(n462), .B(n499), .Z(n501) );
  NOR U1200 ( .A(n517), .B(n499), .Z(n515) );
  IV U1201 ( .A(n472), .Z(n456) );
  XOR U1202 ( .A(n464), .B(n518), .Z(n472) );
  XNOR U1203 ( .A(n510), .B(n519), .Z(n518) );
  OR U1204 ( .A(n482), .B(n520), .Z(n519) );
  OR U1205 ( .A(n521), .B(n479), .Z(n510) );
  XOR U1206 ( .A(n482), .B(n522), .Z(n479) );
  XNOR U1207 ( .A(n508), .B(n523), .Z(n464) );
  XNOR U1208 ( .A(n524), .B(n525), .Z(n523) );
  NAND U1209 ( .A(n496), .B(n526), .Z(n525) );
  XOR U1210 ( .A(n527), .B(n524), .Z(n508) );
  OR U1211 ( .A(n504), .B(n528), .Z(n524) );
  XNOR U1212 ( .A(n506), .B(n496), .Z(n504) );
  XOR U1213 ( .A(n499), .B(n469), .Z(n496) );
  IV U1214 ( .A(n522), .Z(n469) );
  XOR U1215 ( .A(n529), .B(n530), .Z(n522) );
  NANDN U1216 ( .A(n531), .B(n532), .Z(n530) );
  XNOR U1217 ( .A(n533), .B(n534), .Z(n499) );
  OR U1218 ( .A(n531), .B(n535), .Z(n534) );
  ANDN U1219 ( .B(n506), .A(n536), .Z(n527) );
  XOR U1220 ( .A(n462), .B(n482), .Z(n506) );
  XNOR U1221 ( .A(n529), .B(n537), .Z(n482) );
  NANDN U1222 ( .A(n538), .B(n539), .Z(n537) );
  NANDN U1223 ( .A(n540), .B(n541), .Z(n529) );
  OR U1224 ( .A(n543), .B(n540), .Z(n533) );
  XOR U1225 ( .A(n544), .B(n531), .Z(n540) );
  XNOR U1226 ( .A(n545), .B(n546), .Z(n531) );
  XOR U1227 ( .A(n547), .B(n539), .Z(n546) );
  XNOR U1228 ( .A(n548), .B(n549), .Z(n545) );
  XNOR U1229 ( .A(n550), .B(n551), .Z(n549) );
  ANDN U1230 ( .B(n539), .A(n552), .Z(n550) );
  IV U1231 ( .A(n553), .Z(n539) );
  ANDN U1232 ( .B(n544), .A(n552), .Z(n542) );
  IV U1233 ( .A(n538), .Z(n544) );
  XNOR U1234 ( .A(n547), .B(n554), .Z(n538) );
  XNOR U1235 ( .A(n551), .B(n555), .Z(n554) );
  NANDN U1236 ( .A(n535), .B(n532), .Z(n555) );
  NANDN U1237 ( .A(n543), .B(n541), .Z(n551) );
  XNOR U1238 ( .A(n532), .B(n553), .Z(n541) );
  XOR U1239 ( .A(n556), .B(n557), .Z(n553) );
  XOR U1240 ( .A(n558), .B(n559), .Z(n557) );
  XNOR U1241 ( .A(n500), .B(n560), .Z(n559) );
  XNOR U1242 ( .A(n561), .B(n562), .Z(n556) );
  XNOR U1243 ( .A(n563), .B(n564), .Z(n562) );
  ANDN U1244 ( .B(n565), .A(n463), .Z(n563) );
  XNOR U1245 ( .A(n552), .B(n535), .Z(n543) );
  IV U1246 ( .A(n548), .Z(n552) );
  XOR U1247 ( .A(n566), .B(n567), .Z(n548) );
  XNOR U1248 ( .A(n568), .B(n560), .Z(n567) );
  XOR U1249 ( .A(n569), .B(n570), .Z(n560) );
  XNOR U1250 ( .A(n571), .B(n572), .Z(n570) );
  NAND U1251 ( .A(n526), .B(n495), .Z(n572) );
  XNOR U1252 ( .A(n573), .B(n574), .Z(n566) );
  ANDN U1253 ( .B(n575), .A(n520), .Z(n573) );
  XOR U1254 ( .A(n535), .B(n532), .Z(n547) );
  XNOR U1255 ( .A(n576), .B(n577), .Z(n532) );
  XNOR U1256 ( .A(n569), .B(n578), .Z(n577) );
  XOR U1257 ( .A(n568), .B(n491), .Z(n578) );
  XOR U1258 ( .A(n463), .B(n579), .Z(n576) );
  XNOR U1259 ( .A(n580), .B(n564), .Z(n579) );
  OR U1260 ( .A(n502), .B(n516), .Z(n564) );
  XNOR U1261 ( .A(n463), .B(n517), .Z(n516) );
  XOR U1262 ( .A(n491), .B(n500), .Z(n502) );
  ANDN U1263 ( .B(n500), .A(n517), .Z(n580) );
  XOR U1264 ( .A(n581), .B(n582), .Z(n535) );
  XOR U1265 ( .A(n569), .B(n558), .Z(n582) );
  XNOR U1266 ( .A(n512), .B(n468), .Z(n558) );
  XOR U1267 ( .A(n583), .B(n571), .Z(n569) );
  NANDN U1268 ( .A(n528), .B(n505), .Z(n571) );
  XOR U1269 ( .A(n507), .B(n495), .Z(n505) );
  XOR U1270 ( .A(n468), .B(n500), .Z(n495) );
  XNOR U1271 ( .A(n575), .B(n584), .Z(n500) );
  XOR U1272 ( .A(n585), .B(n586), .Z(n584) );
  XOR U1273 ( .A(n536), .B(n526), .Z(n528) );
  XNOR U1274 ( .A(n517), .B(n512), .Z(n526) );
  IV U1275 ( .A(n561), .Z(n517) );
  XOR U1276 ( .A(n587), .B(n588), .Z(n561) );
  XOR U1277 ( .A(n589), .B(n590), .Z(n588) );
  XNOR U1278 ( .A(n463), .B(n591), .Z(n587) );
  ANDN U1279 ( .B(n507), .A(n536), .Z(n583) );
  XNOR U1280 ( .A(n463), .B(n520), .Z(n536) );
  XOR U1281 ( .A(n575), .B(n565), .Z(n507) );
  IV U1282 ( .A(n491), .Z(n565) );
  XOR U1283 ( .A(n592), .B(n593), .Z(n491) );
  XOR U1284 ( .A(n594), .B(n590), .Z(n593) );
  XNOR U1285 ( .A(n595), .B(n596), .Z(n590) );
  XNOR U1286 ( .A(n597), .B(n598), .Z(n596) );
  XNOR U1287 ( .A(key[1164]), .B(n599), .Z(n595) );
  XOR U1288 ( .A(n568), .B(n600), .Z(n581) );
  XNOR U1289 ( .A(n601), .B(n574), .Z(n600) );
  OR U1290 ( .A(n480), .B(n521), .Z(n574) );
  XNOR U1291 ( .A(n602), .B(n512), .Z(n521) );
  XNOR U1292 ( .A(n575), .B(n468), .Z(n480) );
  IV U1293 ( .A(n481), .Z(n575) );
  AND U1294 ( .A(n468), .B(n512), .Z(n601) );
  XOR U1295 ( .A(n594), .B(n592), .Z(n512) );
  XNOR U1296 ( .A(n592), .B(n603), .Z(n468) );
  XNOR U1297 ( .A(n520), .B(n481), .Z(n568) );
  XOR U1298 ( .A(n592), .B(n604), .Z(n481) );
  XNOR U1299 ( .A(n594), .B(n589), .Z(n604) );
  XOR U1300 ( .A(n605), .B(n606), .Z(n589) );
  XNOR U1301 ( .A(n607), .B(n608), .Z(n606) );
  XNOR U1302 ( .A(key[1167]), .B(n609), .Z(n605) );
  XNOR U1303 ( .A(n610), .B(n611), .Z(n592) );
  XOR U1304 ( .A(n612), .B(n613), .Z(n611) );
  XNOR U1305 ( .A(n614), .B(n615), .Z(n610) );
  XNOR U1306 ( .A(key[1165]), .B(n616), .Z(n615) );
  IV U1307 ( .A(n602), .Z(n520) );
  XNOR U1308 ( .A(n586), .B(n617), .Z(n602) );
  XOR U1309 ( .A(n618), .B(n619), .Z(n594) );
  XNOR U1310 ( .A(n463), .B(n620), .Z(n619) );
  XNOR U1311 ( .A(n621), .B(n622), .Z(n463) );
  XNOR U1312 ( .A(n623), .B(n624), .Z(n622) );
  XNOR U1313 ( .A(n625), .B(n626), .Z(n621) );
  XOR U1314 ( .A(key[1160]), .B(n627), .Z(n626) );
  XNOR U1315 ( .A(n628), .B(n629), .Z(n618) );
  XNOR U1316 ( .A(key[1166]), .B(n630), .Z(n629) );
  XOR U1317 ( .A(n631), .B(n632), .Z(n591) );
  XNOR U1318 ( .A(n633), .B(n634), .Z(n632) );
  XOR U1319 ( .A(n635), .B(n585), .Z(n634) );
  XNOR U1320 ( .A(n636), .B(n637), .Z(n585) );
  XNOR U1321 ( .A(n638), .B(n639), .Z(n637) );
  XNOR U1322 ( .A(n640), .B(n641), .Z(n636) );
  XNOR U1323 ( .A(key[1161]), .B(n642), .Z(n641) );
  XNOR U1324 ( .A(n643), .B(n644), .Z(n631) );
  XOR U1325 ( .A(key[1163]), .B(n645), .Z(n644) );
  XOR U1326 ( .A(n646), .B(n647), .Z(n586) );
  XOR U1327 ( .A(n648), .B(n649), .Z(n647) );
  XOR U1328 ( .A(n650), .B(n651), .Z(n646) );
  XNOR U1329 ( .A(key[1162]), .B(n652), .Z(n651) );
  XOR U1330 ( .A(n653), .B(n654), .Z(out[71]) );
  XNOR U1331 ( .A(n655), .B(n656), .Z(n653) );
  XNOR U1332 ( .A(key[1223]), .B(n657), .Z(n656) );
  XOR U1333 ( .A(n658), .B(n659), .Z(out[70]) );
  XNOR U1334 ( .A(n660), .B(n661), .Z(n659) );
  XNOR U1335 ( .A(key[1222]), .B(n662), .Z(n658) );
  XNOR U1336 ( .A(n663), .B(n664), .Z(out[6]) );
  XNOR U1337 ( .A(key[1158]), .B(n665), .Z(n664) );
  XOR U1338 ( .A(n666), .B(n667), .Z(out[69]) );
  XNOR U1339 ( .A(n668), .B(n669), .Z(n667) );
  XNOR U1340 ( .A(n657), .B(n670), .Z(n669) );
  XNOR U1341 ( .A(n671), .B(n672), .Z(n657) );
  XNOR U1342 ( .A(n673), .B(n674), .Z(n672) );
  OR U1343 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U1344 ( .A(n677), .B(n678), .Z(n666) );
  XOR U1345 ( .A(key[1221]), .B(n679), .Z(n678) );
  ANDN U1346 ( .B(n680), .A(n681), .Z(n679) );
  XNOR U1347 ( .A(n682), .B(n683), .Z(out[68]) );
  XNOR U1348 ( .A(key[1220]), .B(n684), .Z(n683) );
  XOR U1349 ( .A(n685), .B(n686), .Z(out[67]) );
  XNOR U1350 ( .A(n687), .B(n661), .Z(n686) );
  XNOR U1351 ( .A(n688), .B(n689), .Z(n661) );
  XNOR U1352 ( .A(n677), .B(n690), .Z(n689) );
  OR U1353 ( .A(n691), .B(n692), .Z(n690) );
  NANDN U1354 ( .A(n693), .B(n694), .Z(n677) );
  XNOR U1355 ( .A(n695), .B(n696), .Z(n685) );
  XNOR U1356 ( .A(key[1219]), .B(n660), .Z(n696) );
  XOR U1357 ( .A(key[1218]), .B(n682), .Z(out[66]) );
  XNOR U1358 ( .A(n662), .B(n687), .Z(n682) );
  XOR U1359 ( .A(n697), .B(n654), .Z(out[65]) );
  XNOR U1360 ( .A(n695), .B(n687), .Z(n654) );
  XNOR U1361 ( .A(n698), .B(n699), .Z(n687) );
  XNOR U1362 ( .A(n700), .B(n701), .Z(n699) );
  NAND U1363 ( .A(n702), .B(n680), .Z(n701) );
  XNOR U1364 ( .A(n688), .B(n703), .Z(n695) );
  XNOR U1365 ( .A(n704), .B(n705), .Z(n703) );
  OR U1366 ( .A(n675), .B(n706), .Z(n705) );
  XNOR U1367 ( .A(n670), .B(n707), .Z(n688) );
  XNOR U1368 ( .A(n708), .B(n709), .Z(n707) );
  NANDN U1369 ( .A(n710), .B(n711), .Z(n709) );
  XNOR U1370 ( .A(key[1217]), .B(n655), .Z(n697) );
  XOR U1371 ( .A(n712), .B(n660), .Z(n655) );
  XNOR U1372 ( .A(n670), .B(n713), .Z(n660) );
  XOR U1373 ( .A(n714), .B(n704), .Z(n713) );
  OR U1374 ( .A(n715), .B(n716), .Z(n704) );
  AND U1375 ( .A(n717), .B(n718), .Z(n714) );
  XOR U1376 ( .A(n719), .B(n708), .Z(n670) );
  NANDN U1377 ( .A(n720), .B(n721), .Z(n708) );
  AND U1378 ( .A(n722), .B(n723), .Z(n719) );
  XNOR U1379 ( .A(n668), .B(n724), .Z(out[64]) );
  XNOR U1380 ( .A(key[1216]), .B(n712), .Z(n724) );
  IV U1381 ( .A(n662), .Z(n712) );
  XNOR U1382 ( .A(n698), .B(n725), .Z(n662) );
  XOR U1383 ( .A(n726), .B(n673), .Z(n725) );
  OR U1384 ( .A(n727), .B(n715), .Z(n673) );
  XOR U1385 ( .A(n675), .B(n718), .Z(n715) );
  ANDN U1386 ( .B(n718), .A(n728), .Z(n726) );
  IV U1387 ( .A(n684), .Z(n668) );
  XOR U1388 ( .A(n671), .B(n729), .Z(n684) );
  XOR U1389 ( .A(n730), .B(n700), .Z(n729) );
  NANDN U1390 ( .A(n731), .B(n694), .Z(n700) );
  XNOR U1391 ( .A(n691), .B(n680), .Z(n694) );
  NOR U1392 ( .A(n732), .B(n691), .Z(n730) );
  XNOR U1393 ( .A(n698), .B(n733), .Z(n671) );
  XNOR U1394 ( .A(n734), .B(n735), .Z(n733) );
  NANDN U1395 ( .A(n710), .B(n736), .Z(n735) );
  XOR U1396 ( .A(n737), .B(n734), .Z(n698) );
  OR U1397 ( .A(n720), .B(n738), .Z(n734) );
  XOR U1398 ( .A(n722), .B(n710), .Z(n720) );
  XNOR U1399 ( .A(n718), .B(n680), .Z(n710) );
  XOR U1400 ( .A(n739), .B(n740), .Z(n680) );
  NANDN U1401 ( .A(n741), .B(n742), .Z(n740) );
  XOR U1402 ( .A(n743), .B(n744), .Z(n718) );
  OR U1403 ( .A(n741), .B(n745), .Z(n744) );
  ANDN U1404 ( .B(n722), .A(n746), .Z(n737) );
  XOR U1405 ( .A(n675), .B(n691), .Z(n722) );
  XOR U1406 ( .A(n747), .B(n739), .Z(n691) );
  NANDN U1407 ( .A(n748), .B(n749), .Z(n739) );
  ANDN U1408 ( .B(n750), .A(n751), .Z(n747) );
  NANDN U1409 ( .A(n748), .B(n753), .Z(n743) );
  XOR U1410 ( .A(n754), .B(n741), .Z(n748) );
  XNOR U1411 ( .A(n755), .B(n756), .Z(n741) );
  XOR U1412 ( .A(n757), .B(n750), .Z(n756) );
  XNOR U1413 ( .A(n758), .B(n759), .Z(n755) );
  XNOR U1414 ( .A(n760), .B(n761), .Z(n759) );
  ANDN U1415 ( .B(n750), .A(n762), .Z(n760) );
  IV U1416 ( .A(n763), .Z(n750) );
  ANDN U1417 ( .B(n754), .A(n762), .Z(n752) );
  IV U1418 ( .A(n758), .Z(n762) );
  IV U1419 ( .A(n751), .Z(n754) );
  XNOR U1420 ( .A(n757), .B(n764), .Z(n751) );
  XOR U1421 ( .A(n765), .B(n761), .Z(n764) );
  NAND U1422 ( .A(n753), .B(n749), .Z(n761) );
  XNOR U1423 ( .A(n742), .B(n763), .Z(n749) );
  XOR U1424 ( .A(n766), .B(n767), .Z(n763) );
  XOR U1425 ( .A(n768), .B(n769), .Z(n767) );
  XNOR U1426 ( .A(n717), .B(n770), .Z(n769) );
  XNOR U1427 ( .A(n771), .B(n772), .Z(n766) );
  XNOR U1428 ( .A(n773), .B(n774), .Z(n772) );
  ANDN U1429 ( .B(n775), .A(n676), .Z(n773) );
  XNOR U1430 ( .A(n758), .B(n745), .Z(n753) );
  XOR U1431 ( .A(n776), .B(n777), .Z(n758) );
  XNOR U1432 ( .A(n778), .B(n770), .Z(n777) );
  XOR U1433 ( .A(n779), .B(n780), .Z(n770) );
  XNOR U1434 ( .A(n781), .B(n782), .Z(n780) );
  NAND U1435 ( .A(n736), .B(n711), .Z(n782) );
  XNOR U1436 ( .A(n783), .B(n784), .Z(n776) );
  ANDN U1437 ( .B(n785), .A(n732), .Z(n783) );
  ANDN U1438 ( .B(n742), .A(n745), .Z(n765) );
  XOR U1439 ( .A(n745), .B(n742), .Z(n757) );
  XNOR U1440 ( .A(n786), .B(n787), .Z(n742) );
  XNOR U1441 ( .A(n779), .B(n788), .Z(n787) );
  XOR U1442 ( .A(n778), .B(n706), .Z(n788) );
  XOR U1443 ( .A(n676), .B(n789), .Z(n786) );
  XNOR U1444 ( .A(n790), .B(n774), .Z(n789) );
  OR U1445 ( .A(n716), .B(n727), .Z(n774) );
  XNOR U1446 ( .A(n676), .B(n728), .Z(n727) );
  XOR U1447 ( .A(n706), .B(n717), .Z(n716) );
  ANDN U1448 ( .B(n717), .A(n728), .Z(n790) );
  XOR U1449 ( .A(n791), .B(n792), .Z(n745) );
  XOR U1450 ( .A(n779), .B(n768), .Z(n792) );
  XOR U1451 ( .A(n702), .B(n681), .Z(n768) );
  XOR U1452 ( .A(n793), .B(n781), .Z(n779) );
  NANDN U1453 ( .A(n738), .B(n721), .Z(n781) );
  XOR U1454 ( .A(n723), .B(n711), .Z(n721) );
  XNOR U1455 ( .A(n785), .B(n794), .Z(n717) );
  XOR U1456 ( .A(n795), .B(n796), .Z(n794) );
  XOR U1457 ( .A(n746), .B(n736), .Z(n738) );
  XNOR U1458 ( .A(n728), .B(n702), .Z(n736) );
  IV U1459 ( .A(n771), .Z(n728) );
  XOR U1460 ( .A(n797), .B(n798), .Z(n771) );
  XOR U1461 ( .A(n799), .B(n800), .Z(n798) );
  XNOR U1462 ( .A(n676), .B(n801), .Z(n797) );
  ANDN U1463 ( .B(n723), .A(n746), .Z(n793) );
  XNOR U1464 ( .A(n676), .B(n732), .Z(n746) );
  XOR U1465 ( .A(n785), .B(n775), .Z(n723) );
  IV U1466 ( .A(n706), .Z(n775) );
  XOR U1467 ( .A(n802), .B(n803), .Z(n706) );
  XOR U1468 ( .A(n804), .B(n800), .Z(n803) );
  XNOR U1469 ( .A(n805), .B(n806), .Z(n800) );
  XNOR U1470 ( .A(n807), .B(n808), .Z(n806) );
  XNOR U1471 ( .A(n809), .B(n810), .Z(n805) );
  XNOR U1472 ( .A(key[1252]), .B(n811), .Z(n810) );
  IV U1473 ( .A(n692), .Z(n785) );
  XOR U1474 ( .A(n778), .B(n812), .Z(n791) );
  XNOR U1475 ( .A(n813), .B(n784), .Z(n812) );
  OR U1476 ( .A(n693), .B(n731), .Z(n784) );
  XNOR U1477 ( .A(n814), .B(n702), .Z(n731) );
  XNOR U1478 ( .A(n692), .B(n681), .Z(n693) );
  ANDN U1479 ( .B(n702), .A(n681), .Z(n813) );
  XOR U1480 ( .A(n802), .B(n815), .Z(n681) );
  XNOR U1481 ( .A(n816), .B(n804), .Z(n815) );
  XOR U1482 ( .A(n804), .B(n802), .Z(n702) );
  XNOR U1483 ( .A(n732), .B(n692), .Z(n778) );
  XOR U1484 ( .A(n802), .B(n817), .Z(n692) );
  XNOR U1485 ( .A(n804), .B(n799), .Z(n817) );
  XOR U1486 ( .A(n818), .B(n819), .Z(n799) );
  XNOR U1487 ( .A(n820), .B(n821), .Z(n819) );
  XOR U1488 ( .A(key[1255]), .B(n822), .Z(n818) );
  XNOR U1489 ( .A(n823), .B(n824), .Z(n802) );
  XNOR U1490 ( .A(n825), .B(n826), .Z(n824) );
  XOR U1491 ( .A(key[1253]), .B(n827), .Z(n823) );
  IV U1492 ( .A(n814), .Z(n732) );
  XNOR U1493 ( .A(n795), .B(n801), .Z(n828) );
  XOR U1494 ( .A(n829), .B(n830), .Z(n801) );
  XOR U1495 ( .A(n831), .B(n832), .Z(n830) );
  XOR U1496 ( .A(n833), .B(n796), .Z(n832) );
  IV U1497 ( .A(n816), .Z(n796) );
  XOR U1498 ( .A(n834), .B(n835), .Z(n816) );
  XNOR U1499 ( .A(n836), .B(n837), .Z(n835) );
  XNOR U1500 ( .A(key[1249]), .B(n838), .Z(n834) );
  XNOR U1501 ( .A(n839), .B(n840), .Z(n829) );
  XNOR U1502 ( .A(key[1251]), .B(n841), .Z(n840) );
  XOR U1503 ( .A(n842), .B(n843), .Z(n795) );
  XOR U1504 ( .A(n844), .B(n845), .Z(n843) );
  XOR U1505 ( .A(key[1250]), .B(n846), .Z(n842) );
  XOR U1506 ( .A(n847), .B(n848), .Z(n804) );
  XNOR U1507 ( .A(n851), .B(n852), .Z(n847) );
  XOR U1508 ( .A(key[1254]), .B(n676), .Z(n852) );
  XNOR U1509 ( .A(n853), .B(n854), .Z(n676) );
  XOR U1510 ( .A(n855), .B(n856), .Z(n854) );
  XNOR U1511 ( .A(key[1248]), .B(n857), .Z(n853) );
  XOR U1512 ( .A(n858), .B(n859), .Z(out[63]) );
  XOR U1513 ( .A(n860), .B(n861), .Z(n858) );
  XNOR U1514 ( .A(key[1215]), .B(n862), .Z(n861) );
  XNOR U1515 ( .A(n863), .B(n864), .Z(out[62]) );
  XNOR U1516 ( .A(key[1214]), .B(n865), .Z(n864) );
  XOR U1517 ( .A(n866), .B(n867), .Z(out[61]) );
  XNOR U1518 ( .A(n868), .B(n869), .Z(n867) );
  XOR U1519 ( .A(n860), .B(n870), .Z(n869) );
  XNOR U1520 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U1521 ( .A(n874), .B(n875), .Z(n873) );
  XOR U1522 ( .A(n877), .B(n878), .Z(n866) );
  XOR U1523 ( .A(key[1213]), .B(n879), .Z(n878) );
  ANDN U1524 ( .B(n880), .A(n881), .Z(n877) );
  XNOR U1525 ( .A(n882), .B(n883), .Z(out[60]) );
  XNOR U1526 ( .A(key[1212]), .B(n884), .Z(n883) );
  XOR U1527 ( .A(n885), .B(n886), .Z(out[5]) );
  XNOR U1528 ( .A(n887), .B(n888), .Z(n886) );
  XOR U1529 ( .A(n441), .B(n889), .Z(n888) );
  XNOR U1530 ( .A(n891), .B(n892), .Z(n890) );
  NANDN U1531 ( .A(n893), .B(n894), .Z(n892) );
  XOR U1532 ( .A(n896), .B(n897), .Z(n885) );
  XOR U1533 ( .A(key[1157]), .B(n898), .Z(n897) );
  ANDN U1534 ( .B(n899), .A(n900), .Z(n896) );
  XOR U1535 ( .A(n901), .B(n902), .Z(out[59]) );
  XNOR U1536 ( .A(n903), .B(n863), .Z(n902) );
  XNOR U1537 ( .A(n904), .B(n905), .Z(n863) );
  XNOR U1538 ( .A(n906), .B(n879), .Z(n905) );
  ANDN U1539 ( .B(n907), .A(n908), .Z(n879) );
  NOR U1540 ( .A(n909), .B(n910), .Z(n906) );
  XNOR U1541 ( .A(n911), .B(n912), .Z(n901) );
  XOR U1542 ( .A(key[1211]), .B(n913), .Z(n912) );
  XOR U1543 ( .A(key[1210]), .B(n882), .Z(out[58]) );
  XNOR U1544 ( .A(n862), .B(n914), .Z(n882) );
  IV U1545 ( .A(n913), .Z(n862) );
  XOR U1546 ( .A(n915), .B(n859), .Z(out[57]) );
  XNOR U1547 ( .A(n904), .B(n916), .Z(n903) );
  XNOR U1548 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U1549 ( .A(n919), .B(n875), .Z(n918) );
  XNOR U1550 ( .A(n870), .B(n920), .Z(n904) );
  XNOR U1551 ( .A(n921), .B(n922), .Z(n920) );
  NANDN U1552 ( .A(n923), .B(n924), .Z(n922) );
  XOR U1553 ( .A(n914), .B(n911), .Z(n865) );
  XNOR U1554 ( .A(n870), .B(n925), .Z(n911) );
  XNOR U1555 ( .A(n917), .B(n926), .Z(n925) );
  NANDN U1556 ( .A(n927), .B(n928), .Z(n926) );
  OR U1557 ( .A(n929), .B(n930), .Z(n917) );
  XOR U1558 ( .A(n931), .B(n921), .Z(n870) );
  NANDN U1559 ( .A(n932), .B(n933), .Z(n921) );
  ANDN U1560 ( .B(n934), .A(n935), .Z(n931) );
  XOR U1561 ( .A(key[1209]), .B(n913), .Z(n915) );
  XOR U1562 ( .A(n936), .B(n937), .Z(n913) );
  XNOR U1563 ( .A(n938), .B(n939), .Z(n937) );
  NANDN U1564 ( .A(n940), .B(n880), .Z(n939) );
  XNOR U1565 ( .A(n868), .B(n941), .Z(out[56]) );
  XOR U1566 ( .A(key[1208]), .B(n914), .Z(n941) );
  XNOR U1567 ( .A(n936), .B(n942), .Z(n914) );
  XOR U1568 ( .A(n943), .B(n872), .Z(n942) );
  OR U1569 ( .A(n944), .B(n929), .Z(n872) );
  XNOR U1570 ( .A(n875), .B(n928), .Z(n929) );
  ANDN U1571 ( .B(n945), .A(n946), .Z(n943) );
  IV U1572 ( .A(n884), .Z(n868) );
  XOR U1573 ( .A(n876), .B(n947), .Z(n884) );
  XOR U1574 ( .A(n948), .B(n938), .Z(n947) );
  XNOR U1575 ( .A(n910), .B(n880), .Z(n907) );
  NOR U1576 ( .A(n950), .B(n910), .Z(n948) );
  XNOR U1577 ( .A(n936), .B(n951), .Z(n876) );
  XNOR U1578 ( .A(n952), .B(n953), .Z(n951) );
  NANDN U1579 ( .A(n923), .B(n954), .Z(n953) );
  XOR U1580 ( .A(n955), .B(n952), .Z(n936) );
  OR U1581 ( .A(n932), .B(n956), .Z(n952) );
  XOR U1582 ( .A(n957), .B(n923), .Z(n932) );
  XNOR U1583 ( .A(n928), .B(n880), .Z(n923) );
  XOR U1584 ( .A(n958), .B(n959), .Z(n880) );
  NANDN U1585 ( .A(n960), .B(n961), .Z(n959) );
  IV U1586 ( .A(n946), .Z(n928) );
  XNOR U1587 ( .A(n962), .B(n963), .Z(n946) );
  NANDN U1588 ( .A(n960), .B(n964), .Z(n963) );
  ANDN U1589 ( .B(n957), .A(n965), .Z(n955) );
  IV U1590 ( .A(n935), .Z(n957) );
  XOR U1591 ( .A(n910), .B(n875), .Z(n935) );
  XNOR U1592 ( .A(n966), .B(n962), .Z(n875) );
  NANDN U1593 ( .A(n967), .B(n968), .Z(n962) );
  XOR U1594 ( .A(n964), .B(n969), .Z(n968) );
  ANDN U1595 ( .B(n969), .A(n970), .Z(n966) );
  XOR U1596 ( .A(n971), .B(n958), .Z(n910) );
  NANDN U1597 ( .A(n967), .B(n972), .Z(n958) );
  XOR U1598 ( .A(n973), .B(n961), .Z(n972) );
  XNOR U1599 ( .A(n974), .B(n975), .Z(n960) );
  XOR U1600 ( .A(n976), .B(n977), .Z(n975) );
  XNOR U1601 ( .A(n978), .B(n979), .Z(n974) );
  XNOR U1602 ( .A(n980), .B(n981), .Z(n979) );
  ANDN U1603 ( .B(n973), .A(n977), .Z(n980) );
  ANDN U1604 ( .B(n973), .A(n970), .Z(n971) );
  XNOR U1605 ( .A(n976), .B(n982), .Z(n970) );
  XOR U1606 ( .A(n983), .B(n981), .Z(n982) );
  NAND U1607 ( .A(n984), .B(n985), .Z(n981) );
  XNOR U1608 ( .A(n978), .B(n961), .Z(n985) );
  IV U1609 ( .A(n973), .Z(n978) );
  XNOR U1610 ( .A(n964), .B(n977), .Z(n984) );
  IV U1611 ( .A(n969), .Z(n977) );
  XOR U1612 ( .A(n986), .B(n987), .Z(n969) );
  XNOR U1613 ( .A(n988), .B(n989), .Z(n987) );
  XNOR U1614 ( .A(n990), .B(n991), .Z(n986) );
  NOR U1615 ( .A(n909), .B(n950), .Z(n990) );
  AND U1616 ( .A(n961), .B(n964), .Z(n983) );
  XNOR U1617 ( .A(n961), .B(n964), .Z(n976) );
  XNOR U1618 ( .A(n992), .B(n993), .Z(n964) );
  XNOR U1619 ( .A(n994), .B(n989), .Z(n993) );
  XOR U1620 ( .A(n995), .B(n996), .Z(n992) );
  XNOR U1621 ( .A(n997), .B(n991), .Z(n996) );
  OR U1622 ( .A(n908), .B(n949), .Z(n991) );
  XNOR U1623 ( .A(n950), .B(n940), .Z(n949) );
  XNOR U1624 ( .A(n909), .B(n881), .Z(n908) );
  ANDN U1625 ( .B(n998), .A(n940), .Z(n997) );
  XNOR U1626 ( .A(n999), .B(n1000), .Z(n961) );
  XNOR U1627 ( .A(n989), .B(n1001), .Z(n1000) );
  XOR U1628 ( .A(n919), .B(n995), .Z(n1001) );
  XNOR U1629 ( .A(n950), .B(n1002), .Z(n989) );
  XNOR U1630 ( .A(n1003), .B(n1004), .Z(n999) );
  XNOR U1631 ( .A(n1005), .B(n1006), .Z(n1004) );
  ANDN U1632 ( .B(n945), .A(n927), .Z(n1005) );
  XNOR U1633 ( .A(n1007), .B(n1008), .Z(n973) );
  XNOR U1634 ( .A(n994), .B(n1009), .Z(n1008) );
  XNOR U1635 ( .A(n927), .B(n988), .Z(n1009) );
  XOR U1636 ( .A(n995), .B(n1010), .Z(n988) );
  XNOR U1637 ( .A(n1011), .B(n1012), .Z(n1010) );
  NAND U1638 ( .A(n954), .B(n924), .Z(n1012) );
  XNOR U1639 ( .A(n1013), .B(n1011), .Z(n995) );
  NANDN U1640 ( .A(n956), .B(n933), .Z(n1011) );
  XOR U1641 ( .A(n934), .B(n924), .Z(n933) );
  XNOR U1642 ( .A(n1014), .B(n881), .Z(n924) );
  XOR U1643 ( .A(n965), .B(n954), .Z(n956) );
  XOR U1644 ( .A(n945), .B(n1015), .Z(n954) );
  ANDN U1645 ( .B(n934), .A(n965), .Z(n1013) );
  XOR U1646 ( .A(n1003), .B(n950), .Z(n965) );
  XOR U1647 ( .A(n1016), .B(n1017), .Z(n950) );
  XNOR U1648 ( .A(n1018), .B(n1019), .Z(n1017) );
  XOR U1649 ( .A(n1020), .B(n1002), .Z(n934) );
  XOR U1650 ( .A(n1015), .B(n998), .Z(n994) );
  IV U1651 ( .A(n881), .Z(n998) );
  XOR U1652 ( .A(n1021), .B(n1022), .Z(n881) );
  XNOR U1653 ( .A(n1023), .B(n1019), .Z(n1022) );
  IV U1654 ( .A(n940), .Z(n1015) );
  XOR U1655 ( .A(n1019), .B(n1024), .Z(n940) );
  XNOR U1656 ( .A(n945), .B(n1025), .Z(n1007) );
  XNOR U1657 ( .A(n1026), .B(n1006), .Z(n1025) );
  OR U1658 ( .A(n930), .B(n944), .Z(n1006) );
  XNOR U1659 ( .A(n1003), .B(n945), .Z(n944) );
  XOR U1660 ( .A(n919), .B(n1014), .Z(n930) );
  IV U1661 ( .A(n927), .Z(n1014) );
  XOR U1662 ( .A(n1002), .B(n1027), .Z(n927) );
  XNOR U1663 ( .A(n1023), .B(n1016), .Z(n1027) );
  XOR U1664 ( .A(n1028), .B(n1029), .Z(n1016) );
  XOR U1665 ( .A(n1030), .B(n1031), .Z(n1029) );
  XOR U1666 ( .A(n429), .B(n1032), .Z(n1028) );
  XNOR U1667 ( .A(key[1210]), .B(n1033), .Z(n1032) );
  IV U1668 ( .A(n909), .Z(n1002) );
  XOR U1669 ( .A(n1021), .B(n1034), .Z(n909) );
  XOR U1670 ( .A(n1019), .B(n1035), .Z(n1034) );
  ANDN U1671 ( .B(n1020), .A(n874), .Z(n1026) );
  IV U1672 ( .A(n919), .Z(n1020) );
  XOR U1673 ( .A(n1021), .B(n1036), .Z(n919) );
  XOR U1674 ( .A(n1019), .B(n1037), .Z(n1036) );
  XOR U1675 ( .A(n1038), .B(n1039), .Z(n1019) );
  XOR U1676 ( .A(n1040), .B(n874), .Z(n1039) );
  IV U1677 ( .A(n1003), .Z(n874) );
  XOR U1678 ( .A(n399), .B(n1041), .Z(n1038) );
  XNOR U1679 ( .A(key[1214]), .B(n1042), .Z(n1041) );
  XNOR U1680 ( .A(n413), .B(n1043), .Z(n399) );
  IV U1681 ( .A(n1024), .Z(n1021) );
  XOR U1682 ( .A(n1044), .B(n1045), .Z(n1024) );
  XOR U1683 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U1684 ( .A(n1048), .B(n1049), .Z(n1044) );
  XNOR U1685 ( .A(key[1213]), .B(n1050), .Z(n1049) );
  XOR U1686 ( .A(n1051), .B(n1052), .Z(n945) );
  XNOR U1687 ( .A(n1037), .B(n1035), .Z(n1052) );
  XNOR U1688 ( .A(n1053), .B(n1054), .Z(n1035) );
  XOR U1689 ( .A(n1055), .B(n1056), .Z(n1054) );
  XNOR U1690 ( .A(key[1215]), .B(n1057), .Z(n1053) );
  XNOR U1691 ( .A(n1058), .B(n1059), .Z(n1037) );
  XNOR U1692 ( .A(n417), .B(n1060), .Z(n1058) );
  XOR U1693 ( .A(key[1212]), .B(n1061), .Z(n1060) );
  XNOR U1694 ( .A(n1062), .B(n1063), .Z(n417) );
  XOR U1695 ( .A(n1003), .B(n1018), .Z(n1051) );
  XOR U1696 ( .A(n1064), .B(n1065), .Z(n1018) );
  XNOR U1697 ( .A(n1023), .B(n1066), .Z(n1065) );
  XOR U1698 ( .A(n1067), .B(n1068), .Z(n1066) );
  XOR U1699 ( .A(n1069), .B(n1070), .Z(n1023) );
  XNOR U1700 ( .A(n1071), .B(n1072), .Z(n1070) );
  XOR U1701 ( .A(n1073), .B(n1074), .Z(n1069) );
  XNOR U1702 ( .A(key[1209]), .B(n436), .Z(n1074) );
  XNOR U1703 ( .A(n423), .B(n1075), .Z(n1064) );
  XNOR U1704 ( .A(key[1211]), .B(n1076), .Z(n1075) );
  XOR U1705 ( .A(n413), .B(n1077), .Z(n423) );
  XOR U1706 ( .A(n1078), .B(n1079), .Z(n1003) );
  XOR U1707 ( .A(n1080), .B(n413), .Z(n1079) );
  XNOR U1708 ( .A(n1081), .B(n1082), .Z(n1078) );
  XNOR U1709 ( .A(key[1208]), .B(n1083), .Z(n1082) );
  XOR U1710 ( .A(n1084), .B(n1085), .Z(out[55]) );
  XOR U1711 ( .A(n1086), .B(n1087), .Z(n1084) );
  XNOR U1712 ( .A(key[1207]), .B(n1088), .Z(n1087) );
  XNOR U1713 ( .A(n1089), .B(n1090), .Z(out[54]) );
  XNOR U1714 ( .A(key[1206]), .B(n1091), .Z(n1090) );
  XOR U1715 ( .A(n1092), .B(n1093), .Z(out[53]) );
  XNOR U1716 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U1717 ( .A(n1086), .B(n1096), .Z(n1095) );
  XNOR U1718 ( .A(n1098), .B(n1099), .Z(n1097) );
  NANDN U1719 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U1720 ( .A(n1103), .B(n1104), .Z(n1092) );
  XOR U1721 ( .A(key[1205]), .B(n1105), .Z(n1104) );
  ANDN U1722 ( .B(n1106), .A(n1107), .Z(n1103) );
  XNOR U1723 ( .A(n1108), .B(n1109), .Z(out[52]) );
  XNOR U1724 ( .A(key[1204]), .B(n1110), .Z(n1109) );
  XOR U1725 ( .A(n1111), .B(n1112), .Z(out[51]) );
  XNOR U1726 ( .A(n1113), .B(n1089), .Z(n1112) );
  XNOR U1727 ( .A(n1114), .B(n1115), .Z(n1089) );
  XNOR U1728 ( .A(n1116), .B(n1105), .Z(n1115) );
  ANDN U1729 ( .B(n1117), .A(n1118), .Z(n1105) );
  NOR U1730 ( .A(n1119), .B(n1120), .Z(n1116) );
  XNOR U1731 ( .A(n1121), .B(n1122), .Z(n1111) );
  XOR U1732 ( .A(key[1203]), .B(n1123), .Z(n1122) );
  XOR U1733 ( .A(key[1202]), .B(n1108), .Z(out[50]) );
  XNOR U1734 ( .A(n1088), .B(n1124), .Z(n1108) );
  IV U1735 ( .A(n1123), .Z(n1088) );
  XNOR U1736 ( .A(n1125), .B(n1126), .Z(out[4]) );
  XNOR U1737 ( .A(key[1156]), .B(n1127), .Z(n1126) );
  XOR U1738 ( .A(n1128), .B(n1085), .Z(out[49]) );
  XNOR U1739 ( .A(n1114), .B(n1129), .Z(n1113) );
  XNOR U1740 ( .A(n1130), .B(n1131), .Z(n1129) );
  NANDN U1741 ( .A(n1132), .B(n1101), .Z(n1131) );
  XNOR U1742 ( .A(n1096), .B(n1133), .Z(n1114) );
  XNOR U1743 ( .A(n1134), .B(n1135), .Z(n1133) );
  NANDN U1744 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U1745 ( .A(n1124), .B(n1121), .Z(n1091) );
  XNOR U1746 ( .A(n1096), .B(n1138), .Z(n1121) );
  XNOR U1747 ( .A(n1130), .B(n1139), .Z(n1138) );
  NANDN U1748 ( .A(n1140), .B(n1141), .Z(n1139) );
  OR U1749 ( .A(n1142), .B(n1143), .Z(n1130) );
  XOR U1750 ( .A(n1144), .B(n1134), .Z(n1096) );
  NANDN U1751 ( .A(n1145), .B(n1146), .Z(n1134) );
  ANDN U1752 ( .B(n1147), .A(n1148), .Z(n1144) );
  XOR U1753 ( .A(key[1201]), .B(n1123), .Z(n1128) );
  XOR U1754 ( .A(n1149), .B(n1150), .Z(n1123) );
  XNOR U1755 ( .A(n1151), .B(n1152), .Z(n1150) );
  NANDN U1756 ( .A(n1153), .B(n1106), .Z(n1152) );
  XNOR U1757 ( .A(n1094), .B(n1154), .Z(out[48]) );
  XOR U1758 ( .A(key[1200]), .B(n1124), .Z(n1154) );
  XNOR U1759 ( .A(n1149), .B(n1155), .Z(n1124) );
  XOR U1760 ( .A(n1156), .B(n1098), .Z(n1155) );
  OR U1761 ( .A(n1157), .B(n1142), .Z(n1098) );
  XNOR U1762 ( .A(n1101), .B(n1141), .Z(n1142) );
  ANDN U1763 ( .B(n1141), .A(n1158), .Z(n1156) );
  IV U1764 ( .A(n1110), .Z(n1094) );
  XOR U1765 ( .A(n1102), .B(n1159), .Z(n1110) );
  XOR U1766 ( .A(n1160), .B(n1151), .Z(n1159) );
  XNOR U1767 ( .A(n1120), .B(n1106), .Z(n1117) );
  NOR U1768 ( .A(n1162), .B(n1120), .Z(n1160) );
  XNOR U1769 ( .A(n1149), .B(n1163), .Z(n1102) );
  XNOR U1770 ( .A(n1164), .B(n1165), .Z(n1163) );
  NANDN U1771 ( .A(n1136), .B(n1166), .Z(n1165) );
  XOR U1772 ( .A(n1167), .B(n1164), .Z(n1149) );
  OR U1773 ( .A(n1145), .B(n1168), .Z(n1164) );
  XOR U1774 ( .A(n1169), .B(n1136), .Z(n1145) );
  XNOR U1775 ( .A(n1141), .B(n1106), .Z(n1136) );
  XOR U1776 ( .A(n1170), .B(n1171), .Z(n1106) );
  NANDN U1777 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U1778 ( .A(n1174), .B(n1175), .Z(n1141) );
  NANDN U1779 ( .A(n1172), .B(n1176), .Z(n1175) );
  ANDN U1780 ( .B(n1169), .A(n1177), .Z(n1167) );
  IV U1781 ( .A(n1148), .Z(n1169) );
  XOR U1782 ( .A(n1120), .B(n1101), .Z(n1148) );
  XNOR U1783 ( .A(n1178), .B(n1174), .Z(n1101) );
  NANDN U1784 ( .A(n1179), .B(n1180), .Z(n1174) );
  XOR U1785 ( .A(n1176), .B(n1181), .Z(n1180) );
  ANDN U1786 ( .B(n1181), .A(n1182), .Z(n1178) );
  XOR U1787 ( .A(n1183), .B(n1170), .Z(n1120) );
  NANDN U1788 ( .A(n1179), .B(n1184), .Z(n1170) );
  XOR U1789 ( .A(n1185), .B(n1173), .Z(n1184) );
  XNOR U1790 ( .A(n1186), .B(n1187), .Z(n1172) );
  XOR U1791 ( .A(n1188), .B(n1189), .Z(n1187) );
  XNOR U1792 ( .A(n1190), .B(n1191), .Z(n1186) );
  XNOR U1793 ( .A(n1192), .B(n1193), .Z(n1191) );
  ANDN U1794 ( .B(n1185), .A(n1189), .Z(n1192) );
  ANDN U1795 ( .B(n1185), .A(n1182), .Z(n1183) );
  XNOR U1796 ( .A(n1188), .B(n1194), .Z(n1182) );
  XOR U1797 ( .A(n1195), .B(n1193), .Z(n1194) );
  NAND U1798 ( .A(n1196), .B(n1197), .Z(n1193) );
  XNOR U1799 ( .A(n1190), .B(n1173), .Z(n1197) );
  IV U1800 ( .A(n1185), .Z(n1190) );
  XNOR U1801 ( .A(n1176), .B(n1189), .Z(n1196) );
  IV U1802 ( .A(n1181), .Z(n1189) );
  XOR U1803 ( .A(n1198), .B(n1199), .Z(n1181) );
  XNOR U1804 ( .A(n1200), .B(n1201), .Z(n1199) );
  XNOR U1805 ( .A(n1202), .B(n1203), .Z(n1198) );
  NOR U1806 ( .A(n1119), .B(n1162), .Z(n1202) );
  AND U1807 ( .A(n1173), .B(n1176), .Z(n1195) );
  XNOR U1808 ( .A(n1173), .B(n1176), .Z(n1188) );
  XNOR U1809 ( .A(n1204), .B(n1205), .Z(n1176) );
  XNOR U1810 ( .A(n1206), .B(n1201), .Z(n1205) );
  XOR U1811 ( .A(n1207), .B(n1208), .Z(n1204) );
  XNOR U1812 ( .A(n1209), .B(n1203), .Z(n1208) );
  OR U1813 ( .A(n1118), .B(n1161), .Z(n1203) );
  XNOR U1814 ( .A(n1162), .B(n1153), .Z(n1161) );
  XNOR U1815 ( .A(n1119), .B(n1107), .Z(n1118) );
  ANDN U1816 ( .B(n1210), .A(n1153), .Z(n1209) );
  XNOR U1817 ( .A(n1211), .B(n1212), .Z(n1173) );
  XNOR U1818 ( .A(n1201), .B(n1213), .Z(n1212) );
  XOR U1819 ( .A(n1132), .B(n1207), .Z(n1213) );
  XNOR U1820 ( .A(n1162), .B(n1214), .Z(n1201) );
  XOR U1821 ( .A(n1100), .B(n1215), .Z(n1211) );
  XNOR U1822 ( .A(n1216), .B(n1217), .Z(n1215) );
  ANDN U1823 ( .B(n1218), .A(n1158), .Z(n1216) );
  XNOR U1824 ( .A(n1219), .B(n1220), .Z(n1185) );
  XNOR U1825 ( .A(n1206), .B(n1221), .Z(n1220) );
  XNOR U1826 ( .A(n1140), .B(n1200), .Z(n1221) );
  XOR U1827 ( .A(n1207), .B(n1222), .Z(n1200) );
  XNOR U1828 ( .A(n1223), .B(n1224), .Z(n1222) );
  NAND U1829 ( .A(n1166), .B(n1137), .Z(n1224) );
  XNOR U1830 ( .A(n1225), .B(n1223), .Z(n1207) );
  NANDN U1831 ( .A(n1168), .B(n1146), .Z(n1223) );
  XOR U1832 ( .A(n1147), .B(n1137), .Z(n1146) );
  XNOR U1833 ( .A(n1218), .B(n1107), .Z(n1137) );
  XOR U1834 ( .A(n1177), .B(n1166), .Z(n1168) );
  XNOR U1835 ( .A(n1158), .B(n1226), .Z(n1166) );
  ANDN U1836 ( .B(n1147), .A(n1177), .Z(n1225) );
  XNOR U1837 ( .A(n1100), .B(n1162), .Z(n1177) );
  XOR U1838 ( .A(n1227), .B(n1228), .Z(n1162) );
  XNOR U1839 ( .A(n1229), .B(n1230), .Z(n1228) );
  XOR U1840 ( .A(n1226), .B(n1210), .Z(n1206) );
  IV U1841 ( .A(n1107), .Z(n1210) );
  XOR U1842 ( .A(n1231), .B(n1232), .Z(n1107) );
  XOR U1843 ( .A(n1233), .B(n1230), .Z(n1232) );
  IV U1844 ( .A(n1153), .Z(n1226) );
  XOR U1845 ( .A(n1230), .B(n1234), .Z(n1153) );
  XNOR U1846 ( .A(n1235), .B(n1236), .Z(n1219) );
  XNOR U1847 ( .A(n1237), .B(n1217), .Z(n1236) );
  OR U1848 ( .A(n1143), .B(n1157), .Z(n1217) );
  XNOR U1849 ( .A(n1100), .B(n1158), .Z(n1157) );
  IV U1850 ( .A(n1235), .Z(n1158) );
  XOR U1851 ( .A(n1132), .B(n1218), .Z(n1143) );
  IV U1852 ( .A(n1140), .Z(n1218) );
  XOR U1853 ( .A(n1214), .B(n1238), .Z(n1140) );
  XNOR U1854 ( .A(n1239), .B(n1227), .Z(n1238) );
  XOR U1855 ( .A(n1240), .B(n1241), .Z(n1227) );
  XNOR U1856 ( .A(n1242), .B(n1243), .Z(n1241) );
  XNOR U1857 ( .A(key[1170]), .B(n640), .Z(n1240) );
  IV U1858 ( .A(n1119), .Z(n1214) );
  XOR U1859 ( .A(n1231), .B(n1244), .Z(n1119) );
  XOR U1860 ( .A(n1230), .B(n1245), .Z(n1244) );
  NOR U1861 ( .A(n1132), .B(n1100), .Z(n1237) );
  XOR U1862 ( .A(n1231), .B(n1246), .Z(n1132) );
  XOR U1863 ( .A(n1230), .B(n1247), .Z(n1246) );
  XOR U1864 ( .A(n1248), .B(n1249), .Z(n1230) );
  XNOR U1865 ( .A(n1100), .B(n1250), .Z(n1249) );
  XOR U1866 ( .A(n620), .B(n1251), .Z(n1248) );
  XNOR U1867 ( .A(key[1174]), .B(n616), .Z(n1251) );
  XNOR U1868 ( .A(n1252), .B(n1253), .Z(n620) );
  IV U1869 ( .A(n1234), .Z(n1231) );
  XOR U1870 ( .A(n1254), .B(n1255), .Z(n1234) );
  XNOR U1871 ( .A(n1256), .B(n613), .Z(n1255) );
  XNOR U1872 ( .A(n1257), .B(n1258), .Z(n613) );
  XNOR U1873 ( .A(key[1173]), .B(n1259), .Z(n1254) );
  XOR U1874 ( .A(n1260), .B(n1261), .Z(n1235) );
  XNOR U1875 ( .A(n1247), .B(n1245), .Z(n1261) );
  XNOR U1876 ( .A(n1262), .B(n1263), .Z(n1245) );
  XOR U1877 ( .A(n1253), .B(n607), .Z(n1263) );
  XNOR U1878 ( .A(n1264), .B(n1265), .Z(n607) );
  XOR U1879 ( .A(n1266), .B(n1267), .Z(n1253) );
  XNOR U1880 ( .A(key[1175]), .B(n1268), .Z(n1262) );
  XNOR U1881 ( .A(n1269), .B(n1270), .Z(n1247) );
  XOR U1882 ( .A(n598), .B(n1271), .Z(n1270) );
  XOR U1883 ( .A(n1272), .B(n1273), .Z(n598) );
  XOR U1884 ( .A(n1274), .B(n1256), .Z(n1273) );
  XOR U1885 ( .A(n1266), .B(n1275), .Z(n1272) );
  XNOR U1886 ( .A(key[1172]), .B(n1276), .Z(n1269) );
  XNOR U1887 ( .A(n1100), .B(n1229), .Z(n1260) );
  XOR U1888 ( .A(n1277), .B(n1278), .Z(n1229) );
  XNOR U1889 ( .A(n1279), .B(n1280), .Z(n1278) );
  XNOR U1890 ( .A(n633), .B(n1239), .Z(n1280) );
  IV U1891 ( .A(n1233), .Z(n1239) );
  XNOR U1892 ( .A(n1281), .B(n1282), .Z(n1233) );
  XNOR U1893 ( .A(n1283), .B(n624), .Z(n1282) );
  XNOR U1894 ( .A(key[1169]), .B(n642), .Z(n1281) );
  XNOR U1895 ( .A(n1266), .B(n1276), .Z(n633) );
  XOR U1896 ( .A(n649), .B(n1284), .Z(n1277) );
  XOR U1897 ( .A(key[1171]), .B(n645), .Z(n1284) );
  XNOR U1898 ( .A(n1285), .B(n1286), .Z(n1100) );
  XOR U1899 ( .A(n1287), .B(n608), .Z(n1286) );
  XNOR U1900 ( .A(key[1168]), .B(n1288), .Z(n1285) );
  XOR U1901 ( .A(n1289), .B(n1290), .Z(out[47]) );
  XOR U1902 ( .A(n1291), .B(n1292), .Z(n1289) );
  XNOR U1903 ( .A(key[1199]), .B(n1293), .Z(n1292) );
  XNOR U1904 ( .A(n1294), .B(n1295), .Z(out[46]) );
  XNOR U1905 ( .A(key[1198]), .B(n1296), .Z(n1295) );
  XOR U1906 ( .A(n1297), .B(n1298), .Z(out[45]) );
  XNOR U1907 ( .A(n1299), .B(n1300), .Z(n1298) );
  XOR U1908 ( .A(n1291), .B(n1301), .Z(n1300) );
  XNOR U1909 ( .A(n1303), .B(n1304), .Z(n1302) );
  NANDN U1910 ( .A(n1305), .B(n1306), .Z(n1304) );
  XOR U1911 ( .A(n1308), .B(n1309), .Z(n1297) );
  XOR U1912 ( .A(key[1197]), .B(n1310), .Z(n1309) );
  ANDN U1913 ( .B(n1311), .A(n1312), .Z(n1308) );
  XNOR U1914 ( .A(n1313), .B(n1314), .Z(out[44]) );
  XNOR U1915 ( .A(key[1196]), .B(n1315), .Z(n1314) );
  XOR U1916 ( .A(n1316), .B(n1317), .Z(out[43]) );
  XNOR U1917 ( .A(n1318), .B(n1294), .Z(n1317) );
  XNOR U1918 ( .A(n1319), .B(n1320), .Z(n1294) );
  XNOR U1919 ( .A(n1321), .B(n1310), .Z(n1320) );
  ANDN U1920 ( .B(n1322), .A(n1323), .Z(n1310) );
  NOR U1921 ( .A(n1324), .B(n1325), .Z(n1321) );
  XNOR U1922 ( .A(n1326), .B(n1327), .Z(n1316) );
  XOR U1923 ( .A(key[1195]), .B(n1328), .Z(n1327) );
  XOR U1924 ( .A(key[1194]), .B(n1313), .Z(out[42]) );
  XNOR U1925 ( .A(n1293), .B(n1329), .Z(n1313) );
  IV U1926 ( .A(n1328), .Z(n1293) );
  XOR U1927 ( .A(n1330), .B(n1290), .Z(out[41]) );
  XNOR U1928 ( .A(n1319), .B(n1331), .Z(n1318) );
  XNOR U1929 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1930 ( .A(n1334), .B(n1306), .Z(n1333) );
  XNOR U1931 ( .A(n1301), .B(n1335), .Z(n1319) );
  XNOR U1932 ( .A(n1336), .B(n1337), .Z(n1335) );
  NANDN U1933 ( .A(n1338), .B(n1339), .Z(n1337) );
  XOR U1934 ( .A(n1329), .B(n1326), .Z(n1296) );
  XNOR U1935 ( .A(n1301), .B(n1340), .Z(n1326) );
  XNOR U1936 ( .A(n1332), .B(n1341), .Z(n1340) );
  NANDN U1937 ( .A(n1342), .B(n1343), .Z(n1341) );
  OR U1938 ( .A(n1344), .B(n1345), .Z(n1332) );
  XOR U1939 ( .A(n1346), .B(n1336), .Z(n1301) );
  NANDN U1940 ( .A(n1347), .B(n1348), .Z(n1336) );
  ANDN U1941 ( .B(n1349), .A(n1350), .Z(n1346) );
  XOR U1942 ( .A(key[1193]), .B(n1328), .Z(n1330) );
  XOR U1943 ( .A(n1351), .B(n1352), .Z(n1328) );
  XNOR U1944 ( .A(n1353), .B(n1354), .Z(n1352) );
  NANDN U1945 ( .A(n1355), .B(n1311), .Z(n1354) );
  XNOR U1946 ( .A(n1299), .B(n1356), .Z(out[40]) );
  XOR U1947 ( .A(key[1192]), .B(n1329), .Z(n1356) );
  XNOR U1948 ( .A(n1351), .B(n1357), .Z(n1329) );
  XOR U1949 ( .A(n1358), .B(n1303), .Z(n1357) );
  OR U1950 ( .A(n1359), .B(n1344), .Z(n1303) );
  XNOR U1951 ( .A(n1306), .B(n1343), .Z(n1344) );
  ANDN U1952 ( .B(n1343), .A(n1360), .Z(n1358) );
  IV U1953 ( .A(n1315), .Z(n1299) );
  XOR U1954 ( .A(n1307), .B(n1361), .Z(n1315) );
  XOR U1955 ( .A(n1362), .B(n1353), .Z(n1361) );
  XNOR U1956 ( .A(n1325), .B(n1311), .Z(n1322) );
  NOR U1957 ( .A(n1364), .B(n1325), .Z(n1362) );
  XNOR U1958 ( .A(n1351), .B(n1365), .Z(n1307) );
  XNOR U1959 ( .A(n1366), .B(n1367), .Z(n1365) );
  NANDN U1960 ( .A(n1338), .B(n1368), .Z(n1367) );
  XOR U1961 ( .A(n1369), .B(n1366), .Z(n1351) );
  OR U1962 ( .A(n1347), .B(n1370), .Z(n1366) );
  XOR U1963 ( .A(n1371), .B(n1338), .Z(n1347) );
  XNOR U1964 ( .A(n1343), .B(n1311), .Z(n1338) );
  XOR U1965 ( .A(n1372), .B(n1373), .Z(n1311) );
  NANDN U1966 ( .A(n1374), .B(n1375), .Z(n1373) );
  XOR U1967 ( .A(n1376), .B(n1377), .Z(n1343) );
  NANDN U1968 ( .A(n1374), .B(n1378), .Z(n1377) );
  ANDN U1969 ( .B(n1371), .A(n1379), .Z(n1369) );
  IV U1970 ( .A(n1350), .Z(n1371) );
  XOR U1971 ( .A(n1325), .B(n1306), .Z(n1350) );
  XNOR U1972 ( .A(n1380), .B(n1376), .Z(n1306) );
  NANDN U1973 ( .A(n1381), .B(n1382), .Z(n1376) );
  XOR U1974 ( .A(n1378), .B(n1383), .Z(n1382) );
  ANDN U1975 ( .B(n1383), .A(n1384), .Z(n1380) );
  XOR U1976 ( .A(n1385), .B(n1372), .Z(n1325) );
  NANDN U1977 ( .A(n1381), .B(n1386), .Z(n1372) );
  XOR U1978 ( .A(n1387), .B(n1375), .Z(n1386) );
  XNOR U1979 ( .A(n1388), .B(n1389), .Z(n1374) );
  XOR U1980 ( .A(n1390), .B(n1391), .Z(n1389) );
  XNOR U1981 ( .A(n1392), .B(n1393), .Z(n1388) );
  XNOR U1982 ( .A(n1394), .B(n1395), .Z(n1393) );
  ANDN U1983 ( .B(n1387), .A(n1391), .Z(n1394) );
  ANDN U1984 ( .B(n1387), .A(n1384), .Z(n1385) );
  XNOR U1985 ( .A(n1390), .B(n1396), .Z(n1384) );
  XOR U1986 ( .A(n1397), .B(n1395), .Z(n1396) );
  NAND U1987 ( .A(n1398), .B(n1399), .Z(n1395) );
  XNOR U1988 ( .A(n1392), .B(n1375), .Z(n1399) );
  IV U1989 ( .A(n1387), .Z(n1392) );
  XNOR U1990 ( .A(n1378), .B(n1391), .Z(n1398) );
  IV U1991 ( .A(n1383), .Z(n1391) );
  XOR U1992 ( .A(n1400), .B(n1401), .Z(n1383) );
  XNOR U1993 ( .A(n1402), .B(n1403), .Z(n1401) );
  XNOR U1994 ( .A(n1404), .B(n1405), .Z(n1400) );
  NOR U1995 ( .A(n1324), .B(n1364), .Z(n1404) );
  AND U1996 ( .A(n1375), .B(n1378), .Z(n1397) );
  XNOR U1997 ( .A(n1375), .B(n1378), .Z(n1390) );
  XNOR U1998 ( .A(n1406), .B(n1407), .Z(n1378) );
  XNOR U1999 ( .A(n1408), .B(n1403), .Z(n1407) );
  XOR U2000 ( .A(n1409), .B(n1410), .Z(n1406) );
  XNOR U2001 ( .A(n1411), .B(n1405), .Z(n1410) );
  OR U2002 ( .A(n1323), .B(n1363), .Z(n1405) );
  XNOR U2003 ( .A(n1364), .B(n1355), .Z(n1363) );
  XNOR U2004 ( .A(n1324), .B(n1312), .Z(n1323) );
  ANDN U2005 ( .B(n1412), .A(n1355), .Z(n1411) );
  XNOR U2006 ( .A(n1413), .B(n1414), .Z(n1375) );
  XNOR U2007 ( .A(n1403), .B(n1415), .Z(n1414) );
  XOR U2008 ( .A(n1334), .B(n1409), .Z(n1415) );
  XNOR U2009 ( .A(n1364), .B(n1416), .Z(n1403) );
  XOR U2010 ( .A(n1305), .B(n1417), .Z(n1413) );
  XNOR U2011 ( .A(n1418), .B(n1419), .Z(n1417) );
  ANDN U2012 ( .B(n1420), .A(n1360), .Z(n1418) );
  XNOR U2013 ( .A(n1421), .B(n1422), .Z(n1387) );
  XNOR U2014 ( .A(n1408), .B(n1423), .Z(n1422) );
  XNOR U2015 ( .A(n1342), .B(n1402), .Z(n1423) );
  XOR U2016 ( .A(n1409), .B(n1424), .Z(n1402) );
  XNOR U2017 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U2018 ( .A(n1368), .B(n1339), .Z(n1426) );
  XNOR U2019 ( .A(n1427), .B(n1425), .Z(n1409) );
  NANDN U2020 ( .A(n1370), .B(n1348), .Z(n1425) );
  XOR U2021 ( .A(n1349), .B(n1339), .Z(n1348) );
  XNOR U2022 ( .A(n1420), .B(n1312), .Z(n1339) );
  XOR U2023 ( .A(n1379), .B(n1368), .Z(n1370) );
  XNOR U2024 ( .A(n1360), .B(n1428), .Z(n1368) );
  ANDN U2025 ( .B(n1349), .A(n1379), .Z(n1427) );
  XNOR U2026 ( .A(n1305), .B(n1364), .Z(n1379) );
  XOR U2027 ( .A(n1429), .B(n1430), .Z(n1364) );
  XNOR U2028 ( .A(n1431), .B(n1432), .Z(n1430) );
  XOR U2029 ( .A(n1428), .B(n1412), .Z(n1408) );
  IV U2030 ( .A(n1312), .Z(n1412) );
  XOR U2031 ( .A(n1433), .B(n1434), .Z(n1312) );
  XOR U2032 ( .A(n1435), .B(n1432), .Z(n1434) );
  IV U2033 ( .A(n1355), .Z(n1428) );
  XOR U2034 ( .A(n1432), .B(n1436), .Z(n1355) );
  XNOR U2035 ( .A(n1437), .B(n1438), .Z(n1421) );
  XNOR U2036 ( .A(n1439), .B(n1419), .Z(n1438) );
  OR U2037 ( .A(n1345), .B(n1359), .Z(n1419) );
  XNOR U2038 ( .A(n1305), .B(n1360), .Z(n1359) );
  IV U2039 ( .A(n1437), .Z(n1360) );
  XOR U2040 ( .A(n1334), .B(n1420), .Z(n1345) );
  IV U2041 ( .A(n1342), .Z(n1420) );
  XOR U2042 ( .A(n1416), .B(n1440), .Z(n1342) );
  XNOR U2043 ( .A(n1441), .B(n1429), .Z(n1440) );
  XOR U2044 ( .A(n1442), .B(n1443), .Z(n1429) );
  XNOR U2045 ( .A(n836), .B(n1444), .Z(n1443) );
  XOR U2046 ( .A(n1445), .B(n1446), .Z(n1442) );
  XNOR U2047 ( .A(key[1258]), .B(n1447), .Z(n1446) );
  IV U2048 ( .A(n1324), .Z(n1416) );
  XOR U2049 ( .A(n1433), .B(n1448), .Z(n1324) );
  XOR U2050 ( .A(n1432), .B(n1449), .Z(n1448) );
  NOR U2051 ( .A(n1334), .B(n1305), .Z(n1439) );
  XOR U2052 ( .A(n1433), .B(n1450), .Z(n1334) );
  XOR U2053 ( .A(n1432), .B(n1451), .Z(n1450) );
  XOR U2054 ( .A(n1452), .B(n1453), .Z(n1432) );
  XNOR U2055 ( .A(n1305), .B(n1454), .Z(n1453) );
  XNOR U2056 ( .A(n1455), .B(n1456), .Z(n1452) );
  XNOR U2057 ( .A(key[1262]), .B(n851), .Z(n1456) );
  XOR U2058 ( .A(n822), .B(n1457), .Z(n851) );
  IV U2059 ( .A(n1436), .Z(n1433) );
  XOR U2060 ( .A(n1458), .B(n1459), .Z(n1436) );
  XOR U2061 ( .A(n1460), .B(n1461), .Z(n1459) );
  XOR U2062 ( .A(n1462), .B(n1463), .Z(n1458) );
  XNOR U2063 ( .A(key[1261]), .B(n1464), .Z(n1463) );
  XOR U2064 ( .A(n1465), .B(n1466), .Z(n1437) );
  XNOR U2065 ( .A(n1451), .B(n1449), .Z(n1466) );
  XNOR U2066 ( .A(n1467), .B(n1468), .Z(n1449) );
  XOR U2067 ( .A(n1469), .B(n1470), .Z(n1468) );
  XNOR U2068 ( .A(key[1263]), .B(n1471), .Z(n1467) );
  XNOR U2069 ( .A(n1472), .B(n1473), .Z(n1451) );
  XOR U2070 ( .A(n1474), .B(n1475), .Z(n1473) );
  XNOR U2071 ( .A(n1476), .B(n1477), .Z(n1472) );
  XNOR U2072 ( .A(key[1260]), .B(n807), .Z(n1477) );
  XNOR U2073 ( .A(n822), .B(n1478), .Z(n807) );
  XNOR U2074 ( .A(n1305), .B(n1431), .Z(n1465) );
  XOR U2075 ( .A(n1479), .B(n1480), .Z(n1431) );
  XNOR U2076 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U2077 ( .A(n1483), .B(n1441), .Z(n1482) );
  IV U2078 ( .A(n1435), .Z(n1441) );
  XNOR U2079 ( .A(n1484), .B(n1485), .Z(n1435) );
  XNOR U2080 ( .A(n1486), .B(n1487), .Z(n1485) );
  XOR U2081 ( .A(n1488), .B(n1489), .Z(n1484) );
  XNOR U2082 ( .A(key[1257]), .B(n857), .Z(n1489) );
  XNOR U2083 ( .A(n833), .B(n1490), .Z(n1479) );
  XNOR U2084 ( .A(key[1259]), .B(n844), .Z(n1490) );
  IV U2085 ( .A(n1491), .Z(n844) );
  XOR U2086 ( .A(n822), .B(n1492), .Z(n833) );
  XNOR U2087 ( .A(n1493), .B(n1494), .Z(n1305) );
  XNOR U2088 ( .A(n822), .B(n1495), .Z(n1494) );
  XNOR U2089 ( .A(n855), .B(n1496), .Z(n1493) );
  XOR U2090 ( .A(key[1256]), .B(n1497), .Z(n1496) );
  XOR U2091 ( .A(n1498), .B(n1499), .Z(out[3]) );
  XNOR U2092 ( .A(n1500), .B(n663), .Z(n1499) );
  XNOR U2093 ( .A(n1501), .B(n1502), .Z(n663) );
  XNOR U2094 ( .A(n1503), .B(n898), .Z(n1502) );
  ANDN U2095 ( .B(n1504), .A(n1505), .Z(n898) );
  NOR U2096 ( .A(n1506), .B(n1507), .Z(n1503) );
  XNOR U2097 ( .A(n1508), .B(n1509), .Z(n1498) );
  XOR U2098 ( .A(key[1155]), .B(n1510), .Z(n1509) );
  XOR U2099 ( .A(n1511), .B(n1512), .Z(out[39]) );
  XOR U2100 ( .A(n1513), .B(n1514), .Z(n1511) );
  XNOR U2101 ( .A(key[1191]), .B(n1515), .Z(n1514) );
  XNOR U2102 ( .A(n1516), .B(n1517), .Z(out[38]) );
  XNOR U2103 ( .A(key[1190]), .B(n1518), .Z(n1517) );
  XOR U2104 ( .A(n1519), .B(n1520), .Z(out[37]) );
  XNOR U2105 ( .A(n1521), .B(n1522), .Z(n1520) );
  XOR U2106 ( .A(n1513), .B(n1523), .Z(n1522) );
  XNOR U2107 ( .A(n1525), .B(n1526), .Z(n1524) );
  NANDN U2108 ( .A(n1527), .B(n1528), .Z(n1526) );
  XOR U2109 ( .A(n1530), .B(n1531), .Z(n1519) );
  XOR U2110 ( .A(key[1189]), .B(n1532), .Z(n1531) );
  ANDN U2111 ( .B(n1533), .A(n1534), .Z(n1530) );
  XNOR U2112 ( .A(n1535), .B(n1536), .Z(out[36]) );
  XNOR U2113 ( .A(key[1188]), .B(n1537), .Z(n1536) );
  XOR U2114 ( .A(n1538), .B(n1539), .Z(out[35]) );
  XNOR U2115 ( .A(n1540), .B(n1516), .Z(n1539) );
  XNOR U2116 ( .A(n1541), .B(n1542), .Z(n1516) );
  XNOR U2117 ( .A(n1543), .B(n1532), .Z(n1542) );
  ANDN U2118 ( .B(n1544), .A(n1545), .Z(n1532) );
  NOR U2119 ( .A(n1546), .B(n1547), .Z(n1543) );
  XNOR U2120 ( .A(n1548), .B(n1549), .Z(n1538) );
  XOR U2121 ( .A(key[1187]), .B(n1550), .Z(n1549) );
  XOR U2122 ( .A(key[1186]), .B(n1535), .Z(out[34]) );
  XNOR U2123 ( .A(n1515), .B(n1551), .Z(n1535) );
  IV U2124 ( .A(n1550), .Z(n1515) );
  XOR U2125 ( .A(n1552), .B(n1512), .Z(out[33]) );
  XNOR U2126 ( .A(n1541), .B(n1553), .Z(n1540) );
  XNOR U2127 ( .A(n1554), .B(n1555), .Z(n1553) );
  NANDN U2128 ( .A(n1556), .B(n1528), .Z(n1555) );
  XNOR U2129 ( .A(n1523), .B(n1557), .Z(n1541) );
  XNOR U2130 ( .A(n1558), .B(n1559), .Z(n1557) );
  NANDN U2131 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U2132 ( .A(n1551), .B(n1548), .Z(n1518) );
  XNOR U2133 ( .A(n1523), .B(n1562), .Z(n1548) );
  XNOR U2134 ( .A(n1554), .B(n1563), .Z(n1562) );
  NANDN U2135 ( .A(n1564), .B(n1565), .Z(n1563) );
  OR U2136 ( .A(n1566), .B(n1567), .Z(n1554) );
  XOR U2137 ( .A(n1568), .B(n1558), .Z(n1523) );
  NANDN U2138 ( .A(n1569), .B(n1570), .Z(n1558) );
  ANDN U2139 ( .B(n1571), .A(n1572), .Z(n1568) );
  XOR U2140 ( .A(key[1185]), .B(n1550), .Z(n1552) );
  XOR U2141 ( .A(n1573), .B(n1574), .Z(n1550) );
  XNOR U2142 ( .A(n1575), .B(n1576), .Z(n1574) );
  NANDN U2143 ( .A(n1577), .B(n1533), .Z(n1576) );
  XNOR U2144 ( .A(n1521), .B(n1578), .Z(out[32]) );
  XOR U2145 ( .A(key[1184]), .B(n1551), .Z(n1578) );
  XNOR U2146 ( .A(n1573), .B(n1579), .Z(n1551) );
  XOR U2147 ( .A(n1580), .B(n1525), .Z(n1579) );
  OR U2148 ( .A(n1581), .B(n1566), .Z(n1525) );
  XNOR U2149 ( .A(n1528), .B(n1565), .Z(n1566) );
  ANDN U2150 ( .B(n1582), .A(n1583), .Z(n1580) );
  IV U2151 ( .A(n1537), .Z(n1521) );
  XOR U2152 ( .A(n1529), .B(n1584), .Z(n1537) );
  XOR U2153 ( .A(n1585), .B(n1575), .Z(n1584) );
  XNOR U2154 ( .A(n1547), .B(n1533), .Z(n1544) );
  NOR U2155 ( .A(n1587), .B(n1547), .Z(n1585) );
  XNOR U2156 ( .A(n1573), .B(n1588), .Z(n1529) );
  XNOR U2157 ( .A(n1589), .B(n1590), .Z(n1588) );
  NANDN U2158 ( .A(n1560), .B(n1591), .Z(n1590) );
  XOR U2159 ( .A(n1592), .B(n1589), .Z(n1573) );
  OR U2160 ( .A(n1569), .B(n1593), .Z(n1589) );
  XOR U2161 ( .A(n1594), .B(n1560), .Z(n1569) );
  XNOR U2162 ( .A(n1565), .B(n1533), .Z(n1560) );
  XOR U2163 ( .A(n1595), .B(n1596), .Z(n1533) );
  NANDN U2164 ( .A(n1597), .B(n1598), .Z(n1596) );
  IV U2165 ( .A(n1583), .Z(n1565) );
  XNOR U2166 ( .A(n1599), .B(n1600), .Z(n1583) );
  NANDN U2167 ( .A(n1597), .B(n1601), .Z(n1600) );
  ANDN U2168 ( .B(n1594), .A(n1602), .Z(n1592) );
  IV U2169 ( .A(n1572), .Z(n1594) );
  XOR U2170 ( .A(n1547), .B(n1528), .Z(n1572) );
  XNOR U2171 ( .A(n1603), .B(n1599), .Z(n1528) );
  NANDN U2172 ( .A(n1604), .B(n1605), .Z(n1599) );
  XOR U2173 ( .A(n1601), .B(n1606), .Z(n1605) );
  ANDN U2174 ( .B(n1606), .A(n1607), .Z(n1603) );
  XOR U2175 ( .A(n1608), .B(n1595), .Z(n1547) );
  NANDN U2176 ( .A(n1604), .B(n1609), .Z(n1595) );
  XOR U2177 ( .A(n1610), .B(n1598), .Z(n1609) );
  XNOR U2178 ( .A(n1611), .B(n1612), .Z(n1597) );
  XOR U2179 ( .A(n1613), .B(n1614), .Z(n1612) );
  XNOR U2180 ( .A(n1615), .B(n1616), .Z(n1611) );
  XNOR U2181 ( .A(n1617), .B(n1618), .Z(n1616) );
  ANDN U2182 ( .B(n1610), .A(n1614), .Z(n1617) );
  ANDN U2183 ( .B(n1610), .A(n1607), .Z(n1608) );
  XNOR U2184 ( .A(n1613), .B(n1619), .Z(n1607) );
  XOR U2185 ( .A(n1620), .B(n1618), .Z(n1619) );
  NAND U2186 ( .A(n1621), .B(n1622), .Z(n1618) );
  XNOR U2187 ( .A(n1615), .B(n1598), .Z(n1622) );
  IV U2188 ( .A(n1610), .Z(n1615) );
  XNOR U2189 ( .A(n1601), .B(n1614), .Z(n1621) );
  IV U2190 ( .A(n1606), .Z(n1614) );
  XOR U2191 ( .A(n1623), .B(n1624), .Z(n1606) );
  XNOR U2192 ( .A(n1625), .B(n1626), .Z(n1624) );
  XNOR U2193 ( .A(n1627), .B(n1628), .Z(n1623) );
  NOR U2194 ( .A(n1546), .B(n1587), .Z(n1627) );
  AND U2195 ( .A(n1598), .B(n1601), .Z(n1620) );
  XNOR U2196 ( .A(n1598), .B(n1601), .Z(n1613) );
  XNOR U2197 ( .A(n1629), .B(n1630), .Z(n1601) );
  XNOR U2198 ( .A(n1631), .B(n1626), .Z(n1630) );
  XOR U2199 ( .A(n1632), .B(n1633), .Z(n1629) );
  XNOR U2200 ( .A(n1634), .B(n1628), .Z(n1633) );
  OR U2201 ( .A(n1545), .B(n1586), .Z(n1628) );
  XNOR U2202 ( .A(n1587), .B(n1577), .Z(n1586) );
  XNOR U2203 ( .A(n1546), .B(n1534), .Z(n1545) );
  ANDN U2204 ( .B(n1635), .A(n1577), .Z(n1634) );
  XNOR U2205 ( .A(n1636), .B(n1637), .Z(n1598) );
  XNOR U2206 ( .A(n1626), .B(n1638), .Z(n1637) );
  XOR U2207 ( .A(n1556), .B(n1632), .Z(n1638) );
  XNOR U2208 ( .A(n1587), .B(n1639), .Z(n1626) );
  XNOR U2209 ( .A(n1640), .B(n1641), .Z(n1636) );
  XNOR U2210 ( .A(n1642), .B(n1643), .Z(n1641) );
  ANDN U2211 ( .B(n1582), .A(n1564), .Z(n1642) );
  XNOR U2212 ( .A(n1644), .B(n1645), .Z(n1610) );
  XNOR U2213 ( .A(n1631), .B(n1646), .Z(n1645) );
  XNOR U2214 ( .A(n1564), .B(n1625), .Z(n1646) );
  XOR U2215 ( .A(n1632), .B(n1647), .Z(n1625) );
  XNOR U2216 ( .A(n1648), .B(n1649), .Z(n1647) );
  NAND U2217 ( .A(n1591), .B(n1561), .Z(n1649) );
  XNOR U2218 ( .A(n1650), .B(n1648), .Z(n1632) );
  NANDN U2219 ( .A(n1593), .B(n1570), .Z(n1648) );
  XOR U2220 ( .A(n1571), .B(n1561), .Z(n1570) );
  XNOR U2221 ( .A(n1651), .B(n1534), .Z(n1561) );
  XOR U2222 ( .A(n1602), .B(n1591), .Z(n1593) );
  XOR U2223 ( .A(n1582), .B(n1652), .Z(n1591) );
  ANDN U2224 ( .B(n1571), .A(n1602), .Z(n1650) );
  XOR U2225 ( .A(n1640), .B(n1587), .Z(n1602) );
  XOR U2226 ( .A(n1653), .B(n1654), .Z(n1587) );
  XNOR U2227 ( .A(n1655), .B(n1656), .Z(n1654) );
  XOR U2228 ( .A(n1657), .B(n1639), .Z(n1571) );
  XOR U2229 ( .A(n1652), .B(n1635), .Z(n1631) );
  IV U2230 ( .A(n1534), .Z(n1635) );
  XOR U2231 ( .A(n1658), .B(n1659), .Z(n1534) );
  XNOR U2232 ( .A(n1660), .B(n1656), .Z(n1659) );
  IV U2233 ( .A(n1577), .Z(n1652) );
  XOR U2234 ( .A(n1656), .B(n1661), .Z(n1577) );
  XNOR U2235 ( .A(n1582), .B(n1662), .Z(n1644) );
  XNOR U2236 ( .A(n1663), .B(n1643), .Z(n1662) );
  OR U2237 ( .A(n1567), .B(n1581), .Z(n1643) );
  XNOR U2238 ( .A(n1640), .B(n1582), .Z(n1581) );
  XOR U2239 ( .A(n1556), .B(n1651), .Z(n1567) );
  IV U2240 ( .A(n1564), .Z(n1651) );
  XOR U2241 ( .A(n1639), .B(n1664), .Z(n1564) );
  XNOR U2242 ( .A(n1660), .B(n1653), .Z(n1664) );
  XOR U2243 ( .A(n1665), .B(n1666), .Z(n1653) );
  XNOR U2244 ( .A(n1667), .B(n178), .Z(n1666) );
  XOR U2245 ( .A(key[1218]), .B(n220), .Z(n1665) );
  IV U2246 ( .A(n1546), .Z(n1639) );
  XOR U2247 ( .A(n1658), .B(n1668), .Z(n1546) );
  XOR U2248 ( .A(n1656), .B(n1669), .Z(n1668) );
  ANDN U2249 ( .B(n1657), .A(n1527), .Z(n1663) );
  IV U2250 ( .A(n1556), .Z(n1657) );
  XOR U2251 ( .A(n1658), .B(n1670), .Z(n1556) );
  XOR U2252 ( .A(n1656), .B(n1671), .Z(n1670) );
  XOR U2253 ( .A(n1672), .B(n1673), .Z(n1656) );
  XNOR U2254 ( .A(n189), .B(n1527), .Z(n1673) );
  IV U2255 ( .A(n1640), .Z(n1527) );
  XOR U2256 ( .A(n1674), .B(n1675), .Z(n189) );
  XNOR U2257 ( .A(n194), .B(n1676), .Z(n1672) );
  XNOR U2258 ( .A(key[1222]), .B(n1677), .Z(n1676) );
  IV U2259 ( .A(n1661), .Z(n1658) );
  XOR U2260 ( .A(n1678), .B(n1679), .Z(n1661) );
  XOR U2261 ( .A(n1680), .B(n195), .Z(n1679) );
  XOR U2262 ( .A(n1681), .B(n1682), .Z(n195) );
  XNOR U2263 ( .A(key[1221]), .B(n1683), .Z(n1678) );
  XOR U2264 ( .A(n1684), .B(n1685), .Z(n1582) );
  XNOR U2265 ( .A(n1671), .B(n1669), .Z(n1685) );
  XNOR U2266 ( .A(n1686), .B(n1687), .Z(n1669) );
  XOR U2267 ( .A(n1675), .B(n204), .Z(n1687) );
  XNOR U2268 ( .A(n1688), .B(n1689), .Z(n204) );
  XNOR U2269 ( .A(n1690), .B(n1691), .Z(n1675) );
  XNOR U2270 ( .A(key[1223]), .B(n1692), .Z(n1686) );
  XNOR U2271 ( .A(n1693), .B(n1694), .Z(n1671) );
  XOR U2272 ( .A(n210), .B(n209), .Z(n1694) );
  XOR U2273 ( .A(n1695), .B(n1696), .Z(n209) );
  XOR U2274 ( .A(n1683), .B(n1690), .Z(n210) );
  XNOR U2275 ( .A(n1697), .B(n1698), .Z(n1693) );
  XNOR U2276 ( .A(key[1220]), .B(n1699), .Z(n1698) );
  XOR U2277 ( .A(n1640), .B(n1655), .Z(n1684) );
  XOR U2278 ( .A(n1700), .B(n1701), .Z(n1655) );
  XNOR U2279 ( .A(n1660), .B(n1702), .Z(n1701) );
  XNOR U2280 ( .A(n225), .B(n215), .Z(n1702) );
  XOR U2281 ( .A(n1690), .B(n1697), .Z(n225) );
  XOR U2282 ( .A(n1703), .B(n1704), .Z(n1660) );
  XNOR U2283 ( .A(n1705), .B(n221), .Z(n1704) );
  XOR U2284 ( .A(key[1217]), .B(n1706), .Z(n1703) );
  XNOR U2285 ( .A(n179), .B(n1707), .Z(n1700) );
  XNOR U2286 ( .A(key[1219]), .B(n1708), .Z(n1707) );
  XOR U2287 ( .A(n1709), .B(n1710), .Z(n1640) );
  XOR U2288 ( .A(n1711), .B(n1712), .Z(n1710) );
  XOR U2289 ( .A(key[1216]), .B(n203), .Z(n1709) );
  XOR U2290 ( .A(n1713), .B(n1714), .Z(out[31]) );
  XOR U2291 ( .A(n1715), .B(n1716), .Z(n1713) );
  XNOR U2292 ( .A(key[1183]), .B(n1717), .Z(n1716) );
  XNOR U2293 ( .A(n1718), .B(n1719), .Z(out[30]) );
  XNOR U2294 ( .A(key[1182]), .B(n1720), .Z(n1719) );
  XOR U2295 ( .A(key[1154]), .B(n1125), .Z(out[2]) );
  XNOR U2296 ( .A(n443), .B(n1721), .Z(n1125) );
  IV U2297 ( .A(n1510), .Z(n443) );
  XOR U2298 ( .A(n1722), .B(n1723), .Z(out[29]) );
  XNOR U2299 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U2300 ( .A(n1715), .B(n1726), .Z(n1725) );
  XNOR U2301 ( .A(n1728), .B(n1729), .Z(n1727) );
  NANDN U2302 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U2303 ( .A(n1733), .B(n1734), .Z(n1722) );
  XOR U2304 ( .A(key[1181]), .B(n1735), .Z(n1734) );
  ANDN U2305 ( .B(n1736), .A(n1737), .Z(n1733) );
  XNOR U2306 ( .A(n1738), .B(n1739), .Z(out[28]) );
  XNOR U2307 ( .A(key[1180]), .B(n1740), .Z(n1739) );
  XOR U2308 ( .A(n1741), .B(n1742), .Z(out[27]) );
  XNOR U2309 ( .A(n1743), .B(n1718), .Z(n1742) );
  XNOR U2310 ( .A(n1744), .B(n1745), .Z(n1718) );
  XNOR U2311 ( .A(n1746), .B(n1735), .Z(n1745) );
  ANDN U2312 ( .B(n1747), .A(n1748), .Z(n1735) );
  NOR U2313 ( .A(n1749), .B(n1750), .Z(n1746) );
  XNOR U2314 ( .A(n1751), .B(n1752), .Z(n1741) );
  XOR U2315 ( .A(key[1179]), .B(n1753), .Z(n1752) );
  XOR U2316 ( .A(key[1178]), .B(n1738), .Z(out[26]) );
  XNOR U2317 ( .A(n1717), .B(n1754), .Z(n1738) );
  IV U2318 ( .A(n1753), .Z(n1717) );
  XOR U2319 ( .A(n1755), .B(n1714), .Z(out[25]) );
  XNOR U2320 ( .A(n1744), .B(n1756), .Z(n1743) );
  XNOR U2321 ( .A(n1757), .B(n1758), .Z(n1756) );
  NANDN U2322 ( .A(n1759), .B(n1731), .Z(n1758) );
  XNOR U2323 ( .A(n1726), .B(n1760), .Z(n1744) );
  XNOR U2324 ( .A(n1761), .B(n1762), .Z(n1760) );
  NANDN U2325 ( .A(n1763), .B(n1764), .Z(n1762) );
  XOR U2326 ( .A(n1754), .B(n1751), .Z(n1720) );
  XNOR U2327 ( .A(n1726), .B(n1765), .Z(n1751) );
  XNOR U2328 ( .A(n1757), .B(n1766), .Z(n1765) );
  NANDN U2329 ( .A(n1767), .B(n1768), .Z(n1766) );
  OR U2330 ( .A(n1769), .B(n1770), .Z(n1757) );
  XOR U2331 ( .A(n1771), .B(n1761), .Z(n1726) );
  NANDN U2332 ( .A(n1772), .B(n1773), .Z(n1761) );
  ANDN U2333 ( .B(n1774), .A(n1775), .Z(n1771) );
  XOR U2334 ( .A(key[1177]), .B(n1753), .Z(n1755) );
  XOR U2335 ( .A(n1776), .B(n1777), .Z(n1753) );
  XNOR U2336 ( .A(n1778), .B(n1779), .Z(n1777) );
  NANDN U2337 ( .A(n1780), .B(n1736), .Z(n1779) );
  XNOR U2338 ( .A(n1724), .B(n1781), .Z(out[24]) );
  XOR U2339 ( .A(key[1176]), .B(n1754), .Z(n1781) );
  XNOR U2340 ( .A(n1776), .B(n1782), .Z(n1754) );
  XOR U2341 ( .A(n1783), .B(n1728), .Z(n1782) );
  OR U2342 ( .A(n1784), .B(n1769), .Z(n1728) );
  XNOR U2343 ( .A(n1731), .B(n1768), .Z(n1769) );
  ANDN U2344 ( .B(n1785), .A(n1786), .Z(n1783) );
  IV U2345 ( .A(n1740), .Z(n1724) );
  XOR U2346 ( .A(n1732), .B(n1787), .Z(n1740) );
  XOR U2347 ( .A(n1788), .B(n1778), .Z(n1787) );
  XNOR U2348 ( .A(n1750), .B(n1736), .Z(n1747) );
  NOR U2349 ( .A(n1790), .B(n1750), .Z(n1788) );
  XNOR U2350 ( .A(n1776), .B(n1791), .Z(n1732) );
  XNOR U2351 ( .A(n1792), .B(n1793), .Z(n1791) );
  NANDN U2352 ( .A(n1763), .B(n1794), .Z(n1793) );
  XOR U2353 ( .A(n1795), .B(n1792), .Z(n1776) );
  OR U2354 ( .A(n1772), .B(n1796), .Z(n1792) );
  XOR U2355 ( .A(n1797), .B(n1763), .Z(n1772) );
  XNOR U2356 ( .A(n1768), .B(n1736), .Z(n1763) );
  XOR U2357 ( .A(n1798), .B(n1799), .Z(n1736) );
  NANDN U2358 ( .A(n1800), .B(n1801), .Z(n1799) );
  IV U2359 ( .A(n1786), .Z(n1768) );
  XNOR U2360 ( .A(n1802), .B(n1803), .Z(n1786) );
  NANDN U2361 ( .A(n1800), .B(n1804), .Z(n1803) );
  ANDN U2362 ( .B(n1797), .A(n1805), .Z(n1795) );
  IV U2363 ( .A(n1775), .Z(n1797) );
  XOR U2364 ( .A(n1750), .B(n1731), .Z(n1775) );
  XNOR U2365 ( .A(n1806), .B(n1802), .Z(n1731) );
  NANDN U2366 ( .A(n1807), .B(n1808), .Z(n1802) );
  XOR U2367 ( .A(n1804), .B(n1809), .Z(n1808) );
  ANDN U2368 ( .B(n1809), .A(n1810), .Z(n1806) );
  XOR U2369 ( .A(n1811), .B(n1798), .Z(n1750) );
  NANDN U2370 ( .A(n1807), .B(n1812), .Z(n1798) );
  XOR U2371 ( .A(n1813), .B(n1801), .Z(n1812) );
  XNOR U2372 ( .A(n1814), .B(n1815), .Z(n1800) );
  XOR U2373 ( .A(n1816), .B(n1817), .Z(n1815) );
  XNOR U2374 ( .A(n1818), .B(n1819), .Z(n1814) );
  XNOR U2375 ( .A(n1820), .B(n1821), .Z(n1819) );
  ANDN U2376 ( .B(n1813), .A(n1817), .Z(n1820) );
  ANDN U2377 ( .B(n1813), .A(n1810), .Z(n1811) );
  XNOR U2378 ( .A(n1816), .B(n1822), .Z(n1810) );
  XOR U2379 ( .A(n1823), .B(n1821), .Z(n1822) );
  NAND U2380 ( .A(n1824), .B(n1825), .Z(n1821) );
  XNOR U2381 ( .A(n1818), .B(n1801), .Z(n1825) );
  IV U2382 ( .A(n1813), .Z(n1818) );
  XNOR U2383 ( .A(n1804), .B(n1817), .Z(n1824) );
  IV U2384 ( .A(n1809), .Z(n1817) );
  XOR U2385 ( .A(n1826), .B(n1827), .Z(n1809) );
  XNOR U2386 ( .A(n1828), .B(n1829), .Z(n1827) );
  XNOR U2387 ( .A(n1830), .B(n1831), .Z(n1826) );
  NOR U2388 ( .A(n1749), .B(n1790), .Z(n1830) );
  AND U2389 ( .A(n1801), .B(n1804), .Z(n1823) );
  XNOR U2390 ( .A(n1801), .B(n1804), .Z(n1816) );
  XNOR U2391 ( .A(n1832), .B(n1833), .Z(n1804) );
  XNOR U2392 ( .A(n1834), .B(n1829), .Z(n1833) );
  XOR U2393 ( .A(n1835), .B(n1836), .Z(n1832) );
  XNOR U2394 ( .A(n1837), .B(n1831), .Z(n1836) );
  OR U2395 ( .A(n1748), .B(n1789), .Z(n1831) );
  XNOR U2396 ( .A(n1790), .B(n1780), .Z(n1789) );
  XNOR U2397 ( .A(n1749), .B(n1737), .Z(n1748) );
  ANDN U2398 ( .B(n1838), .A(n1780), .Z(n1837) );
  XNOR U2399 ( .A(n1839), .B(n1840), .Z(n1801) );
  XNOR U2400 ( .A(n1829), .B(n1841), .Z(n1840) );
  XOR U2401 ( .A(n1759), .B(n1835), .Z(n1841) );
  XNOR U2402 ( .A(n1790), .B(n1842), .Z(n1829) );
  XNOR U2403 ( .A(n1843), .B(n1844), .Z(n1839) );
  XNOR U2404 ( .A(n1845), .B(n1846), .Z(n1844) );
  ANDN U2405 ( .B(n1785), .A(n1767), .Z(n1845) );
  XNOR U2406 ( .A(n1847), .B(n1848), .Z(n1813) );
  XNOR U2407 ( .A(n1834), .B(n1849), .Z(n1848) );
  XNOR U2408 ( .A(n1767), .B(n1828), .Z(n1849) );
  XOR U2409 ( .A(n1835), .B(n1850), .Z(n1828) );
  XNOR U2410 ( .A(n1851), .B(n1852), .Z(n1850) );
  NAND U2411 ( .A(n1794), .B(n1764), .Z(n1852) );
  XNOR U2412 ( .A(n1853), .B(n1851), .Z(n1835) );
  NANDN U2413 ( .A(n1796), .B(n1773), .Z(n1851) );
  XOR U2414 ( .A(n1774), .B(n1764), .Z(n1773) );
  XNOR U2415 ( .A(n1854), .B(n1737), .Z(n1764) );
  XOR U2416 ( .A(n1805), .B(n1794), .Z(n1796) );
  XOR U2417 ( .A(n1785), .B(n1855), .Z(n1794) );
  ANDN U2418 ( .B(n1774), .A(n1805), .Z(n1853) );
  XOR U2419 ( .A(n1843), .B(n1790), .Z(n1805) );
  XOR U2420 ( .A(n1856), .B(n1857), .Z(n1790) );
  XNOR U2421 ( .A(n1858), .B(n1859), .Z(n1857) );
  XOR U2422 ( .A(n1860), .B(n1842), .Z(n1774) );
  XOR U2423 ( .A(n1855), .B(n1838), .Z(n1834) );
  IV U2424 ( .A(n1737), .Z(n1838) );
  XOR U2425 ( .A(n1861), .B(n1862), .Z(n1737) );
  XNOR U2426 ( .A(n1863), .B(n1859), .Z(n1862) );
  IV U2427 ( .A(n1780), .Z(n1855) );
  XOR U2428 ( .A(n1859), .B(n1864), .Z(n1780) );
  XNOR U2429 ( .A(n1785), .B(n1865), .Z(n1847) );
  XNOR U2430 ( .A(n1866), .B(n1846), .Z(n1865) );
  OR U2431 ( .A(n1770), .B(n1784), .Z(n1846) );
  XNOR U2432 ( .A(n1843), .B(n1785), .Z(n1784) );
  XOR U2433 ( .A(n1759), .B(n1854), .Z(n1770) );
  IV U2434 ( .A(n1767), .Z(n1854) );
  XOR U2435 ( .A(n1842), .B(n1867), .Z(n1767) );
  XNOR U2436 ( .A(n1863), .B(n1856), .Z(n1867) );
  XOR U2437 ( .A(n1868), .B(n1869), .Z(n1856) );
  XNOR U2438 ( .A(n638), .B(n1870), .Z(n1869) );
  XOR U2439 ( .A(n1871), .B(n1872), .Z(n1868) );
  XNOR U2440 ( .A(key[1178]), .B(n1873), .Z(n1872) );
  IV U2441 ( .A(n1749), .Z(n1842) );
  XOR U2442 ( .A(n1861), .B(n1874), .Z(n1749) );
  XOR U2443 ( .A(n1859), .B(n1875), .Z(n1874) );
  ANDN U2444 ( .B(n1860), .A(n1730), .Z(n1866) );
  IV U2445 ( .A(n1759), .Z(n1860) );
  XOR U2446 ( .A(n1861), .B(n1876), .Z(n1759) );
  XOR U2447 ( .A(n1859), .B(n1877), .Z(n1876) );
  XOR U2448 ( .A(n1878), .B(n1879), .Z(n1859) );
  XNOR U2449 ( .A(n1250), .B(n1730), .Z(n1879) );
  IV U2450 ( .A(n1843), .Z(n1730) );
  XOR U2451 ( .A(n1880), .B(n1881), .Z(n1250) );
  XNOR U2452 ( .A(n612), .B(n1882), .Z(n1878) );
  XNOR U2453 ( .A(key[1182]), .B(n1883), .Z(n1882) );
  IV U2454 ( .A(n1864), .Z(n1861) );
  XOR U2455 ( .A(n1884), .B(n1885), .Z(n1864) );
  XOR U2456 ( .A(n1886), .B(n1258), .Z(n1885) );
  XNOR U2457 ( .A(n630), .B(n1887), .Z(n1884) );
  XOR U2458 ( .A(key[1181]), .B(n1888), .Z(n1887) );
  XOR U2459 ( .A(n1889), .B(n1890), .Z(n1785) );
  XNOR U2460 ( .A(n1877), .B(n1875), .Z(n1890) );
  XNOR U2461 ( .A(n1891), .B(n1892), .Z(n1875) );
  XOR U2462 ( .A(n1265), .B(n1893), .Z(n1892) );
  XOR U2463 ( .A(key[1183]), .B(n1894), .Z(n1891) );
  XNOR U2464 ( .A(n1895), .B(n1896), .Z(n1877) );
  XNOR U2465 ( .A(n1897), .B(n1271), .Z(n1896) );
  XOR U2466 ( .A(n1880), .B(n1898), .Z(n1271) );
  XNOR U2467 ( .A(n1899), .B(n1900), .Z(n1895) );
  XNOR U2468 ( .A(key[1180]), .B(n1275), .Z(n1900) );
  XOR U2469 ( .A(n1843), .B(n1858), .Z(n1889) );
  XOR U2470 ( .A(n1901), .B(n1902), .Z(n1858) );
  XNOR U2471 ( .A(n1863), .B(n1903), .Z(n1902) );
  XNOR U2472 ( .A(n1904), .B(n1279), .Z(n1903) );
  XNOR U2473 ( .A(n1268), .B(n597), .Z(n1279) );
  IV U2474 ( .A(n1880), .Z(n1268) );
  XOR U2475 ( .A(n1905), .B(n1906), .Z(n1863) );
  XOR U2476 ( .A(n650), .B(n1287), .Z(n1906) );
  XNOR U2477 ( .A(n1907), .B(n1908), .Z(n1905) );
  XOR U2478 ( .A(key[1177]), .B(n627), .Z(n1908) );
  XOR U2479 ( .A(n1243), .B(n1909), .Z(n1901) );
  XNOR U2480 ( .A(key[1179]), .B(n652), .Z(n1909) );
  XOR U2481 ( .A(n1910), .B(n1911), .Z(n1843) );
  XNOR U2482 ( .A(n639), .B(n608), .Z(n1911) );
  XOR U2483 ( .A(n1266), .B(n623), .Z(n608) );
  XOR U2484 ( .A(n1880), .B(n1912), .Z(n1910) );
  XOR U2485 ( .A(key[1176]), .B(n1913), .Z(n1912) );
  XOR U2486 ( .A(n1914), .B(n1915), .Z(out[23]) );
  XOR U2487 ( .A(n1916), .B(n1917), .Z(n1914) );
  XNOR U2488 ( .A(key[1175]), .B(n1918), .Z(n1917) );
  XNOR U2489 ( .A(n1919), .B(n1920), .Z(out[22]) );
  XNOR U2490 ( .A(key[1174]), .B(n1921), .Z(n1920) );
  XOR U2491 ( .A(n1922), .B(n1923), .Z(out[21]) );
  XNOR U2492 ( .A(n1924), .B(n1925), .Z(n1923) );
  XOR U2493 ( .A(n1916), .B(n1926), .Z(n1925) );
  XNOR U2494 ( .A(n1928), .B(n1929), .Z(n1927) );
  NANDN U2495 ( .A(n1930), .B(n1931), .Z(n1929) );
  XOR U2496 ( .A(n1933), .B(n1934), .Z(n1922) );
  XOR U2497 ( .A(key[1173]), .B(n1935), .Z(n1934) );
  ANDN U2498 ( .B(n1936), .A(n1937), .Z(n1933) );
  XNOR U2499 ( .A(n1938), .B(n1939), .Z(out[20]) );
  XNOR U2500 ( .A(key[1172]), .B(n1940), .Z(n1939) );
  XOR U2501 ( .A(n1941), .B(n440), .Z(out[1]) );
  XNOR U2502 ( .A(n1501), .B(n1942), .Z(n1500) );
  XNOR U2503 ( .A(n1943), .B(n1944), .Z(n1942) );
  NANDN U2504 ( .A(n1945), .B(n894), .Z(n1944) );
  XNOR U2505 ( .A(n889), .B(n1946), .Z(n1501) );
  XNOR U2506 ( .A(n1947), .B(n1948), .Z(n1946) );
  NANDN U2507 ( .A(n1949), .B(n1950), .Z(n1948) );
  XOR U2508 ( .A(n1721), .B(n1508), .Z(n665) );
  XNOR U2509 ( .A(n889), .B(n1951), .Z(n1508) );
  XNOR U2510 ( .A(n1943), .B(n1952), .Z(n1951) );
  NANDN U2511 ( .A(n1953), .B(n1954), .Z(n1952) );
  OR U2512 ( .A(n1955), .B(n1956), .Z(n1943) );
  XOR U2513 ( .A(n1957), .B(n1947), .Z(n889) );
  NANDN U2514 ( .A(n1958), .B(n1959), .Z(n1947) );
  ANDN U2515 ( .B(n1960), .A(n1961), .Z(n1957) );
  XOR U2516 ( .A(key[1153]), .B(n1510), .Z(n1941) );
  XOR U2517 ( .A(n1962), .B(n1963), .Z(n1510) );
  XNOR U2518 ( .A(n1964), .B(n1965), .Z(n1963) );
  NANDN U2519 ( .A(n1966), .B(n899), .Z(n1965) );
  XOR U2520 ( .A(n1967), .B(n1968), .Z(out[19]) );
  XNOR U2521 ( .A(n1969), .B(n1919), .Z(n1968) );
  XNOR U2522 ( .A(n1970), .B(n1971), .Z(n1919) );
  XNOR U2523 ( .A(n1972), .B(n1935), .Z(n1971) );
  ANDN U2524 ( .B(n1973), .A(n1974), .Z(n1935) );
  NOR U2525 ( .A(n1975), .B(n1976), .Z(n1972) );
  XNOR U2526 ( .A(n1977), .B(n1978), .Z(n1967) );
  XOR U2527 ( .A(key[1171]), .B(n1979), .Z(n1978) );
  XOR U2528 ( .A(key[1170]), .B(n1938), .Z(out[18]) );
  XNOR U2529 ( .A(n1918), .B(n1980), .Z(n1938) );
  IV U2530 ( .A(n1979), .Z(n1918) );
  XOR U2531 ( .A(n1981), .B(n1915), .Z(out[17]) );
  XNOR U2532 ( .A(n1970), .B(n1982), .Z(n1969) );
  XNOR U2533 ( .A(n1983), .B(n1984), .Z(n1982) );
  NANDN U2534 ( .A(n1985), .B(n1931), .Z(n1984) );
  XNOR U2535 ( .A(n1926), .B(n1986), .Z(n1970) );
  XNOR U2536 ( .A(n1987), .B(n1988), .Z(n1986) );
  NANDN U2537 ( .A(n1989), .B(n1990), .Z(n1988) );
  XOR U2538 ( .A(n1980), .B(n1977), .Z(n1921) );
  XNOR U2539 ( .A(n1926), .B(n1991), .Z(n1977) );
  XNOR U2540 ( .A(n1983), .B(n1992), .Z(n1991) );
  NANDN U2541 ( .A(n1993), .B(n1994), .Z(n1992) );
  OR U2542 ( .A(n1995), .B(n1996), .Z(n1983) );
  XOR U2543 ( .A(n1997), .B(n1987), .Z(n1926) );
  NANDN U2544 ( .A(n1998), .B(n1999), .Z(n1987) );
  ANDN U2545 ( .B(n2000), .A(n2001), .Z(n1997) );
  XOR U2546 ( .A(key[1169]), .B(n1979), .Z(n1981) );
  XOR U2547 ( .A(n2002), .B(n2003), .Z(n1979) );
  XNOR U2548 ( .A(n2004), .B(n2005), .Z(n2003) );
  NANDN U2549 ( .A(n2006), .B(n1936), .Z(n2005) );
  XNOR U2550 ( .A(n1924), .B(n2007), .Z(out[16]) );
  XOR U2551 ( .A(key[1168]), .B(n1980), .Z(n2007) );
  XNOR U2552 ( .A(n2002), .B(n2008), .Z(n1980) );
  XOR U2553 ( .A(n2009), .B(n1928), .Z(n2008) );
  OR U2554 ( .A(n2010), .B(n1995), .Z(n1928) );
  XNOR U2555 ( .A(n1931), .B(n1994), .Z(n1995) );
  ANDN U2556 ( .B(n1994), .A(n2011), .Z(n2009) );
  IV U2557 ( .A(n1940), .Z(n1924) );
  XOR U2558 ( .A(n1932), .B(n2012), .Z(n1940) );
  XOR U2559 ( .A(n2013), .B(n2004), .Z(n2012) );
  XNOR U2560 ( .A(n1976), .B(n1936), .Z(n1973) );
  NOR U2561 ( .A(n2015), .B(n1976), .Z(n2013) );
  XNOR U2562 ( .A(n2002), .B(n2016), .Z(n1932) );
  XNOR U2563 ( .A(n2017), .B(n2018), .Z(n2016) );
  NANDN U2564 ( .A(n1989), .B(n2019), .Z(n2018) );
  XOR U2565 ( .A(n2020), .B(n2017), .Z(n2002) );
  OR U2566 ( .A(n1998), .B(n2021), .Z(n2017) );
  XOR U2567 ( .A(n2022), .B(n1989), .Z(n1998) );
  XNOR U2568 ( .A(n1994), .B(n1936), .Z(n1989) );
  XOR U2569 ( .A(n2023), .B(n2024), .Z(n1936) );
  NANDN U2570 ( .A(n2025), .B(n2026), .Z(n2024) );
  XOR U2571 ( .A(n2027), .B(n2028), .Z(n1994) );
  NANDN U2572 ( .A(n2025), .B(n2029), .Z(n2028) );
  ANDN U2573 ( .B(n2022), .A(n2030), .Z(n2020) );
  IV U2574 ( .A(n2001), .Z(n2022) );
  XOR U2575 ( .A(n1976), .B(n1931), .Z(n2001) );
  XNOR U2576 ( .A(n2031), .B(n2027), .Z(n1931) );
  NANDN U2577 ( .A(n2032), .B(n2033), .Z(n2027) );
  XOR U2578 ( .A(n2029), .B(n2034), .Z(n2033) );
  ANDN U2579 ( .B(n2034), .A(n2035), .Z(n2031) );
  XOR U2580 ( .A(n2036), .B(n2023), .Z(n1976) );
  NANDN U2581 ( .A(n2032), .B(n2037), .Z(n2023) );
  XOR U2582 ( .A(n2038), .B(n2026), .Z(n2037) );
  XNOR U2583 ( .A(n2039), .B(n2040), .Z(n2025) );
  XOR U2584 ( .A(n2041), .B(n2042), .Z(n2040) );
  XNOR U2585 ( .A(n2043), .B(n2044), .Z(n2039) );
  XNOR U2586 ( .A(n2045), .B(n2046), .Z(n2044) );
  ANDN U2587 ( .B(n2038), .A(n2042), .Z(n2045) );
  ANDN U2588 ( .B(n2038), .A(n2035), .Z(n2036) );
  XNOR U2589 ( .A(n2041), .B(n2047), .Z(n2035) );
  XOR U2590 ( .A(n2048), .B(n2046), .Z(n2047) );
  NAND U2591 ( .A(n2049), .B(n2050), .Z(n2046) );
  XNOR U2592 ( .A(n2043), .B(n2026), .Z(n2050) );
  IV U2593 ( .A(n2038), .Z(n2043) );
  XNOR U2594 ( .A(n2029), .B(n2042), .Z(n2049) );
  IV U2595 ( .A(n2034), .Z(n2042) );
  XOR U2596 ( .A(n2051), .B(n2052), .Z(n2034) );
  XNOR U2597 ( .A(n2053), .B(n2054), .Z(n2052) );
  XNOR U2598 ( .A(n2055), .B(n2056), .Z(n2051) );
  NOR U2599 ( .A(n1975), .B(n2015), .Z(n2055) );
  AND U2600 ( .A(n2026), .B(n2029), .Z(n2048) );
  XNOR U2601 ( .A(n2026), .B(n2029), .Z(n2041) );
  XNOR U2602 ( .A(n2057), .B(n2058), .Z(n2029) );
  XNOR U2603 ( .A(n2059), .B(n2054), .Z(n2058) );
  XOR U2604 ( .A(n2060), .B(n2061), .Z(n2057) );
  XNOR U2605 ( .A(n2062), .B(n2056), .Z(n2061) );
  OR U2606 ( .A(n1974), .B(n2014), .Z(n2056) );
  XNOR U2607 ( .A(n2015), .B(n2006), .Z(n2014) );
  XNOR U2608 ( .A(n1975), .B(n1937), .Z(n1974) );
  ANDN U2609 ( .B(n2063), .A(n2006), .Z(n2062) );
  XNOR U2610 ( .A(n2064), .B(n2065), .Z(n2026) );
  XNOR U2611 ( .A(n2054), .B(n2066), .Z(n2065) );
  XOR U2612 ( .A(n1985), .B(n2060), .Z(n2066) );
  XNOR U2613 ( .A(n2015), .B(n2067), .Z(n2054) );
  XOR U2614 ( .A(n1930), .B(n2068), .Z(n2064) );
  XNOR U2615 ( .A(n2069), .B(n2070), .Z(n2068) );
  ANDN U2616 ( .B(n2071), .A(n2011), .Z(n2069) );
  XNOR U2617 ( .A(n2072), .B(n2073), .Z(n2038) );
  XNOR U2618 ( .A(n2059), .B(n2074), .Z(n2073) );
  XNOR U2619 ( .A(n1993), .B(n2053), .Z(n2074) );
  XOR U2620 ( .A(n2060), .B(n2075), .Z(n2053) );
  XNOR U2621 ( .A(n2076), .B(n2077), .Z(n2075) );
  NAND U2622 ( .A(n2019), .B(n1990), .Z(n2077) );
  XNOR U2623 ( .A(n2078), .B(n2076), .Z(n2060) );
  NANDN U2624 ( .A(n2021), .B(n1999), .Z(n2076) );
  XOR U2625 ( .A(n2000), .B(n1990), .Z(n1999) );
  XNOR U2626 ( .A(n2071), .B(n1937), .Z(n1990) );
  XOR U2627 ( .A(n2030), .B(n2019), .Z(n2021) );
  XNOR U2628 ( .A(n2011), .B(n2079), .Z(n2019) );
  ANDN U2629 ( .B(n2000), .A(n2030), .Z(n2078) );
  XNOR U2630 ( .A(n1930), .B(n2015), .Z(n2030) );
  XOR U2631 ( .A(n2080), .B(n2081), .Z(n2015) );
  XNOR U2632 ( .A(n2082), .B(n2083), .Z(n2081) );
  XOR U2633 ( .A(n2079), .B(n2063), .Z(n2059) );
  IV U2634 ( .A(n1937), .Z(n2063) );
  XOR U2635 ( .A(n2084), .B(n2085), .Z(n1937) );
  XOR U2636 ( .A(n2086), .B(n2083), .Z(n2085) );
  IV U2637 ( .A(n2006), .Z(n2079) );
  XOR U2638 ( .A(n2083), .B(n2087), .Z(n2006) );
  XNOR U2639 ( .A(n2088), .B(n2089), .Z(n2072) );
  XNOR U2640 ( .A(n2090), .B(n2070), .Z(n2089) );
  OR U2641 ( .A(n1996), .B(n2010), .Z(n2070) );
  XNOR U2642 ( .A(n1930), .B(n2011), .Z(n2010) );
  IV U2643 ( .A(n2088), .Z(n2011) );
  XOR U2644 ( .A(n1985), .B(n2071), .Z(n1996) );
  IV U2645 ( .A(n1993), .Z(n2071) );
  XOR U2646 ( .A(n2067), .B(n2091), .Z(n1993) );
  XNOR U2647 ( .A(n2092), .B(n2080), .Z(n2091) );
  XOR U2648 ( .A(n2093), .B(n2094), .Z(n2080) );
  XNOR U2649 ( .A(n836), .B(n831), .Z(n2094) );
  XOR U2650 ( .A(n846), .B(n1486), .Z(n836) );
  XOR U2651 ( .A(key[1266]), .B(n1488), .Z(n2093) );
  IV U2652 ( .A(n1975), .Z(n2067) );
  XOR U2653 ( .A(n2084), .B(n2095), .Z(n1975) );
  XOR U2654 ( .A(n2083), .B(n2096), .Z(n2095) );
  NOR U2655 ( .A(n1985), .B(n1930), .Z(n2090) );
  XOR U2656 ( .A(n2084), .B(n2097), .Z(n1985) );
  XOR U2657 ( .A(n2083), .B(n2098), .Z(n2097) );
  XOR U2658 ( .A(n2099), .B(n2100), .Z(n2083) );
  XNOR U2659 ( .A(n1930), .B(n2101), .Z(n2100) );
  XOR U2660 ( .A(n1454), .B(n2102), .Z(n2099) );
  XNOR U2661 ( .A(key[1270]), .B(n1464), .Z(n2102) );
  XOR U2662 ( .A(n826), .B(n2103), .Z(n1454) );
  XOR U2663 ( .A(n850), .B(n1460), .Z(n826) );
  IV U2664 ( .A(n2104), .Z(n1460) );
  IV U2665 ( .A(n2087), .Z(n2084) );
  XOR U2666 ( .A(n2105), .B(n2106), .Z(n2087) );
  XNOR U2667 ( .A(n2107), .B(n1461), .Z(n2106) );
  XOR U2668 ( .A(n827), .B(n1478), .Z(n1461) );
  XNOR U2669 ( .A(key[1269]), .B(n2108), .Z(n2105) );
  XOR U2670 ( .A(n2109), .B(n2110), .Z(n2088) );
  XNOR U2671 ( .A(n2098), .B(n2096), .Z(n2110) );
  XNOR U2672 ( .A(n2111), .B(n2112), .Z(n2096) );
  XNOR U2673 ( .A(n2103), .B(n1469), .Z(n2112) );
  XOR U2674 ( .A(n1457), .B(n2113), .Z(n1469) );
  XNOR U2675 ( .A(n856), .B(n2114), .Z(n2103) );
  XNOR U2676 ( .A(key[1271]), .B(n2115), .Z(n2111) );
  XNOR U2677 ( .A(n2116), .B(n2117), .Z(n2098) );
  XNOR U2678 ( .A(n1475), .B(n2118), .Z(n2117) );
  XOR U2679 ( .A(n811), .B(n1492), .Z(n1475) );
  XNOR U2680 ( .A(n1474), .B(n2119), .Z(n2116) );
  XOR U2681 ( .A(key[1268]), .B(n2120), .Z(n2119) );
  XNOR U2682 ( .A(n856), .B(n2107), .Z(n1474) );
  XNOR U2683 ( .A(n1930), .B(n2082), .Z(n2109) );
  XOR U2684 ( .A(n2121), .B(n2122), .Z(n2082) );
  XNOR U2685 ( .A(n2123), .B(n2124), .Z(n2122) );
  XNOR U2686 ( .A(n1481), .B(n2092), .Z(n2124) );
  IV U2687 ( .A(n2086), .Z(n2092) );
  XNOR U2688 ( .A(n2125), .B(n2126), .Z(n2086) );
  XNOR U2689 ( .A(n845), .B(n1495), .Z(n2126) );
  XNOR U2690 ( .A(key[1265]), .B(n857), .Z(n2125) );
  XNOR U2691 ( .A(n2127), .B(n1497), .Z(n857) );
  XNOR U2692 ( .A(n856), .B(n2120), .Z(n1481) );
  XNOR U2693 ( .A(n2128), .B(n2129), .Z(n2121) );
  XOR U2694 ( .A(key[1267]), .B(n1491), .Z(n2129) );
  XOR U2695 ( .A(n841), .B(n1447), .Z(n1491) );
  XNOR U2696 ( .A(n2130), .B(n2131), .Z(n1930) );
  XNOR U2697 ( .A(n837), .B(n1470), .Z(n2131) );
  XOR U2698 ( .A(key[1264]), .B(n2132), .Z(n2130) );
  XOR U2699 ( .A(n2133), .B(n2134), .Z(out[15]) );
  XNOR U2700 ( .A(n4), .B(n2135), .Z(n2134) );
  XNOR U2701 ( .A(n3), .B(n2136), .Z(n2133) );
  XOR U2702 ( .A(key[1167]), .B(n5), .Z(n2136) );
  XNOR U2703 ( .A(n2137), .B(n2138), .Z(out[14]) );
  XOR U2704 ( .A(key[1166]), .B(n3), .Z(n2138) );
  XOR U2705 ( .A(n63), .B(n2139), .Z(n3) );
  IV U2706 ( .A(n2140), .Z(n63) );
  XOR U2707 ( .A(n2141), .B(n2142), .Z(out[13]) );
  XNOR U2708 ( .A(n2135), .B(n2143), .Z(n2142) );
  XNOR U2709 ( .A(n2144), .B(n61), .Z(n2143) );
  XNOR U2710 ( .A(n2145), .B(n2146), .Z(n2135) );
  XNOR U2711 ( .A(n2147), .B(n2148), .Z(n2146) );
  NANDN U2712 ( .A(n2149), .B(n2150), .Z(n2148) );
  XOR U2713 ( .A(n2151), .B(n2152), .Z(n2141) );
  XOR U2714 ( .A(key[1165]), .B(n2153), .Z(n2152) );
  ANDN U2715 ( .B(n2154), .A(n2155), .Z(n2151) );
  XNOR U2716 ( .A(n2156), .B(n2157), .Z(out[12]) );
  XOR U2717 ( .A(key[1164]), .B(n61), .Z(n2157) );
  XNOR U2718 ( .A(n2145), .B(n2158), .Z(n61) );
  XOR U2719 ( .A(n2159), .B(n2160), .Z(n2158) );
  ANDN U2720 ( .B(n2161), .A(n2162), .Z(n2159) );
  XNOR U2721 ( .A(n2163), .B(n2164), .Z(n2145) );
  XNOR U2722 ( .A(n2165), .B(n2166), .Z(n2164) );
  NAND U2723 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U2724 ( .A(n2169), .B(n2170), .Z(out[127]) );
  XOR U2725 ( .A(n2171), .B(n2172), .Z(n2169) );
  XNOR U2726 ( .A(key[1279]), .B(n2173), .Z(n2172) );
  XNOR U2727 ( .A(n2174), .B(n2175), .Z(out[126]) );
  XNOR U2728 ( .A(key[1278]), .B(n2176), .Z(n2175) );
  XOR U2729 ( .A(n2177), .B(n2178), .Z(out[125]) );
  XNOR U2730 ( .A(n2179), .B(n2180), .Z(n2178) );
  XOR U2731 ( .A(n2171), .B(n2181), .Z(n2180) );
  XNOR U2732 ( .A(n2183), .B(n2184), .Z(n2182) );
  NANDN U2733 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U2734 ( .A(n2188), .B(n2189), .Z(n2177) );
  XOR U2735 ( .A(key[1277]), .B(n2190), .Z(n2189) );
  ANDN U2736 ( .B(n2191), .A(n2192), .Z(n2188) );
  XNOR U2737 ( .A(n2193), .B(n2194), .Z(out[124]) );
  XNOR U2738 ( .A(key[1276]), .B(n2195), .Z(n2194) );
  XOR U2739 ( .A(n2196), .B(n2197), .Z(out[123]) );
  XNOR U2740 ( .A(n2198), .B(n2174), .Z(n2197) );
  XNOR U2741 ( .A(n2199), .B(n2200), .Z(n2174) );
  XNOR U2742 ( .A(n2201), .B(n2190), .Z(n2200) );
  ANDN U2743 ( .B(n2202), .A(n2203), .Z(n2190) );
  NOR U2744 ( .A(n2204), .B(n2205), .Z(n2201) );
  XNOR U2745 ( .A(n2206), .B(n2207), .Z(n2196) );
  XOR U2746 ( .A(key[1275]), .B(n2208), .Z(n2207) );
  XOR U2747 ( .A(key[1274]), .B(n2193), .Z(out[122]) );
  XNOR U2748 ( .A(n2173), .B(n2209), .Z(n2193) );
  IV U2749 ( .A(n2208), .Z(n2173) );
  XOR U2750 ( .A(n2210), .B(n2170), .Z(out[121]) );
  XNOR U2751 ( .A(n2199), .B(n2211), .Z(n2198) );
  XNOR U2752 ( .A(n2212), .B(n2213), .Z(n2211) );
  NANDN U2753 ( .A(n2214), .B(n2186), .Z(n2213) );
  XNOR U2754 ( .A(n2181), .B(n2215), .Z(n2199) );
  XNOR U2755 ( .A(n2216), .B(n2217), .Z(n2215) );
  NANDN U2756 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U2757 ( .A(n2209), .B(n2206), .Z(n2176) );
  XNOR U2758 ( .A(n2181), .B(n2220), .Z(n2206) );
  XNOR U2759 ( .A(n2212), .B(n2221), .Z(n2220) );
  NANDN U2760 ( .A(n2222), .B(n2223), .Z(n2221) );
  OR U2761 ( .A(n2224), .B(n2225), .Z(n2212) );
  XOR U2762 ( .A(n2226), .B(n2216), .Z(n2181) );
  NANDN U2763 ( .A(n2227), .B(n2228), .Z(n2216) );
  ANDN U2764 ( .B(n2229), .A(n2230), .Z(n2226) );
  XOR U2765 ( .A(key[1273]), .B(n2208), .Z(n2210) );
  XOR U2766 ( .A(n2231), .B(n2232), .Z(n2208) );
  XNOR U2767 ( .A(n2233), .B(n2234), .Z(n2232) );
  NANDN U2768 ( .A(n2235), .B(n2191), .Z(n2234) );
  XNOR U2769 ( .A(n2179), .B(n2236), .Z(out[120]) );
  XOR U2770 ( .A(key[1272]), .B(n2209), .Z(n2236) );
  XNOR U2771 ( .A(n2231), .B(n2237), .Z(n2209) );
  XOR U2772 ( .A(n2238), .B(n2183), .Z(n2237) );
  OR U2773 ( .A(n2239), .B(n2224), .Z(n2183) );
  XNOR U2774 ( .A(n2186), .B(n2223), .Z(n2224) );
  ANDN U2775 ( .B(n2240), .A(n2241), .Z(n2238) );
  IV U2776 ( .A(n2195), .Z(n2179) );
  XOR U2777 ( .A(n2187), .B(n2242), .Z(n2195) );
  XOR U2778 ( .A(n2243), .B(n2233), .Z(n2242) );
  XNOR U2779 ( .A(n2205), .B(n2191), .Z(n2202) );
  NOR U2780 ( .A(n2245), .B(n2205), .Z(n2243) );
  XNOR U2781 ( .A(n2231), .B(n2246), .Z(n2187) );
  XNOR U2782 ( .A(n2247), .B(n2248), .Z(n2246) );
  NANDN U2783 ( .A(n2218), .B(n2249), .Z(n2248) );
  XOR U2784 ( .A(n2250), .B(n2247), .Z(n2231) );
  OR U2785 ( .A(n2227), .B(n2251), .Z(n2247) );
  XOR U2786 ( .A(n2252), .B(n2218), .Z(n2227) );
  XNOR U2787 ( .A(n2223), .B(n2191), .Z(n2218) );
  XOR U2788 ( .A(n2253), .B(n2254), .Z(n2191) );
  NANDN U2789 ( .A(n2255), .B(n2256), .Z(n2254) );
  IV U2790 ( .A(n2241), .Z(n2223) );
  XNOR U2791 ( .A(n2257), .B(n2258), .Z(n2241) );
  NANDN U2792 ( .A(n2255), .B(n2259), .Z(n2258) );
  ANDN U2793 ( .B(n2252), .A(n2260), .Z(n2250) );
  IV U2794 ( .A(n2230), .Z(n2252) );
  XOR U2795 ( .A(n2205), .B(n2186), .Z(n2230) );
  XNOR U2796 ( .A(n2261), .B(n2257), .Z(n2186) );
  NANDN U2797 ( .A(n2262), .B(n2263), .Z(n2257) );
  XOR U2798 ( .A(n2259), .B(n2264), .Z(n2263) );
  ANDN U2799 ( .B(n2264), .A(n2265), .Z(n2261) );
  XOR U2800 ( .A(n2266), .B(n2253), .Z(n2205) );
  NANDN U2801 ( .A(n2262), .B(n2267), .Z(n2253) );
  XOR U2802 ( .A(n2268), .B(n2256), .Z(n2267) );
  XNOR U2803 ( .A(n2269), .B(n2270), .Z(n2255) );
  XOR U2804 ( .A(n2271), .B(n2272), .Z(n2270) );
  XNOR U2805 ( .A(n2273), .B(n2274), .Z(n2269) );
  XNOR U2806 ( .A(n2275), .B(n2276), .Z(n2274) );
  ANDN U2807 ( .B(n2268), .A(n2272), .Z(n2275) );
  ANDN U2808 ( .B(n2268), .A(n2265), .Z(n2266) );
  XNOR U2809 ( .A(n2271), .B(n2277), .Z(n2265) );
  XOR U2810 ( .A(n2278), .B(n2276), .Z(n2277) );
  NAND U2811 ( .A(n2279), .B(n2280), .Z(n2276) );
  XNOR U2812 ( .A(n2273), .B(n2256), .Z(n2280) );
  IV U2813 ( .A(n2268), .Z(n2273) );
  XNOR U2814 ( .A(n2259), .B(n2272), .Z(n2279) );
  IV U2815 ( .A(n2264), .Z(n2272) );
  XOR U2816 ( .A(n2281), .B(n2282), .Z(n2264) );
  XNOR U2817 ( .A(n2283), .B(n2284), .Z(n2282) );
  XNOR U2818 ( .A(n2285), .B(n2286), .Z(n2281) );
  NOR U2819 ( .A(n2204), .B(n2245), .Z(n2285) );
  AND U2820 ( .A(n2256), .B(n2259), .Z(n2278) );
  XNOR U2821 ( .A(n2256), .B(n2259), .Z(n2271) );
  XNOR U2822 ( .A(n2287), .B(n2288), .Z(n2259) );
  XNOR U2823 ( .A(n2289), .B(n2284), .Z(n2288) );
  XOR U2824 ( .A(n2290), .B(n2291), .Z(n2287) );
  XNOR U2825 ( .A(n2292), .B(n2286), .Z(n2291) );
  OR U2826 ( .A(n2203), .B(n2244), .Z(n2286) );
  XNOR U2827 ( .A(n2245), .B(n2235), .Z(n2244) );
  XNOR U2828 ( .A(n2204), .B(n2192), .Z(n2203) );
  ANDN U2829 ( .B(n2293), .A(n2235), .Z(n2292) );
  XNOR U2830 ( .A(n2294), .B(n2295), .Z(n2256) );
  XNOR U2831 ( .A(n2284), .B(n2296), .Z(n2295) );
  XOR U2832 ( .A(n2214), .B(n2290), .Z(n2296) );
  XNOR U2833 ( .A(n2245), .B(n2297), .Z(n2284) );
  XNOR U2834 ( .A(n2298), .B(n2299), .Z(n2294) );
  XNOR U2835 ( .A(n2300), .B(n2301), .Z(n2299) );
  ANDN U2836 ( .B(n2240), .A(n2222), .Z(n2300) );
  XNOR U2837 ( .A(n2302), .B(n2303), .Z(n2268) );
  XNOR U2838 ( .A(n2289), .B(n2304), .Z(n2303) );
  XNOR U2839 ( .A(n2222), .B(n2283), .Z(n2304) );
  XOR U2840 ( .A(n2290), .B(n2305), .Z(n2283) );
  XNOR U2841 ( .A(n2306), .B(n2307), .Z(n2305) );
  NAND U2842 ( .A(n2249), .B(n2219), .Z(n2307) );
  XNOR U2843 ( .A(n2308), .B(n2306), .Z(n2290) );
  NANDN U2844 ( .A(n2251), .B(n2228), .Z(n2306) );
  XOR U2845 ( .A(n2229), .B(n2219), .Z(n2228) );
  XNOR U2846 ( .A(n2309), .B(n2192), .Z(n2219) );
  XOR U2847 ( .A(n2260), .B(n2249), .Z(n2251) );
  XOR U2848 ( .A(n2240), .B(n2310), .Z(n2249) );
  ANDN U2849 ( .B(n2229), .A(n2260), .Z(n2308) );
  XOR U2850 ( .A(n2298), .B(n2245), .Z(n2260) );
  XOR U2851 ( .A(n2311), .B(n2312), .Z(n2245) );
  XNOR U2852 ( .A(n2313), .B(n2314), .Z(n2312) );
  XOR U2853 ( .A(n2315), .B(n2297), .Z(n2229) );
  XOR U2854 ( .A(n2310), .B(n2293), .Z(n2289) );
  IV U2855 ( .A(n2192), .Z(n2293) );
  XOR U2856 ( .A(n2316), .B(n2317), .Z(n2192) );
  XNOR U2857 ( .A(n2318), .B(n2314), .Z(n2317) );
  IV U2858 ( .A(n2235), .Z(n2310) );
  XOR U2859 ( .A(n2314), .B(n2319), .Z(n2235) );
  XNOR U2860 ( .A(n2240), .B(n2320), .Z(n2302) );
  XNOR U2861 ( .A(n2321), .B(n2301), .Z(n2320) );
  OR U2862 ( .A(n2225), .B(n2239), .Z(n2301) );
  XNOR U2863 ( .A(n2298), .B(n2240), .Z(n2239) );
  XOR U2864 ( .A(n2214), .B(n2309), .Z(n2225) );
  IV U2865 ( .A(n2222), .Z(n2309) );
  XOR U2866 ( .A(n2297), .B(n2322), .Z(n2222) );
  XNOR U2867 ( .A(n2318), .B(n2311), .Z(n2322) );
  XOR U2868 ( .A(n2323), .B(n2324), .Z(n2311) );
  XNOR U2869 ( .A(n1486), .B(n1483), .Z(n2324) );
  XOR U2870 ( .A(n845), .B(n2325), .Z(n2323) );
  XNOR U2871 ( .A(key[1274]), .B(n841), .Z(n2325) );
  XOR U2872 ( .A(n2326), .B(n2327), .Z(n841) );
  XOR U2873 ( .A(n2328), .B(n2329), .Z(n2327) );
  XNOR U2874 ( .A(n2330), .B(n2331), .Z(n2326) );
  XOR U2875 ( .A(n1445), .B(n1488), .Z(n845) );
  IV U2876 ( .A(n2204), .Z(n2297) );
  XOR U2877 ( .A(n2316), .B(n2332), .Z(n2204) );
  XOR U2878 ( .A(n2314), .B(n2333), .Z(n2332) );
  ANDN U2879 ( .B(n2315), .A(n2185), .Z(n2321) );
  IV U2880 ( .A(n2214), .Z(n2315) );
  XOR U2881 ( .A(n2316), .B(n2334), .Z(n2214) );
  XOR U2882 ( .A(n2314), .B(n2335), .Z(n2334) );
  XOR U2883 ( .A(n2336), .B(n2337), .Z(n2314) );
  XNOR U2884 ( .A(n2101), .B(n2185), .Z(n2337) );
  IV U2885 ( .A(n2298), .Z(n2185) );
  XOR U2886 ( .A(n2338), .B(n2339), .Z(n2101) );
  XOR U2887 ( .A(n2104), .B(n2340), .Z(n2336) );
  XOR U2888 ( .A(key[1278]), .B(n849), .Z(n2340) );
  XOR U2889 ( .A(n820), .B(n2108), .Z(n849) );
  XNOR U2890 ( .A(n1455), .B(n1464), .Z(n2108) );
  XOR U2891 ( .A(n2341), .B(n2342), .Z(n1464) );
  XOR U2892 ( .A(n2343), .B(n2113), .Z(n820) );
  XNOR U2893 ( .A(n2344), .B(n2345), .Z(n2113) );
  XNOR U2894 ( .A(n2346), .B(n2347), .Z(n2345) );
  XOR U2895 ( .A(n2330), .B(n2348), .Z(n2344) );
  XOR U2896 ( .A(n2349), .B(n2350), .Z(n2104) );
  IV U2897 ( .A(n2319), .Z(n2316) );
  XOR U2898 ( .A(n2351), .B(n2352), .Z(n2319) );
  XOR U2899 ( .A(n1478), .B(n825), .Z(n2352) );
  XNOR U2900 ( .A(n1462), .B(n2107), .Z(n825) );
  XNOR U2901 ( .A(n2353), .B(n2354), .Z(n2107) );
  XNOR U2902 ( .A(n2355), .B(n2356), .Z(n2354) );
  XNOR U2903 ( .A(n2357), .B(n2358), .Z(n2353) );
  XOR U2904 ( .A(n2359), .B(n2360), .Z(n2358) );
  ANDN U2905 ( .B(n2361), .A(n2362), .Z(n2360) );
  XNOR U2906 ( .A(n2363), .B(n2364), .Z(n1478) );
  XNOR U2907 ( .A(n2365), .B(n2366), .Z(n2364) );
  XNOR U2908 ( .A(n2367), .B(n2368), .Z(n2363) );
  XOR U2909 ( .A(n2369), .B(n2370), .Z(n2368) );
  ANDN U2910 ( .B(n2371), .A(n2372), .Z(n2370) );
  XOR U2911 ( .A(n850), .B(n2373), .Z(n2351) );
  XNOR U2912 ( .A(key[1277]), .B(n1455), .Z(n2373) );
  XOR U2913 ( .A(n2374), .B(n2375), .Z(n1455) );
  XNOR U2914 ( .A(n2346), .B(n2329), .Z(n850) );
  XOR U2915 ( .A(n2376), .B(n2377), .Z(n2329) );
  XNOR U2916 ( .A(n2378), .B(n2379), .Z(n2377) );
  NOR U2917 ( .A(n2380), .B(n2381), .Z(n2378) );
  XOR U2918 ( .A(n2382), .B(n2383), .Z(n2240) );
  XNOR U2919 ( .A(n2335), .B(n2333), .Z(n2383) );
  XNOR U2920 ( .A(n2384), .B(n2385), .Z(n2333) );
  XNOR U2921 ( .A(n1457), .B(n821), .Z(n2385) );
  XNOR U2922 ( .A(n2339), .B(n2114), .Z(n821) );
  XNOR U2923 ( .A(n2386), .B(n2387), .Z(n2114) );
  XNOR U2924 ( .A(n2388), .B(n2356), .Z(n2387) );
  XNOR U2925 ( .A(n2389), .B(n2390), .Z(n2356) );
  XNOR U2926 ( .A(n2391), .B(n2392), .Z(n2390) );
  NANDN U2927 ( .A(n2393), .B(n2394), .Z(n2392) );
  XNOR U2928 ( .A(n2395), .B(n2341), .Z(n2386) );
  IV U2929 ( .A(n1471), .Z(n2339) );
  XOR U2930 ( .A(n2396), .B(n2397), .Z(n1471) );
  XNOR U2931 ( .A(n2374), .B(n2398), .Z(n2397) );
  XOR U2932 ( .A(n2399), .B(n2400), .Z(n2396) );
  XOR U2933 ( .A(n2401), .B(n2402), .Z(n1457) );
  XNOR U2934 ( .A(n2349), .B(n2366), .Z(n2402) );
  XNOR U2935 ( .A(n2403), .B(n2404), .Z(n2366) );
  XNOR U2936 ( .A(n2405), .B(n2406), .Z(n2404) );
  NANDN U2937 ( .A(n2407), .B(n2408), .Z(n2406) );
  IV U2938 ( .A(n2409), .Z(n2349) );
  XNOR U2939 ( .A(n2410), .B(n2411), .Z(n2401) );
  XNOR U2940 ( .A(key[1279]), .B(n855), .Z(n2384) );
  XNOR U2941 ( .A(n2132), .B(n2338), .Z(n855) );
  XNOR U2942 ( .A(n2412), .B(n2413), .Z(n2335) );
  XOR U2943 ( .A(n808), .B(n2118), .Z(n2413) );
  XOR U2944 ( .A(n2338), .B(n1462), .Z(n2118) );
  XNOR U2945 ( .A(n2414), .B(n2415), .Z(n1462) );
  XNOR U2946 ( .A(n2416), .B(n2398), .Z(n2415) );
  XNOR U2947 ( .A(n2417), .B(n2418), .Z(n2398) );
  XNOR U2948 ( .A(n2419), .B(n2420), .Z(n2418) );
  NANDN U2949 ( .A(n2421), .B(n2422), .Z(n2420) );
  XNOR U2950 ( .A(n2423), .B(n2424), .Z(n2414) );
  XOR U2951 ( .A(n2425), .B(n2426), .Z(n2424) );
  ANDN U2952 ( .B(n2427), .A(n2428), .Z(n2426) );
  XOR U2953 ( .A(n1476), .B(n2120), .Z(n808) );
  XNOR U2954 ( .A(n2357), .B(n1488), .Z(n2120) );
  XOR U2955 ( .A(n2429), .B(n2430), .Z(n1488) );
  XNOR U2956 ( .A(n809), .B(n2431), .Z(n2412) );
  XNOR U2957 ( .A(key[1276]), .B(n1492), .Z(n2431) );
  XOR U2958 ( .A(n2365), .B(n1486), .Z(n1492) );
  XNOR U2959 ( .A(n2432), .B(n2433), .Z(n1486) );
  XOR U2960 ( .A(n2343), .B(n827), .Z(n809) );
  XNOR U2961 ( .A(n2434), .B(n2435), .Z(n827) );
  XNOR U2962 ( .A(n2436), .B(n2347), .Z(n2435) );
  XNOR U2963 ( .A(n2437), .B(n2438), .Z(n2347) );
  XNOR U2964 ( .A(n2439), .B(n2440), .Z(n2438) );
  NANDN U2965 ( .A(n2441), .B(n2442), .Z(n2440) );
  XNOR U2966 ( .A(n2443), .B(n2444), .Z(n2434) );
  XOR U2967 ( .A(n2379), .B(n2445), .Z(n2444) );
  ANDN U2968 ( .B(n2446), .A(n2447), .Z(n2445) );
  NOR U2969 ( .A(n2448), .B(n2449), .Z(n2379) );
  XOR U2970 ( .A(n2298), .B(n2313), .Z(n2382) );
  XOR U2971 ( .A(n2450), .B(n2451), .Z(n2313) );
  XNOR U2972 ( .A(n2318), .B(n2452), .Z(n2451) );
  XOR U2973 ( .A(n831), .B(n2123), .Z(n2452) );
  XNOR U2974 ( .A(n2115), .B(n1476), .Z(n2123) );
  XOR U2975 ( .A(n2423), .B(n1445), .Z(n1476) );
  XOR U2976 ( .A(n1444), .B(n1483), .Z(n831) );
  XNOR U2977 ( .A(n2453), .B(n2454), .Z(n1483) );
  XOR U2978 ( .A(n2455), .B(n2375), .Z(n2454) );
  XOR U2979 ( .A(n2456), .B(n2457), .Z(n2375) );
  XNOR U2980 ( .A(n2458), .B(n2425), .Z(n2457) );
  ANDN U2981 ( .B(n2459), .A(n2460), .Z(n2425) );
  ANDN U2982 ( .B(n2461), .A(n2462), .Z(n2458) );
  IV U2983 ( .A(n2128), .Z(n1444) );
  XOR U2984 ( .A(n2463), .B(n2464), .Z(n2128) );
  XOR U2985 ( .A(n2388), .B(n2342), .Z(n2464) );
  XOR U2986 ( .A(n2465), .B(n2466), .Z(n2342) );
  XNOR U2987 ( .A(n2467), .B(n2359), .Z(n2466) );
  ANDN U2988 ( .B(n2468), .A(n2469), .Z(n2359) );
  ANDN U2989 ( .B(n2470), .A(n2471), .Z(n2467) );
  XOR U2990 ( .A(n2430), .B(n2472), .Z(n2463) );
  XOR U2991 ( .A(n2473), .B(n2474), .Z(n2318) );
  XNOR U2992 ( .A(n1445), .B(n837), .Z(n2474) );
  XOR U2993 ( .A(n1487), .B(n1495), .Z(n837) );
  XOR U2994 ( .A(n2388), .B(n2475), .Z(n1495) );
  XNOR U2995 ( .A(n2430), .B(n2341), .Z(n2475) );
  XNOR U2996 ( .A(n2355), .B(n2476), .Z(n2472) );
  XNOR U2997 ( .A(n2477), .B(n2478), .Z(n2476) );
  NANDN U2998 ( .A(n2479), .B(n2480), .Z(n2478) );
  IV U2999 ( .A(n2395), .Z(n2430) );
  XOR U3000 ( .A(n2481), .B(n2482), .Z(n2395) );
  XOR U3001 ( .A(n2483), .B(n2484), .Z(n2482) );
  NANDN U3002 ( .A(n2485), .B(n2361), .Z(n2484) );
  XNOR U3003 ( .A(n2465), .B(n2486), .Z(n2388) );
  XNOR U3004 ( .A(n2477), .B(n2487), .Z(n2486) );
  NANDN U3005 ( .A(n2488), .B(n2394), .Z(n2487) );
  OR U3006 ( .A(n2489), .B(n2490), .Z(n2477) );
  XNOR U3007 ( .A(n2355), .B(n2491), .Z(n2465) );
  XNOR U3008 ( .A(n2492), .B(n2493), .Z(n2491) );
  NANDN U3009 ( .A(n2494), .B(n2495), .Z(n2493) );
  XOR U3010 ( .A(n2496), .B(n2492), .Z(n2355) );
  NANDN U3011 ( .A(n2497), .B(n2498), .Z(n2492) );
  ANDN U3012 ( .B(n2499), .A(n2500), .Z(n2496) );
  IV U3013 ( .A(n2501), .Z(n1487) );
  XNOR U3014 ( .A(n2502), .B(n2399), .Z(n1445) );
  XOR U3015 ( .A(n846), .B(n2503), .Z(n2473) );
  XOR U3016 ( .A(key[1273]), .B(n1497), .Z(n2503) );
  XNOR U3017 ( .A(n2409), .B(n2504), .Z(n1497) );
  XOR U3018 ( .A(n2410), .B(n2411), .Z(n2504) );
  IV U3019 ( .A(n2432), .Z(n2410) );
  XOR U3020 ( .A(n2433), .B(n2505), .Z(n2409) );
  XNOR U3021 ( .A(n839), .B(n2506), .Z(n2450) );
  XNOR U3022 ( .A(key[1275]), .B(n1447), .Z(n2506) );
  XOR U3023 ( .A(n2507), .B(n2508), .Z(n1447) );
  XNOR U3024 ( .A(n2505), .B(n2350), .Z(n2508) );
  XNOR U3025 ( .A(n2509), .B(n2510), .Z(n2350) );
  XNOR U3026 ( .A(n2511), .B(n2369), .Z(n2510) );
  ANDN U3027 ( .B(n2512), .A(n2513), .Z(n2369) );
  ANDN U3028 ( .B(n2514), .A(n2515), .Z(n2511) );
  XNOR U3029 ( .A(n2367), .B(n2516), .Z(n2505) );
  XNOR U3030 ( .A(n2517), .B(n2518), .Z(n2516) );
  NANDN U3031 ( .A(n2519), .B(n2520), .Z(n2518) );
  XOR U3032 ( .A(n2432), .B(n2411), .Z(n2507) );
  XNOR U3033 ( .A(n2517), .B(n2522), .Z(n2521) );
  NANDN U3034 ( .A(n2523), .B(n2408), .Z(n2522) );
  OR U3035 ( .A(n2524), .B(n2525), .Z(n2517) );
  XNOR U3036 ( .A(n2367), .B(n2526), .Z(n2509) );
  XNOR U3037 ( .A(n2527), .B(n2528), .Z(n2526) );
  NANDN U3038 ( .A(n2529), .B(n2530), .Z(n2528) );
  XOR U3039 ( .A(n2531), .B(n2527), .Z(n2367) );
  NANDN U3040 ( .A(n2532), .B(n2533), .Z(n2527) );
  ANDN U3041 ( .B(n2534), .A(n2535), .Z(n2531) );
  XOR U3042 ( .A(n2536), .B(n2537), .Z(n2432) );
  XOR U3043 ( .A(n2538), .B(n2539), .Z(n2537) );
  NANDN U3044 ( .A(n2540), .B(n2371), .Z(n2539) );
  XOR U3045 ( .A(n2132), .B(n811), .Z(n839) );
  XOR U3046 ( .A(n2436), .B(n846), .Z(n811) );
  XOR U3047 ( .A(n2331), .B(n2541), .Z(n846) );
  IV U3048 ( .A(n2343), .Z(n2132) );
  XOR U3049 ( .A(n2541), .B(n2436), .Z(n2343) );
  XNOR U3050 ( .A(n2437), .B(n2542), .Z(n2436) );
  XOR U3051 ( .A(n2543), .B(n2544), .Z(n2542) );
  NOR U3052 ( .A(n2545), .B(n2381), .Z(n2543) );
  XNOR U3053 ( .A(n2546), .B(n2547), .Z(n2437) );
  XNOR U3054 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U3055 ( .A(n2550), .B(n2551), .Z(n2549) );
  XOR U3056 ( .A(n2552), .B(n2553), .Z(n2298) );
  XOR U3057 ( .A(n2501), .B(n1470), .Z(n2553) );
  XOR U3058 ( .A(n856), .B(n822), .Z(n1470) );
  XOR U3059 ( .A(n2433), .B(n2365), .Z(n822) );
  XNOR U3060 ( .A(n2403), .B(n2554), .Z(n2365) );
  XNOR U3061 ( .A(n2555), .B(n2538), .Z(n2554) );
  XOR U3062 ( .A(n2557), .B(n2371), .Z(n2512) );
  ANDN U3063 ( .B(n2558), .A(n2515), .Z(n2555) );
  IV U3064 ( .A(n2557), .Z(n2515) );
  XNOR U3065 ( .A(n2536), .B(n2559), .Z(n2403) );
  XNOR U3066 ( .A(n2560), .B(n2561), .Z(n2559) );
  NANDN U3067 ( .A(n2529), .B(n2562), .Z(n2561) );
  XNOR U3068 ( .A(n2536), .B(n2563), .Z(n2433) );
  XOR U3069 ( .A(n2564), .B(n2405), .Z(n2563) );
  OR U3070 ( .A(n2565), .B(n2524), .Z(n2405) );
  XNOR U3071 ( .A(n2408), .B(n2520), .Z(n2524) );
  ANDN U3072 ( .B(n2566), .A(n2567), .Z(n2564) );
  XOR U3073 ( .A(n2568), .B(n2560), .Z(n2536) );
  OR U3074 ( .A(n2532), .B(n2569), .Z(n2560) );
  XNOR U3075 ( .A(n2535), .B(n2529), .Z(n2532) );
  XNOR U3076 ( .A(n2520), .B(n2371), .Z(n2529) );
  XOR U3077 ( .A(n2570), .B(n2571), .Z(n2371) );
  NANDN U3078 ( .A(n2572), .B(n2573), .Z(n2571) );
  IV U3079 ( .A(n2567), .Z(n2520) );
  XNOR U3080 ( .A(n2574), .B(n2575), .Z(n2567) );
  NANDN U3081 ( .A(n2572), .B(n2576), .Z(n2575) );
  NOR U3082 ( .A(n2535), .B(n2577), .Z(n2568) );
  XNOR U3083 ( .A(n2557), .B(n2408), .Z(n2535) );
  XNOR U3084 ( .A(n2578), .B(n2574), .Z(n2408) );
  NANDN U3085 ( .A(n2579), .B(n2580), .Z(n2574) );
  XOR U3086 ( .A(n2576), .B(n2581), .Z(n2580) );
  ANDN U3087 ( .B(n2581), .A(n2582), .Z(n2578) );
  XNOR U3088 ( .A(n2583), .B(n2570), .Z(n2557) );
  NANDN U3089 ( .A(n2579), .B(n2584), .Z(n2570) );
  XOR U3090 ( .A(n2585), .B(n2573), .Z(n2584) );
  XNOR U3091 ( .A(n2586), .B(n2587), .Z(n2572) );
  XOR U3092 ( .A(n2588), .B(n2589), .Z(n2587) );
  XNOR U3093 ( .A(n2590), .B(n2591), .Z(n2586) );
  XNOR U3094 ( .A(n2592), .B(n2593), .Z(n2591) );
  ANDN U3095 ( .B(n2585), .A(n2589), .Z(n2592) );
  ANDN U3096 ( .B(n2585), .A(n2582), .Z(n2583) );
  XNOR U3097 ( .A(n2588), .B(n2594), .Z(n2582) );
  XOR U3098 ( .A(n2595), .B(n2593), .Z(n2594) );
  NAND U3099 ( .A(n2596), .B(n2597), .Z(n2593) );
  XNOR U3100 ( .A(n2590), .B(n2573), .Z(n2597) );
  IV U3101 ( .A(n2585), .Z(n2590) );
  XNOR U3102 ( .A(n2576), .B(n2589), .Z(n2596) );
  IV U3103 ( .A(n2581), .Z(n2589) );
  XOR U3104 ( .A(n2598), .B(n2599), .Z(n2581) );
  XNOR U3105 ( .A(n2600), .B(n2601), .Z(n2599) );
  XNOR U3106 ( .A(n2602), .B(n2603), .Z(n2598) );
  ANDN U3107 ( .B(n2558), .A(n2604), .Z(n2602) );
  AND U3108 ( .A(n2573), .B(n2576), .Z(n2595) );
  XNOR U3109 ( .A(n2573), .B(n2576), .Z(n2588) );
  XNOR U3110 ( .A(n2605), .B(n2606), .Z(n2576) );
  XNOR U3111 ( .A(n2607), .B(n2601), .Z(n2606) );
  XOR U3112 ( .A(n2608), .B(n2609), .Z(n2605) );
  XNOR U3113 ( .A(n2610), .B(n2603), .Z(n2609) );
  OR U3114 ( .A(n2513), .B(n2556), .Z(n2603) );
  XNOR U3115 ( .A(n2558), .B(n2611), .Z(n2556) );
  XNOR U3116 ( .A(n2604), .B(n2372), .Z(n2513) );
  ANDN U3117 ( .B(n2612), .A(n2540), .Z(n2610) );
  XNOR U3118 ( .A(n2613), .B(n2614), .Z(n2573) );
  XNOR U3119 ( .A(n2601), .B(n2615), .Z(n2614) );
  XOR U3120 ( .A(n2523), .B(n2608), .Z(n2615) );
  XNOR U3121 ( .A(n2558), .B(n2604), .Z(n2601) );
  XNOR U3122 ( .A(n2616), .B(n2617), .Z(n2613) );
  XNOR U3123 ( .A(n2618), .B(n2619), .Z(n2617) );
  ANDN U3124 ( .B(n2566), .A(n2519), .Z(n2618) );
  XNOR U3125 ( .A(n2620), .B(n2621), .Z(n2585) );
  XNOR U3126 ( .A(n2607), .B(n2622), .Z(n2621) );
  XNOR U3127 ( .A(n2519), .B(n2600), .Z(n2622) );
  XOR U3128 ( .A(n2608), .B(n2623), .Z(n2600) );
  XNOR U3129 ( .A(n2624), .B(n2625), .Z(n2623) );
  NAND U3130 ( .A(n2562), .B(n2530), .Z(n2625) );
  XNOR U3131 ( .A(n2626), .B(n2624), .Z(n2608) );
  NANDN U3132 ( .A(n2569), .B(n2533), .Z(n2624) );
  XOR U3133 ( .A(n2534), .B(n2530), .Z(n2533) );
  XNOR U3134 ( .A(n2627), .B(n2372), .Z(n2530) );
  XOR U3135 ( .A(n2577), .B(n2562), .Z(n2569) );
  XOR U3136 ( .A(n2566), .B(n2611), .Z(n2562) );
  ANDN U3137 ( .B(n2534), .A(n2577), .Z(n2626) );
  XNOR U3138 ( .A(n2616), .B(n2558), .Z(n2577) );
  XNOR U3139 ( .A(n2628), .B(n2629), .Z(n2558) );
  XNOR U3140 ( .A(n2630), .B(n2631), .Z(n2629) );
  XOR U3141 ( .A(n2632), .B(n2514), .Z(n2534) );
  XOR U3142 ( .A(n2611), .B(n2612), .Z(n2607) );
  IV U3143 ( .A(n2372), .Z(n2612) );
  XOR U3144 ( .A(n2633), .B(n2634), .Z(n2372) );
  XNOR U3145 ( .A(n2635), .B(n2631), .Z(n2634) );
  IV U3146 ( .A(n2540), .Z(n2611) );
  XOR U3147 ( .A(n2631), .B(n2636), .Z(n2540) );
  XNOR U3148 ( .A(n2566), .B(n2637), .Z(n2620) );
  XNOR U3149 ( .A(n2638), .B(n2619), .Z(n2637) );
  OR U3150 ( .A(n2525), .B(n2565), .Z(n2619) );
  XNOR U3151 ( .A(n2616), .B(n2566), .Z(n2565) );
  XOR U3152 ( .A(n2523), .B(n2627), .Z(n2525) );
  IV U3153 ( .A(n2519), .Z(n2627) );
  XOR U3154 ( .A(n2514), .B(n2639), .Z(n2519) );
  XNOR U3155 ( .A(n2635), .B(n2628), .Z(n2639) );
  XOR U3156 ( .A(n2640), .B(n2641), .Z(n2628) );
  XNOR U3157 ( .A(n2642), .B(n2643), .Z(n2641) );
  XOR U3158 ( .A(key[1026]), .B(n2644), .Z(n2640) );
  IV U3159 ( .A(n2604), .Z(n2514) );
  XOR U3160 ( .A(n2633), .B(n2645), .Z(n2604) );
  XOR U3161 ( .A(n2631), .B(n2646), .Z(n2645) );
  ANDN U3162 ( .B(n2632), .A(n2407), .Z(n2638) );
  IV U3163 ( .A(n2523), .Z(n2632) );
  XOR U3164 ( .A(n2633), .B(n2647), .Z(n2523) );
  XOR U3165 ( .A(n2631), .B(n2648), .Z(n2647) );
  XOR U3166 ( .A(n2649), .B(n2650), .Z(n2631) );
  XNOR U3167 ( .A(n2651), .B(n2407), .Z(n2650) );
  IV U3168 ( .A(n2616), .Z(n2407) );
  XOR U3169 ( .A(n2652), .B(n2653), .Z(n2649) );
  XNOR U3170 ( .A(key[1030]), .B(n2654), .Z(n2653) );
  IV U3171 ( .A(n2636), .Z(n2633) );
  XOR U3172 ( .A(n2655), .B(n2656), .Z(n2636) );
  XNOR U3173 ( .A(n2657), .B(n2658), .Z(n2656) );
  XNOR U3174 ( .A(key[1029]), .B(n2659), .Z(n2655) );
  XOR U3175 ( .A(n2660), .B(n2661), .Z(n2566) );
  XNOR U3176 ( .A(n2648), .B(n2646), .Z(n2661) );
  XNOR U3177 ( .A(n2662), .B(n2663), .Z(n2646) );
  XOR U3178 ( .A(n2664), .B(n2665), .Z(n2663) );
  XNOR U3179 ( .A(key[1031]), .B(n2666), .Z(n2662) );
  XNOR U3180 ( .A(n2667), .B(n2668), .Z(n2648) );
  XNOR U3181 ( .A(n2669), .B(n2670), .Z(n2667) );
  XOR U3182 ( .A(key[1028]), .B(n2671), .Z(n2670) );
  XOR U3183 ( .A(n2616), .B(n2630), .Z(n2660) );
  XOR U3184 ( .A(n2672), .B(n2673), .Z(n2630) );
  XNOR U3185 ( .A(n2635), .B(n2674), .Z(n2673) );
  XOR U3186 ( .A(n2675), .B(n2676), .Z(n2674) );
  XOR U3187 ( .A(n2677), .B(n2678), .Z(n2635) );
  XNOR U3188 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR U3189 ( .A(key[1025]), .B(n2681), .Z(n2677) );
  XNOR U3190 ( .A(n2682), .B(n2683), .Z(n2672) );
  XNOR U3191 ( .A(key[1027]), .B(n2684), .Z(n2683) );
  XOR U3192 ( .A(n2685), .B(n2686), .Z(n2616) );
  XOR U3193 ( .A(n2687), .B(n2688), .Z(n2686) );
  XOR U3194 ( .A(key[1024]), .B(n2689), .Z(n2685) );
  XOR U3195 ( .A(n2429), .B(n2357), .Z(n856) );
  XNOR U3196 ( .A(n2389), .B(n2690), .Z(n2357) );
  XNOR U3197 ( .A(n2691), .B(n2483), .Z(n2690) );
  XOR U3198 ( .A(n2693), .B(n2361), .Z(n2468) );
  ANDN U3199 ( .B(n2694), .A(n2471), .Z(n2691) );
  IV U3200 ( .A(n2693), .Z(n2471) );
  XNOR U3201 ( .A(n2481), .B(n2695), .Z(n2389) );
  XNOR U3202 ( .A(n2696), .B(n2697), .Z(n2695) );
  NANDN U3203 ( .A(n2494), .B(n2698), .Z(n2697) );
  XNOR U3204 ( .A(n2481), .B(n2699), .Z(n2429) );
  XOR U3205 ( .A(n2700), .B(n2391), .Z(n2699) );
  OR U3206 ( .A(n2701), .B(n2489), .Z(n2391) );
  XNOR U3207 ( .A(n2394), .B(n2480), .Z(n2489) );
  ANDN U3208 ( .B(n2702), .A(n2703), .Z(n2700) );
  XOR U3209 ( .A(n2704), .B(n2696), .Z(n2481) );
  OR U3210 ( .A(n2497), .B(n2705), .Z(n2696) );
  XNOR U3211 ( .A(n2500), .B(n2494), .Z(n2497) );
  XNOR U3212 ( .A(n2480), .B(n2361), .Z(n2494) );
  XOR U3213 ( .A(n2706), .B(n2707), .Z(n2361) );
  NANDN U3214 ( .A(n2708), .B(n2709), .Z(n2707) );
  IV U3215 ( .A(n2703), .Z(n2480) );
  XNOR U3216 ( .A(n2710), .B(n2711), .Z(n2703) );
  NANDN U3217 ( .A(n2708), .B(n2712), .Z(n2711) );
  NOR U3218 ( .A(n2500), .B(n2713), .Z(n2704) );
  XNOR U3219 ( .A(n2693), .B(n2394), .Z(n2500) );
  XNOR U3220 ( .A(n2714), .B(n2710), .Z(n2394) );
  NANDN U3221 ( .A(n2715), .B(n2716), .Z(n2710) );
  XOR U3222 ( .A(n2712), .B(n2717), .Z(n2716) );
  ANDN U3223 ( .B(n2717), .A(n2718), .Z(n2714) );
  XNOR U3224 ( .A(n2719), .B(n2706), .Z(n2693) );
  NANDN U3225 ( .A(n2715), .B(n2720), .Z(n2706) );
  XOR U3226 ( .A(n2721), .B(n2709), .Z(n2720) );
  XNOR U3227 ( .A(n2722), .B(n2723), .Z(n2708) );
  XOR U3228 ( .A(n2724), .B(n2725), .Z(n2723) );
  XNOR U3229 ( .A(n2726), .B(n2727), .Z(n2722) );
  XNOR U3230 ( .A(n2728), .B(n2729), .Z(n2727) );
  ANDN U3231 ( .B(n2721), .A(n2725), .Z(n2728) );
  ANDN U3232 ( .B(n2721), .A(n2718), .Z(n2719) );
  XNOR U3233 ( .A(n2724), .B(n2730), .Z(n2718) );
  XOR U3234 ( .A(n2731), .B(n2729), .Z(n2730) );
  NAND U3235 ( .A(n2732), .B(n2733), .Z(n2729) );
  XNOR U3236 ( .A(n2726), .B(n2709), .Z(n2733) );
  IV U3237 ( .A(n2721), .Z(n2726) );
  XNOR U3238 ( .A(n2712), .B(n2725), .Z(n2732) );
  IV U3239 ( .A(n2717), .Z(n2725) );
  XOR U3240 ( .A(n2734), .B(n2735), .Z(n2717) );
  XNOR U3241 ( .A(n2736), .B(n2737), .Z(n2735) );
  XNOR U3242 ( .A(n2738), .B(n2739), .Z(n2734) );
  ANDN U3243 ( .B(n2694), .A(n2740), .Z(n2738) );
  AND U3244 ( .A(n2709), .B(n2712), .Z(n2731) );
  XNOR U3245 ( .A(n2709), .B(n2712), .Z(n2724) );
  XNOR U3246 ( .A(n2741), .B(n2742), .Z(n2712) );
  XNOR U3247 ( .A(n2743), .B(n2737), .Z(n2742) );
  XOR U3248 ( .A(n2744), .B(n2745), .Z(n2741) );
  XNOR U3249 ( .A(n2746), .B(n2739), .Z(n2745) );
  OR U3250 ( .A(n2469), .B(n2692), .Z(n2739) );
  XNOR U3251 ( .A(n2694), .B(n2747), .Z(n2692) );
  XNOR U3252 ( .A(n2740), .B(n2362), .Z(n2469) );
  ANDN U3253 ( .B(n2748), .A(n2485), .Z(n2746) );
  XNOR U3254 ( .A(n2749), .B(n2750), .Z(n2709) );
  XNOR U3255 ( .A(n2737), .B(n2751), .Z(n2750) );
  XOR U3256 ( .A(n2488), .B(n2744), .Z(n2751) );
  XNOR U3257 ( .A(n2694), .B(n2740), .Z(n2737) );
  XNOR U3258 ( .A(n2752), .B(n2753), .Z(n2749) );
  XNOR U3259 ( .A(n2754), .B(n2755), .Z(n2753) );
  ANDN U3260 ( .B(n2702), .A(n2479), .Z(n2754) );
  XNOR U3261 ( .A(n2756), .B(n2757), .Z(n2721) );
  XNOR U3262 ( .A(n2743), .B(n2758), .Z(n2757) );
  XNOR U3263 ( .A(n2479), .B(n2736), .Z(n2758) );
  XOR U3264 ( .A(n2744), .B(n2759), .Z(n2736) );
  XNOR U3265 ( .A(n2760), .B(n2761), .Z(n2759) );
  NAND U3266 ( .A(n2698), .B(n2495), .Z(n2761) );
  XNOR U3267 ( .A(n2762), .B(n2760), .Z(n2744) );
  NANDN U3268 ( .A(n2705), .B(n2498), .Z(n2760) );
  XOR U3269 ( .A(n2499), .B(n2495), .Z(n2498) );
  XNOR U3270 ( .A(n2763), .B(n2362), .Z(n2495) );
  XOR U3271 ( .A(n2713), .B(n2698), .Z(n2705) );
  XOR U3272 ( .A(n2702), .B(n2747), .Z(n2698) );
  ANDN U3273 ( .B(n2499), .A(n2713), .Z(n2762) );
  XNOR U3274 ( .A(n2752), .B(n2694), .Z(n2713) );
  XNOR U3275 ( .A(n2764), .B(n2765), .Z(n2694) );
  XNOR U3276 ( .A(n2766), .B(n2767), .Z(n2765) );
  XOR U3277 ( .A(n2768), .B(n2470), .Z(n2499) );
  XOR U3278 ( .A(n2747), .B(n2748), .Z(n2743) );
  IV U3279 ( .A(n2362), .Z(n2748) );
  XOR U3280 ( .A(n2769), .B(n2770), .Z(n2362) );
  XNOR U3281 ( .A(n2771), .B(n2767), .Z(n2770) );
  IV U3282 ( .A(n2485), .Z(n2747) );
  XOR U3283 ( .A(n2767), .B(n2772), .Z(n2485) );
  XNOR U3284 ( .A(n2702), .B(n2773), .Z(n2756) );
  XNOR U3285 ( .A(n2774), .B(n2755), .Z(n2773) );
  OR U3286 ( .A(n2490), .B(n2701), .Z(n2755) );
  XNOR U3287 ( .A(n2752), .B(n2702), .Z(n2701) );
  XOR U3288 ( .A(n2488), .B(n2763), .Z(n2490) );
  IV U3289 ( .A(n2479), .Z(n2763) );
  XOR U3290 ( .A(n2470), .B(n2775), .Z(n2479) );
  XNOR U3291 ( .A(n2771), .B(n2764), .Z(n2775) );
  XOR U3292 ( .A(n2776), .B(n2777), .Z(n2764) );
  XOR U3293 ( .A(n2778), .B(n2779), .Z(n2777) );
  XNOR U3294 ( .A(n2780), .B(n2781), .Z(n2776) );
  XNOR U3295 ( .A(key[1066]), .B(n2782), .Z(n2781) );
  IV U3296 ( .A(n2740), .Z(n2470) );
  XOR U3297 ( .A(n2769), .B(n2783), .Z(n2740) );
  XOR U3298 ( .A(n2767), .B(n2784), .Z(n2783) );
  ANDN U3299 ( .B(n2768), .A(n2393), .Z(n2774) );
  IV U3300 ( .A(n2488), .Z(n2768) );
  XOR U3301 ( .A(n2769), .B(n2785), .Z(n2488) );
  XOR U3302 ( .A(n2767), .B(n2786), .Z(n2785) );
  XOR U3303 ( .A(n2787), .B(n2788), .Z(n2767) );
  XOR U3304 ( .A(n2789), .B(n2393), .Z(n2788) );
  IV U3305 ( .A(n2752), .Z(n2393) );
  XNOR U3306 ( .A(n2790), .B(n2791), .Z(n2787) );
  XNOR U3307 ( .A(key[1070]), .B(n2792), .Z(n2791) );
  IV U3308 ( .A(n2772), .Z(n2769) );
  XOR U3309 ( .A(n2793), .B(n2794), .Z(n2772) );
  XOR U3310 ( .A(n2795), .B(n2796), .Z(n2794) );
  XNOR U3311 ( .A(n2797), .B(n2798), .Z(n2793) );
  XNOR U3312 ( .A(key[1069]), .B(n2799), .Z(n2798) );
  XOR U3313 ( .A(n2800), .B(n2801), .Z(n2702) );
  XNOR U3314 ( .A(n2786), .B(n2784), .Z(n2801) );
  XNOR U3315 ( .A(n2802), .B(n2803), .Z(n2784) );
  XOR U3316 ( .A(n2804), .B(n2805), .Z(n2803) );
  XOR U3317 ( .A(key[1071]), .B(n2806), .Z(n2802) );
  XNOR U3318 ( .A(n2807), .B(n2808), .Z(n2786) );
  XNOR U3319 ( .A(n2809), .B(n2810), .Z(n2808) );
  XNOR U3320 ( .A(n2811), .B(n2812), .Z(n2807) );
  XOR U3321 ( .A(key[1068]), .B(n2813), .Z(n2812) );
  XOR U3322 ( .A(n2752), .B(n2766), .Z(n2800) );
  XOR U3323 ( .A(n2814), .B(n2815), .Z(n2766) );
  XNOR U3324 ( .A(n2771), .B(n2816), .Z(n2815) );
  XOR U3325 ( .A(n2817), .B(n2818), .Z(n2816) );
  XOR U3326 ( .A(n2819), .B(n2820), .Z(n2771) );
  XNOR U3327 ( .A(n2821), .B(n2822), .Z(n2820) );
  XNOR U3328 ( .A(n2823), .B(n2824), .Z(n2819) );
  XOR U3329 ( .A(key[1065]), .B(n2825), .Z(n2824) );
  XNOR U3330 ( .A(n2826), .B(n2827), .Z(n2814) );
  XOR U3331 ( .A(key[1067]), .B(n2828), .Z(n2827) );
  XOR U3332 ( .A(n2829), .B(n2830), .Z(n2752) );
  XNOR U3333 ( .A(n2831), .B(n2832), .Z(n2830) );
  XOR U3334 ( .A(n2833), .B(n2834), .Z(n2829) );
  XOR U3335 ( .A(key[1064]), .B(n2835), .Z(n2834) );
  XNOR U3336 ( .A(n2374), .B(n2836), .Z(n2501) );
  XNOR U3337 ( .A(n2399), .B(n2400), .Z(n2836) );
  XOR U3338 ( .A(n2456), .B(n2837), .Z(n2400) );
  XNOR U3339 ( .A(n2838), .B(n2839), .Z(n2837) );
  NANDN U3340 ( .A(n2840), .B(n2422), .Z(n2839) );
  XNOR U3341 ( .A(n2416), .B(n2841), .Z(n2456) );
  XNOR U3342 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U3343 ( .A(n2844), .B(n2845), .Z(n2843) );
  XOR U3344 ( .A(n2846), .B(n2847), .Z(n2399) );
  XOR U3345 ( .A(n2848), .B(n2849), .Z(n2847) );
  NANDN U3346 ( .A(n2850), .B(n2427), .Z(n2849) );
  XOR U3347 ( .A(n2851), .B(n2455), .Z(n2374) );
  XNOR U3348 ( .A(n2416), .B(n2852), .Z(n2455) );
  XNOR U3349 ( .A(n2838), .B(n2853), .Z(n2852) );
  NANDN U3350 ( .A(n2854), .B(n2855), .Z(n2853) );
  OR U3351 ( .A(n2856), .B(n2857), .Z(n2838) );
  XOR U3352 ( .A(n2858), .B(n2842), .Z(n2416) );
  NANDN U3353 ( .A(n2859), .B(n2860), .Z(n2842) );
  ANDN U3354 ( .B(n2861), .A(n2862), .Z(n2858) );
  XOR U3355 ( .A(n2338), .B(n2863), .Z(n2552) );
  XOR U3356 ( .A(key[1272]), .B(n2127), .Z(n2863) );
  IV U3357 ( .A(n838), .Z(n2127) );
  XNOR U3358 ( .A(n2346), .B(n2864), .Z(n838) );
  XNOR U3359 ( .A(n2330), .B(n2348), .Z(n2864) );
  IV U3360 ( .A(n2331), .Z(n2348) );
  XOR U3361 ( .A(n2546), .B(n2865), .Z(n2331) );
  XNOR U3362 ( .A(n2544), .B(n2866), .Z(n2865) );
  NANDN U3363 ( .A(n2867), .B(n2446), .Z(n2866) );
  OR U3364 ( .A(n2868), .B(n2448), .Z(n2544) );
  XOR U3365 ( .A(n2381), .B(n2446), .Z(n2448) );
  XNOR U3366 ( .A(n2376), .B(n2869), .Z(n2330) );
  XNOR U3367 ( .A(n2870), .B(n2871), .Z(n2869) );
  NAND U3368 ( .A(n2872), .B(n2442), .Z(n2871) );
  XNOR U3369 ( .A(n2443), .B(n2873), .Z(n2376) );
  XNOR U3370 ( .A(n2874), .B(n2875), .Z(n2873) );
  NANDN U3371 ( .A(n2876), .B(n2877), .Z(n2875) );
  XOR U3372 ( .A(n2541), .B(n2328), .Z(n2346) );
  XNOR U3373 ( .A(n2443), .B(n2878), .Z(n2328) );
  XNOR U3374 ( .A(n2870), .B(n2879), .Z(n2878) );
  NANDN U3375 ( .A(n2880), .B(n2881), .Z(n2879) );
  OR U3376 ( .A(n2882), .B(n2883), .Z(n2870) );
  XOR U3377 ( .A(n2884), .B(n2874), .Z(n2443) );
  OR U3378 ( .A(n2885), .B(n2886), .Z(n2874) );
  ANDN U3379 ( .B(n2887), .A(n2888), .Z(n2884) );
  XOR U3380 ( .A(n2546), .B(n2889), .Z(n2541) );
  XOR U3381 ( .A(n2890), .B(n2439), .Z(n2889) );
  OR U3382 ( .A(n2891), .B(n2882), .Z(n2439) );
  XNOR U3383 ( .A(n2442), .B(n2881), .Z(n2882) );
  ANDN U3384 ( .B(n2881), .A(n2892), .Z(n2890) );
  XOR U3385 ( .A(n2893), .B(n2548), .Z(n2546) );
  OR U3386 ( .A(n2885), .B(n2894), .Z(n2548) );
  XNOR U3387 ( .A(n2887), .B(n2877), .Z(n2885) );
  IV U3388 ( .A(n2550), .Z(n2877) );
  XNOR U3389 ( .A(n2881), .B(n2446), .Z(n2550) );
  XOR U3390 ( .A(n2895), .B(n2896), .Z(n2446) );
  NANDN U3391 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR U3392 ( .A(n2899), .B(n2900), .Z(n2881) );
  NANDN U3393 ( .A(n2897), .B(n2901), .Z(n2900) );
  AND U3394 ( .A(n2902), .B(n2887), .Z(n2893) );
  XNOR U3395 ( .A(n2381), .B(n2442), .Z(n2887) );
  XNOR U3396 ( .A(n2903), .B(n2899), .Z(n2442) );
  NANDN U3397 ( .A(n2904), .B(n2905), .Z(n2899) );
  XOR U3398 ( .A(n2901), .B(n2906), .Z(n2905) );
  ANDN U3399 ( .B(n2906), .A(n2907), .Z(n2903) );
  NANDN U3400 ( .A(n2904), .B(n2909), .Z(n2895) );
  XOR U3401 ( .A(n2910), .B(n2898), .Z(n2909) );
  XNOR U3402 ( .A(n2911), .B(n2912), .Z(n2897) );
  XOR U3403 ( .A(n2913), .B(n2914), .Z(n2912) );
  XNOR U3404 ( .A(n2915), .B(n2916), .Z(n2911) );
  XNOR U3405 ( .A(n2917), .B(n2918), .Z(n2916) );
  ANDN U3406 ( .B(n2910), .A(n2914), .Z(n2917) );
  ANDN U3407 ( .B(n2910), .A(n2907), .Z(n2908) );
  XNOR U3408 ( .A(n2913), .B(n2919), .Z(n2907) );
  XOR U3409 ( .A(n2920), .B(n2918), .Z(n2919) );
  NAND U3410 ( .A(n2921), .B(n2922), .Z(n2918) );
  XNOR U3411 ( .A(n2915), .B(n2898), .Z(n2922) );
  IV U3412 ( .A(n2910), .Z(n2915) );
  XNOR U3413 ( .A(n2901), .B(n2914), .Z(n2921) );
  IV U3414 ( .A(n2906), .Z(n2914) );
  XOR U3415 ( .A(n2923), .B(n2924), .Z(n2906) );
  XNOR U3416 ( .A(n2925), .B(n2926), .Z(n2924) );
  XNOR U3417 ( .A(n2927), .B(n2928), .Z(n2923) );
  ANDN U3418 ( .B(n2929), .A(n2545), .Z(n2927) );
  AND U3419 ( .A(n2898), .B(n2901), .Z(n2920) );
  XNOR U3420 ( .A(n2898), .B(n2901), .Z(n2913) );
  XNOR U3421 ( .A(n2930), .B(n2931), .Z(n2901) );
  XNOR U3422 ( .A(n2932), .B(n2926), .Z(n2931) );
  XOR U3423 ( .A(n2933), .B(n2934), .Z(n2930) );
  XNOR U3424 ( .A(n2935), .B(n2928), .Z(n2934) );
  OR U3425 ( .A(n2449), .B(n2868), .Z(n2928) );
  XNOR U3426 ( .A(n2936), .B(n2967), .Z(n2868) );
  XNOR U3427 ( .A(n2380), .B(n2447), .Z(n2449) );
  ANDN U3428 ( .B(n2937), .A(n2867), .Z(n2935) );
  XNOR U3429 ( .A(n2938), .B(n2939), .Z(n2898) );
  XNOR U3430 ( .A(n2926), .B(n2940), .Z(n2939) );
  XNOR U3431 ( .A(n2872), .B(n2933), .Z(n2940) );
  XNOR U3432 ( .A(n2380), .B(n2936), .Z(n2926) );
  XNOR U3433 ( .A(n2941), .B(n2942), .Z(n2938) );
  XNOR U3434 ( .A(n2943), .B(n2944), .Z(n2942) );
  ANDN U3435 ( .B(n2945), .A(n2892), .Z(n2943) );
  XNOR U3436 ( .A(n2946), .B(n2947), .Z(n2910) );
  XNOR U3437 ( .A(n2932), .B(n2948), .Z(n2947) );
  XNOR U3438 ( .A(n2949), .B(n2925), .Z(n2948) );
  XOR U3439 ( .A(n2933), .B(n2950), .Z(n2925) );
  XNOR U3440 ( .A(n2951), .B(n2952), .Z(n2950) );
  NANDN U3441 ( .A(n2876), .B(n2551), .Z(n2952) );
  XNOR U3442 ( .A(n2953), .B(n2951), .Z(n2933) );
  OR U3443 ( .A(n2894), .B(n2886), .Z(n2951) );
  XOR U3444 ( .A(n2954), .B(n2876), .Z(n2886) );
  XNOR U3445 ( .A(n2937), .B(n2945), .Z(n2876) );
  IV U3446 ( .A(n2447), .Z(n2937) );
  XNOR U3447 ( .A(n2902), .B(n2551), .Z(n2894) );
  XNOR U3448 ( .A(n2892), .B(n2967), .Z(n2551) );
  IV U3449 ( .A(n2949), .Z(n2892) );
  ANDN U3450 ( .B(n2902), .A(n2888), .Z(n2953) );
  IV U3451 ( .A(n2954), .Z(n2888) );
  XOR U3452 ( .A(n2929), .B(n2872), .Z(n2954) );
  XOR U3453 ( .A(n2447), .B(n2867), .Z(n2932) );
  XOR U3454 ( .A(n2955), .B(n2956), .Z(n2867) );
  XOR U3455 ( .A(n2957), .B(n2958), .Z(n2447) );
  XOR U3456 ( .A(n2959), .B(n2956), .Z(n2958) );
  XNOR U3457 ( .A(n2880), .B(n2960), .Z(n2946) );
  XNOR U3458 ( .A(n2961), .B(n2944), .Z(n2960) );
  OR U3459 ( .A(n2883), .B(n2891), .Z(n2944) );
  XNOR U3460 ( .A(n2941), .B(n2949), .Z(n2891) );
  XOR U3461 ( .A(n2962), .B(n2963), .Z(n2949) );
  XNOR U3462 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR U3463 ( .A(n2941), .B(n2966), .Z(n2962) );
  XNOR U3464 ( .A(n2872), .B(n2945), .Z(n2883) );
  IV U3465 ( .A(n2880), .Z(n2945) );
  ANDN U3466 ( .B(n2872), .A(n2441), .Z(n2961) );
  XOR U3467 ( .A(n2964), .B(n2967), .Z(n2872) );
  XOR U3468 ( .A(n2968), .B(n2969), .Z(n2964) );
  XOR U3469 ( .A(n2970), .B(n2971), .Z(n2969) );
  XNOR U3470 ( .A(n2972), .B(n2973), .Z(n2968) );
  XNOR U3471 ( .A(key[1148]), .B(n2974), .Z(n2973) );
  XNOR U3472 ( .A(n2975), .B(n2976), .Z(n2880) );
  XOR U3473 ( .A(n2380), .B(n2957), .Z(n2976) );
  IV U3474 ( .A(n2929), .Z(n2380) );
  XOR U3475 ( .A(n2966), .B(n2967), .Z(n2929) );
  XNOR U3476 ( .A(n2955), .B(n2956), .Z(n2967) );
  IV U3477 ( .A(n2959), .Z(n2955) );
  XNOR U3478 ( .A(n2977), .B(n2978), .Z(n2959) );
  XOR U3479 ( .A(n2979), .B(n2980), .Z(n2978) );
  XOR U3480 ( .A(n2981), .B(n2982), .Z(n2977) );
  XNOR U3481 ( .A(key[1149]), .B(n2983), .Z(n2982) );
  XOR U3482 ( .A(n2984), .B(n2985), .Z(n2966) );
  XNOR U3483 ( .A(n2986), .B(n2987), .Z(n2985) );
  XOR U3484 ( .A(key[1151]), .B(n2988), .Z(n2984) );
  XOR U3485 ( .A(n2441), .B(n2545), .Z(n2902) );
  IV U3486 ( .A(n2936), .Z(n2545) );
  XNOR U3487 ( .A(n2965), .B(n2989), .Z(n2936) );
  XNOR U3488 ( .A(n2956), .B(n2975), .Z(n2989) );
  XOR U3489 ( .A(n2990), .B(n2991), .Z(n2975) );
  XNOR U3490 ( .A(n2992), .B(n2993), .Z(n2991) );
  XOR U3491 ( .A(n2994), .B(n2995), .Z(n2990) );
  XNOR U3492 ( .A(key[1146]), .B(n2996), .Z(n2995) );
  XOR U3493 ( .A(n2997), .B(n2998), .Z(n2956) );
  XOR U3494 ( .A(n2999), .B(n2441), .Z(n2998) );
  XOR U3495 ( .A(n3000), .B(n3001), .Z(n2997) );
  XOR U3496 ( .A(key[1150]), .B(n3002), .Z(n3001) );
  XOR U3497 ( .A(n3003), .B(n3004), .Z(n2965) );
  XOR U3498 ( .A(n2957), .B(n3005), .Z(n3004) );
  XOR U3499 ( .A(n3006), .B(n3007), .Z(n3005) );
  XNOR U3500 ( .A(n3008), .B(n3009), .Z(n2957) );
  XOR U3501 ( .A(n3010), .B(n3011), .Z(n3009) );
  XNOR U3502 ( .A(n3012), .B(n3013), .Z(n3008) );
  XOR U3503 ( .A(key[1145]), .B(n3014), .Z(n3013) );
  XNOR U3504 ( .A(n3015), .B(n3016), .Z(n3003) );
  XNOR U3505 ( .A(key[1147]), .B(n3017), .Z(n3016) );
  IV U3506 ( .A(n2941), .Z(n2441) );
  XOR U3507 ( .A(n3018), .B(n3019), .Z(n2941) );
  XNOR U3508 ( .A(n3020), .B(n3021), .Z(n3019) );
  XOR U3509 ( .A(n3022), .B(n3023), .Z(n3018) );
  XOR U3510 ( .A(key[1144]), .B(n3024), .Z(n3023) );
  IV U3511 ( .A(n2115), .Z(n2338) );
  XOR U3512 ( .A(n2851), .B(n2423), .Z(n2115) );
  XNOR U3513 ( .A(n2417), .B(n3025), .Z(n2423) );
  XNOR U3514 ( .A(n3026), .B(n2848), .Z(n3025) );
  XOR U3515 ( .A(n3028), .B(n2427), .Z(n2459) );
  ANDN U3516 ( .B(n3029), .A(n2462), .Z(n3026) );
  IV U3517 ( .A(n3028), .Z(n2462) );
  XNOR U3518 ( .A(n2846), .B(n3030), .Z(n2417) );
  XNOR U3519 ( .A(n3031), .B(n3032), .Z(n3030) );
  NANDN U3520 ( .A(n2844), .B(n3033), .Z(n3032) );
  IV U3521 ( .A(n2502), .Z(n2851) );
  XNOR U3522 ( .A(n2846), .B(n3034), .Z(n2502) );
  XOR U3523 ( .A(n3035), .B(n2419), .Z(n3034) );
  OR U3524 ( .A(n3036), .B(n2856), .Z(n2419) );
  XNOR U3525 ( .A(n2422), .B(n2855), .Z(n2856) );
  ANDN U3526 ( .B(n3037), .A(n3038), .Z(n3035) );
  XOR U3527 ( .A(n3039), .B(n3031), .Z(n2846) );
  OR U3528 ( .A(n2859), .B(n3040), .Z(n3031) );
  XNOR U3529 ( .A(n2862), .B(n2844), .Z(n2859) );
  XNOR U3530 ( .A(n2855), .B(n2427), .Z(n2844) );
  XOR U3531 ( .A(n3041), .B(n3042), .Z(n2427) );
  NANDN U3532 ( .A(n3043), .B(n3044), .Z(n3042) );
  IV U3533 ( .A(n3038), .Z(n2855) );
  XNOR U3534 ( .A(n3045), .B(n3046), .Z(n3038) );
  NANDN U3535 ( .A(n3043), .B(n3047), .Z(n3046) );
  NOR U3536 ( .A(n2862), .B(n3048), .Z(n3039) );
  XNOR U3537 ( .A(n3028), .B(n2422), .Z(n2862) );
  XNOR U3538 ( .A(n3049), .B(n3045), .Z(n2422) );
  NANDN U3539 ( .A(n3050), .B(n3051), .Z(n3045) );
  XOR U3540 ( .A(n3047), .B(n3052), .Z(n3051) );
  ANDN U3541 ( .B(n3052), .A(n3053), .Z(n3049) );
  XNOR U3542 ( .A(n3054), .B(n3041), .Z(n3028) );
  NANDN U3543 ( .A(n3050), .B(n3055), .Z(n3041) );
  XOR U3544 ( .A(n3056), .B(n3044), .Z(n3055) );
  XNOR U3545 ( .A(n3057), .B(n3058), .Z(n3043) );
  XOR U3546 ( .A(n3059), .B(n3060), .Z(n3058) );
  XNOR U3547 ( .A(n3061), .B(n3062), .Z(n3057) );
  XNOR U3548 ( .A(n3063), .B(n3064), .Z(n3062) );
  ANDN U3549 ( .B(n3056), .A(n3060), .Z(n3063) );
  ANDN U3550 ( .B(n3056), .A(n3053), .Z(n3054) );
  XNOR U3551 ( .A(n3059), .B(n3065), .Z(n3053) );
  XOR U3552 ( .A(n3066), .B(n3064), .Z(n3065) );
  NAND U3553 ( .A(n3067), .B(n3068), .Z(n3064) );
  XNOR U3554 ( .A(n3061), .B(n3044), .Z(n3068) );
  IV U3555 ( .A(n3056), .Z(n3061) );
  XNOR U3556 ( .A(n3047), .B(n3060), .Z(n3067) );
  IV U3557 ( .A(n3052), .Z(n3060) );
  XOR U3558 ( .A(n3069), .B(n3070), .Z(n3052) );
  XNOR U3559 ( .A(n3071), .B(n3072), .Z(n3070) );
  XNOR U3560 ( .A(n3073), .B(n3074), .Z(n3069) );
  ANDN U3561 ( .B(n3029), .A(n3075), .Z(n3073) );
  AND U3562 ( .A(n3044), .B(n3047), .Z(n3066) );
  XNOR U3563 ( .A(n3044), .B(n3047), .Z(n3059) );
  XNOR U3564 ( .A(n3076), .B(n3077), .Z(n3047) );
  XNOR U3565 ( .A(n3078), .B(n3072), .Z(n3077) );
  XOR U3566 ( .A(n3079), .B(n3080), .Z(n3076) );
  XNOR U3567 ( .A(n3081), .B(n3074), .Z(n3080) );
  OR U3568 ( .A(n2460), .B(n3027), .Z(n3074) );
  XNOR U3569 ( .A(n3029), .B(n3082), .Z(n3027) );
  XNOR U3570 ( .A(n3075), .B(n2428), .Z(n2460) );
  ANDN U3571 ( .B(n3083), .A(n2850), .Z(n3081) );
  XNOR U3572 ( .A(n3084), .B(n3085), .Z(n3044) );
  XNOR U3573 ( .A(n3072), .B(n3086), .Z(n3085) );
  XOR U3574 ( .A(n2840), .B(n3079), .Z(n3086) );
  XNOR U3575 ( .A(n3029), .B(n3075), .Z(n3072) );
  XNOR U3576 ( .A(n3087), .B(n3088), .Z(n3084) );
  XNOR U3577 ( .A(n3089), .B(n3090), .Z(n3088) );
  ANDN U3578 ( .B(n3037), .A(n2854), .Z(n3089) );
  XNOR U3579 ( .A(n3091), .B(n3092), .Z(n3056) );
  XNOR U3580 ( .A(n3078), .B(n3093), .Z(n3092) );
  XNOR U3581 ( .A(n2854), .B(n3071), .Z(n3093) );
  XOR U3582 ( .A(n3079), .B(n3094), .Z(n3071) );
  XNOR U3583 ( .A(n3095), .B(n3096), .Z(n3094) );
  NAND U3584 ( .A(n3033), .B(n2845), .Z(n3096) );
  XNOR U3585 ( .A(n3097), .B(n3095), .Z(n3079) );
  NANDN U3586 ( .A(n3040), .B(n2860), .Z(n3095) );
  XOR U3587 ( .A(n2861), .B(n2845), .Z(n2860) );
  XNOR U3588 ( .A(n3098), .B(n2428), .Z(n2845) );
  XOR U3589 ( .A(n3048), .B(n3033), .Z(n3040) );
  XOR U3590 ( .A(n3037), .B(n3082), .Z(n3033) );
  ANDN U3591 ( .B(n2861), .A(n3048), .Z(n3097) );
  XNOR U3592 ( .A(n3087), .B(n3029), .Z(n3048) );
  XNOR U3593 ( .A(n3099), .B(n3100), .Z(n3029) );
  XNOR U3594 ( .A(n3101), .B(n3102), .Z(n3100) );
  XOR U3595 ( .A(n3103), .B(n2461), .Z(n2861) );
  XOR U3596 ( .A(n3082), .B(n3083), .Z(n3078) );
  IV U3597 ( .A(n2428), .Z(n3083) );
  XOR U3598 ( .A(n3104), .B(n3105), .Z(n2428) );
  XNOR U3599 ( .A(n3106), .B(n3102), .Z(n3105) );
  IV U3600 ( .A(n2850), .Z(n3082) );
  XOR U3601 ( .A(n3102), .B(n3107), .Z(n2850) );
  XNOR U3602 ( .A(n3037), .B(n3108), .Z(n3091) );
  XNOR U3603 ( .A(n3109), .B(n3090), .Z(n3108) );
  OR U3604 ( .A(n2857), .B(n3036), .Z(n3090) );
  XNOR U3605 ( .A(n3087), .B(n3037), .Z(n3036) );
  XOR U3606 ( .A(n2840), .B(n3098), .Z(n2857) );
  IV U3607 ( .A(n2854), .Z(n3098) );
  XOR U3608 ( .A(n2461), .B(n3110), .Z(n2854) );
  XNOR U3609 ( .A(n3106), .B(n3099), .Z(n3110) );
  XOR U3610 ( .A(n3111), .B(n3112), .Z(n3099) );
  XNOR U3611 ( .A(n3113), .B(n3114), .Z(n3112) );
  XOR U3612 ( .A(key[1106]), .B(n3115), .Z(n3111) );
  IV U3613 ( .A(n3075), .Z(n2461) );
  XOR U3614 ( .A(n3104), .B(n3116), .Z(n3075) );
  XOR U3615 ( .A(n3102), .B(n3117), .Z(n3116) );
  ANDN U3616 ( .B(n3103), .A(n2421), .Z(n3109) );
  IV U3617 ( .A(n2840), .Z(n3103) );
  XOR U3618 ( .A(n3104), .B(n3118), .Z(n2840) );
  XOR U3619 ( .A(n3102), .B(n3119), .Z(n3118) );
  XOR U3620 ( .A(n3120), .B(n3121), .Z(n3102) );
  XOR U3621 ( .A(n3122), .B(n2421), .Z(n3121) );
  IV U3622 ( .A(n3087), .Z(n2421) );
  XNOR U3623 ( .A(n3123), .B(n3124), .Z(n3120) );
  XNOR U3624 ( .A(key[1110]), .B(n3125), .Z(n3124) );
  IV U3625 ( .A(n3107), .Z(n3104) );
  XOR U3626 ( .A(n3126), .B(n3127), .Z(n3107) );
  XNOR U3627 ( .A(n3128), .B(n3129), .Z(n3127) );
  XNOR U3628 ( .A(key[1109]), .B(n3130), .Z(n3126) );
  XOR U3629 ( .A(n3131), .B(n3132), .Z(n3037) );
  XNOR U3630 ( .A(n3119), .B(n3117), .Z(n3132) );
  XNOR U3631 ( .A(n3133), .B(n3134), .Z(n3117) );
  XOR U3632 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U3633 ( .A(key[1111]), .B(n3137), .Z(n3133) );
  XNOR U3634 ( .A(n3138), .B(n3139), .Z(n3119) );
  XOR U3635 ( .A(n3140), .B(n3141), .Z(n3138) );
  XNOR U3636 ( .A(key[1108]), .B(n3142), .Z(n3141) );
  XOR U3637 ( .A(n3087), .B(n3101), .Z(n3131) );
  XOR U3638 ( .A(n3143), .B(n3144), .Z(n3101) );
  XNOR U3639 ( .A(n3106), .B(n3145), .Z(n3144) );
  XNOR U3640 ( .A(n3146), .B(n3147), .Z(n3145) );
  XOR U3641 ( .A(n3148), .B(n3149), .Z(n3106) );
  XNOR U3642 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U3643 ( .A(key[1105]), .B(n3152), .Z(n3148) );
  XNOR U3644 ( .A(n3153), .B(n3154), .Z(n3143) );
  XNOR U3645 ( .A(key[1107]), .B(n3155), .Z(n3154) );
  XOR U3646 ( .A(n3156), .B(n3157), .Z(n3087) );
  XNOR U3647 ( .A(n3158), .B(n3159), .Z(n3157) );
  XNOR U3648 ( .A(key[1104]), .B(n3160), .Z(n3156) );
  XOR U3649 ( .A(n3161), .B(n3162), .Z(out[11]) );
  XNOR U3650 ( .A(n4), .B(n2137), .Z(n3162) );
  XNOR U3651 ( .A(n3163), .B(n3164), .Z(n2137) );
  XNOR U3652 ( .A(n3165), .B(n2153), .Z(n3164) );
  ANDN U3653 ( .B(n3166), .A(n3167), .Z(n2153) );
  NOR U3654 ( .A(n2162), .B(n3168), .Z(n3165) );
  XNOR U3655 ( .A(n2139), .B(n3169), .Z(n3161) );
  XOR U3656 ( .A(key[1163]), .B(n5), .Z(n3169) );
  XOR U3657 ( .A(n3163), .B(n3170), .Z(n5) );
  XNOR U3658 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3659 ( .A(n2149), .B(n3173), .Z(n3172) );
  XNOR U3660 ( .A(n2144), .B(n3174), .Z(n3163) );
  XNOR U3661 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3662 ( .A(n3177), .B(n2167), .Z(n3176) );
  XNOR U3663 ( .A(n2144), .B(n3178), .Z(n2139) );
  XNOR U3664 ( .A(n3171), .B(n3179), .Z(n3178) );
  NANDN U3665 ( .A(n3180), .B(n3181), .Z(n3179) );
  OR U3666 ( .A(n3182), .B(n3183), .Z(n3171) );
  XOR U3667 ( .A(n3184), .B(n3175), .Z(n2144) );
  OR U3668 ( .A(n3185), .B(n3186), .Z(n3175) );
  ANDN U3669 ( .B(n3187), .A(n3188), .Z(n3184) );
  XOR U3670 ( .A(n3189), .B(n3190), .Z(out[119]) );
  XOR U3671 ( .A(n3191), .B(n3192), .Z(n3189) );
  XNOR U3672 ( .A(key[1271]), .B(n3193), .Z(n3192) );
  XNOR U3673 ( .A(n3194), .B(n3195), .Z(out[118]) );
  XNOR U3674 ( .A(key[1270]), .B(n3196), .Z(n3195) );
  XOR U3675 ( .A(n3197), .B(n3198), .Z(out[117]) );
  XNOR U3676 ( .A(n3199), .B(n3200), .Z(n3198) );
  XOR U3677 ( .A(n3191), .B(n3201), .Z(n3200) );
  XNOR U3678 ( .A(n3203), .B(n3204), .Z(n3202) );
  NANDN U3679 ( .A(n3205), .B(n3206), .Z(n3204) );
  XOR U3680 ( .A(n3208), .B(n3209), .Z(n3197) );
  XOR U3681 ( .A(key[1269]), .B(n3210), .Z(n3209) );
  ANDN U3682 ( .B(n3211), .A(n3212), .Z(n3208) );
  XNOR U3683 ( .A(n3213), .B(n3214), .Z(out[116]) );
  XNOR U3684 ( .A(key[1268]), .B(n3215), .Z(n3214) );
  XOR U3685 ( .A(n3216), .B(n3217), .Z(out[115]) );
  XNOR U3686 ( .A(n3218), .B(n3194), .Z(n3217) );
  XNOR U3687 ( .A(n3219), .B(n3220), .Z(n3194) );
  XNOR U3688 ( .A(n3221), .B(n3210), .Z(n3220) );
  ANDN U3689 ( .B(n3222), .A(n3223), .Z(n3210) );
  NOR U3690 ( .A(n3224), .B(n3225), .Z(n3221) );
  XNOR U3691 ( .A(n3226), .B(n3227), .Z(n3216) );
  XOR U3692 ( .A(key[1267]), .B(n3228), .Z(n3227) );
  XOR U3693 ( .A(key[1266]), .B(n3213), .Z(out[114]) );
  XNOR U3694 ( .A(n3193), .B(n3229), .Z(n3213) );
  IV U3695 ( .A(n3228), .Z(n3193) );
  XOR U3696 ( .A(n3230), .B(n3190), .Z(out[113]) );
  XNOR U3697 ( .A(n3219), .B(n3231), .Z(n3218) );
  XNOR U3698 ( .A(n3232), .B(n3233), .Z(n3231) );
  NANDN U3699 ( .A(n3234), .B(n3206), .Z(n3233) );
  XNOR U3700 ( .A(n3201), .B(n3235), .Z(n3219) );
  XNOR U3701 ( .A(n3236), .B(n3237), .Z(n3235) );
  NANDN U3702 ( .A(n3238), .B(n3239), .Z(n3237) );
  XOR U3703 ( .A(n3229), .B(n3226), .Z(n3196) );
  XNOR U3704 ( .A(n3201), .B(n3240), .Z(n3226) );
  XNOR U3705 ( .A(n3232), .B(n3241), .Z(n3240) );
  NANDN U3706 ( .A(n3242), .B(n3243), .Z(n3241) );
  OR U3707 ( .A(n3244), .B(n3245), .Z(n3232) );
  XOR U3708 ( .A(n3246), .B(n3236), .Z(n3201) );
  NANDN U3709 ( .A(n3247), .B(n3248), .Z(n3236) );
  ANDN U3710 ( .B(n3249), .A(n3250), .Z(n3246) );
  XOR U3711 ( .A(key[1265]), .B(n3228), .Z(n3230) );
  XOR U3712 ( .A(n3251), .B(n3252), .Z(n3228) );
  XNOR U3713 ( .A(n3253), .B(n3254), .Z(n3252) );
  NANDN U3714 ( .A(n3255), .B(n3211), .Z(n3254) );
  XNOR U3715 ( .A(n3199), .B(n3256), .Z(out[112]) );
  XOR U3716 ( .A(key[1264]), .B(n3229), .Z(n3256) );
  XNOR U3717 ( .A(n3251), .B(n3257), .Z(n3229) );
  XOR U3718 ( .A(n3258), .B(n3203), .Z(n3257) );
  OR U3719 ( .A(n3259), .B(n3244), .Z(n3203) );
  XNOR U3720 ( .A(n3206), .B(n3243), .Z(n3244) );
  ANDN U3721 ( .B(n3260), .A(n3261), .Z(n3258) );
  IV U3722 ( .A(n3215), .Z(n3199) );
  XOR U3723 ( .A(n3207), .B(n3262), .Z(n3215) );
  XOR U3724 ( .A(n3263), .B(n3253), .Z(n3262) );
  XNOR U3725 ( .A(n3225), .B(n3211), .Z(n3222) );
  NOR U3726 ( .A(n3265), .B(n3225), .Z(n3263) );
  XNOR U3727 ( .A(n3251), .B(n3266), .Z(n3207) );
  XNOR U3728 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3729 ( .A(n3238), .B(n3269), .Z(n3268) );
  XOR U3730 ( .A(n3270), .B(n3267), .Z(n3251) );
  OR U3731 ( .A(n3247), .B(n3271), .Z(n3267) );
  XOR U3732 ( .A(n3272), .B(n3238), .Z(n3247) );
  XNOR U3733 ( .A(n3243), .B(n3211), .Z(n3238) );
  XOR U3734 ( .A(n3273), .B(n3274), .Z(n3211) );
  NANDN U3735 ( .A(n3275), .B(n3276), .Z(n3274) );
  IV U3736 ( .A(n3261), .Z(n3243) );
  XNOR U3737 ( .A(n3277), .B(n3278), .Z(n3261) );
  NANDN U3738 ( .A(n3275), .B(n3279), .Z(n3278) );
  ANDN U3739 ( .B(n3272), .A(n3280), .Z(n3270) );
  IV U3740 ( .A(n3250), .Z(n3272) );
  XOR U3741 ( .A(n3225), .B(n3206), .Z(n3250) );
  XNOR U3742 ( .A(n3281), .B(n3277), .Z(n3206) );
  NANDN U3743 ( .A(n3282), .B(n3283), .Z(n3277) );
  XOR U3744 ( .A(n3279), .B(n3284), .Z(n3283) );
  ANDN U3745 ( .B(n3284), .A(n3285), .Z(n3281) );
  XOR U3746 ( .A(n3286), .B(n3273), .Z(n3225) );
  NANDN U3747 ( .A(n3282), .B(n3287), .Z(n3273) );
  XOR U3748 ( .A(n3288), .B(n3276), .Z(n3287) );
  XNOR U3749 ( .A(n3289), .B(n3290), .Z(n3275) );
  XOR U3750 ( .A(n3291), .B(n3292), .Z(n3290) );
  XNOR U3751 ( .A(n3293), .B(n3294), .Z(n3289) );
  XNOR U3752 ( .A(n3295), .B(n3296), .Z(n3294) );
  ANDN U3753 ( .B(n3288), .A(n3292), .Z(n3295) );
  ANDN U3754 ( .B(n3288), .A(n3285), .Z(n3286) );
  XNOR U3755 ( .A(n3291), .B(n3297), .Z(n3285) );
  XOR U3756 ( .A(n3298), .B(n3296), .Z(n3297) );
  NAND U3757 ( .A(n3299), .B(n3300), .Z(n3296) );
  XNOR U3758 ( .A(n3293), .B(n3276), .Z(n3300) );
  IV U3759 ( .A(n3288), .Z(n3293) );
  XNOR U3760 ( .A(n3279), .B(n3292), .Z(n3299) );
  IV U3761 ( .A(n3284), .Z(n3292) );
  XOR U3762 ( .A(n3301), .B(n3302), .Z(n3284) );
  XNOR U3763 ( .A(n3303), .B(n3304), .Z(n3302) );
  XNOR U3764 ( .A(n3305), .B(n3306), .Z(n3301) );
  NOR U3765 ( .A(n3224), .B(n3265), .Z(n3305) );
  AND U3766 ( .A(n3276), .B(n3279), .Z(n3298) );
  XNOR U3767 ( .A(n3276), .B(n3279), .Z(n3291) );
  XNOR U3768 ( .A(n3307), .B(n3308), .Z(n3279) );
  XNOR U3769 ( .A(n3309), .B(n3304), .Z(n3308) );
  XOR U3770 ( .A(n3310), .B(n3311), .Z(n3307) );
  XNOR U3771 ( .A(n3312), .B(n3306), .Z(n3311) );
  OR U3772 ( .A(n3223), .B(n3264), .Z(n3306) );
  XNOR U3773 ( .A(n3265), .B(n3255), .Z(n3264) );
  XNOR U3774 ( .A(n3224), .B(n3212), .Z(n3223) );
  ANDN U3775 ( .B(n3313), .A(n3255), .Z(n3312) );
  XNOR U3776 ( .A(n3314), .B(n3315), .Z(n3276) );
  XNOR U3777 ( .A(n3304), .B(n3316), .Z(n3315) );
  XOR U3778 ( .A(n3234), .B(n3310), .Z(n3316) );
  XNOR U3779 ( .A(n3265), .B(n3317), .Z(n3304) );
  XNOR U3780 ( .A(n3318), .B(n3319), .Z(n3314) );
  XNOR U3781 ( .A(n3320), .B(n3321), .Z(n3319) );
  ANDN U3782 ( .B(n3260), .A(n3242), .Z(n3320) );
  XNOR U3783 ( .A(n3322), .B(n3323), .Z(n3288) );
  XNOR U3784 ( .A(n3309), .B(n3324), .Z(n3323) );
  XNOR U3785 ( .A(n3242), .B(n3303), .Z(n3324) );
  XOR U3786 ( .A(n3310), .B(n3325), .Z(n3303) );
  XNOR U3787 ( .A(n3326), .B(n3327), .Z(n3325) );
  NAND U3788 ( .A(n3269), .B(n3239), .Z(n3327) );
  XNOR U3789 ( .A(n3328), .B(n3326), .Z(n3310) );
  NANDN U3790 ( .A(n3271), .B(n3248), .Z(n3326) );
  XOR U3791 ( .A(n3249), .B(n3239), .Z(n3248) );
  XNOR U3792 ( .A(n3329), .B(n3212), .Z(n3239) );
  XOR U3793 ( .A(n3280), .B(n3269), .Z(n3271) );
  XOR U3794 ( .A(n3260), .B(n3330), .Z(n3269) );
  ANDN U3795 ( .B(n3249), .A(n3280), .Z(n3328) );
  XOR U3796 ( .A(n3318), .B(n3265), .Z(n3280) );
  XOR U3797 ( .A(n3331), .B(n3332), .Z(n3265) );
  XNOR U3798 ( .A(n3333), .B(n3334), .Z(n3332) );
  XOR U3799 ( .A(n3335), .B(n3317), .Z(n3249) );
  XOR U3800 ( .A(n3330), .B(n3313), .Z(n3309) );
  IV U3801 ( .A(n3212), .Z(n3313) );
  XOR U3802 ( .A(n3336), .B(n3337), .Z(n3212) );
  XNOR U3803 ( .A(n3338), .B(n3334), .Z(n3337) );
  IV U3804 ( .A(n3255), .Z(n3330) );
  XOR U3805 ( .A(n3334), .B(n3339), .Z(n3255) );
  XNOR U3806 ( .A(n3260), .B(n3340), .Z(n3322) );
  XNOR U3807 ( .A(n3341), .B(n3321), .Z(n3340) );
  OR U3808 ( .A(n3245), .B(n3259), .Z(n3321) );
  XNOR U3809 ( .A(n3318), .B(n3260), .Z(n3259) );
  XOR U3810 ( .A(n3234), .B(n3329), .Z(n3245) );
  IV U3811 ( .A(n3242), .Z(n3329) );
  XOR U3812 ( .A(n3317), .B(n3342), .Z(n3242) );
  XNOR U3813 ( .A(n3338), .B(n3331), .Z(n3342) );
  XOR U3814 ( .A(n3343), .B(n3344), .Z(n3331) );
  XOR U3815 ( .A(n1705), .B(n215), .Z(n3344) );
  XOR U3816 ( .A(n3345), .B(n177), .Z(n215) );
  XOR U3817 ( .A(key[1234]), .B(n3346), .Z(n3343) );
  IV U3818 ( .A(n3224), .Z(n3317) );
  XOR U3819 ( .A(n3336), .B(n3347), .Z(n3224) );
  XOR U3820 ( .A(n3334), .B(n3348), .Z(n3347) );
  ANDN U3821 ( .B(n3335), .A(n3205), .Z(n3341) );
  IV U3822 ( .A(n3234), .Z(n3335) );
  XOR U3823 ( .A(n3336), .B(n3349), .Z(n3234) );
  XOR U3824 ( .A(n3334), .B(n3350), .Z(n3349) );
  XOR U3825 ( .A(n3351), .B(n3352), .Z(n3334) );
  XOR U3826 ( .A(n188), .B(n3205), .Z(n3352) );
  IV U3827 ( .A(n3318), .Z(n3205) );
  XNOR U3828 ( .A(n3353), .B(n1689), .Z(n188) );
  XNOR U3829 ( .A(n3354), .B(n3355), .Z(n3351) );
  XOR U3830 ( .A(key[1238]), .B(n3356), .Z(n3355) );
  IV U3831 ( .A(n3339), .Z(n3336) );
  XOR U3832 ( .A(n3357), .B(n3358), .Z(n3339) );
  XOR U3833 ( .A(n1682), .B(n1674), .Z(n3358) );
  XNOR U3834 ( .A(n3356), .B(n3359), .Z(n1674) );
  XNOR U3835 ( .A(key[1237]), .B(n3360), .Z(n3357) );
  XOR U3836 ( .A(n3361), .B(n3362), .Z(n3260) );
  XNOR U3837 ( .A(n3350), .B(n3348), .Z(n3362) );
  XNOR U3838 ( .A(n3363), .B(n3364), .Z(n3348) );
  XNOR U3839 ( .A(n3365), .B(n3366), .Z(n3364) );
  XNOR U3840 ( .A(key[1239]), .B(n234), .Z(n3363) );
  XNOR U3841 ( .A(n3367), .B(n3368), .Z(n3350) );
  XOR U3842 ( .A(n1696), .B(n208), .Z(n3368) );
  XNOR U3843 ( .A(n3369), .B(n234), .Z(n208) );
  XOR U3844 ( .A(n3370), .B(n3371), .Z(n3367) );
  XNOR U3845 ( .A(key[1236]), .B(n3372), .Z(n3371) );
  XOR U3846 ( .A(n3318), .B(n3333), .Z(n3361) );
  XOR U3847 ( .A(n3373), .B(n3374), .Z(n3333) );
  XNOR U3848 ( .A(n3338), .B(n3375), .Z(n3374) );
  XNOR U3849 ( .A(n3376), .B(n217), .Z(n3375) );
  XOR U3850 ( .A(n3353), .B(n1695), .Z(n217) );
  XOR U3851 ( .A(n3377), .B(n3378), .Z(n3338) );
  XNOR U3852 ( .A(n1712), .B(n178), .Z(n3378) );
  XNOR U3853 ( .A(n222), .B(n3346), .Z(n178) );
  XOR U3854 ( .A(key[1233]), .B(n3379), .Z(n3377) );
  XNOR U3855 ( .A(n3380), .B(n3381), .Z(n3373) );
  XOR U3856 ( .A(key[1235]), .B(n3382), .Z(n3381) );
  XOR U3857 ( .A(n3383), .B(n3384), .Z(n3318) );
  XNOR U3858 ( .A(n232), .B(n221), .Z(n3384) );
  XOR U3859 ( .A(n3379), .B(n231), .Z(n221) );
  XOR U3860 ( .A(key[1232]), .B(n1690), .Z(n3383) );
  XOR U3861 ( .A(n3385), .B(n3386), .Z(out[111]) );
  XOR U3862 ( .A(n3387), .B(n3388), .Z(n3385) );
  XNOR U3863 ( .A(key[1263]), .B(n3389), .Z(n3388) );
  XNOR U3864 ( .A(n3390), .B(n3391), .Z(out[110]) );
  XNOR U3865 ( .A(key[1262]), .B(n3392), .Z(n3391) );
  XOR U3866 ( .A(key[1162]), .B(n2156), .Z(out[10]) );
  XNOR U3867 ( .A(n2140), .B(n4), .Z(n2156) );
  XNOR U3868 ( .A(n2163), .B(n3393), .Z(n4) );
  XNOR U3869 ( .A(n2160), .B(n3394), .Z(n3393) );
  NANDN U3870 ( .A(n3395), .B(n2154), .Z(n3394) );
  XNOR U3871 ( .A(n2162), .B(n2154), .Z(n3166) );
  XNOR U3872 ( .A(n2163), .B(n3397), .Z(n2140) );
  XOR U3873 ( .A(n3398), .B(n2147), .Z(n3397) );
  OR U3874 ( .A(n3182), .B(n3399), .Z(n2147) );
  XNOR U3875 ( .A(n2149), .B(n3180), .Z(n3182) );
  NOR U3876 ( .A(n3400), .B(n3180), .Z(n3398) );
  XOR U3877 ( .A(n3401), .B(n2165), .Z(n2163) );
  NANDN U3878 ( .A(n3186), .B(n3402), .Z(n2165) );
  XNOR U3879 ( .A(n3187), .B(n2167), .Z(n3186) );
  XNOR U3880 ( .A(n3180), .B(n2154), .Z(n2167) );
  XOR U3881 ( .A(n3403), .B(n3404), .Z(n2154) );
  NANDN U3882 ( .A(n3405), .B(n3406), .Z(n3404) );
  XNOR U3883 ( .A(n3407), .B(n3408), .Z(n3180) );
  OR U3884 ( .A(n3405), .B(n3409), .Z(n3408) );
  AND U3885 ( .A(n3187), .B(n3410), .Z(n3401) );
  XOR U3886 ( .A(n2149), .B(n2162), .Z(n3187) );
  XOR U3887 ( .A(n3411), .B(n3403), .Z(n2162) );
  NANDN U3888 ( .A(n3412), .B(n3413), .Z(n3403) );
  ANDN U3889 ( .B(n3414), .A(n3415), .Z(n3411) );
  NANDN U3890 ( .A(n3412), .B(n3417), .Z(n3407) );
  XOR U3891 ( .A(n3418), .B(n3405), .Z(n3412) );
  XNOR U3892 ( .A(n3419), .B(n3420), .Z(n3405) );
  XOR U3893 ( .A(n3421), .B(n3414), .Z(n3420) );
  XNOR U3894 ( .A(n3422), .B(n3423), .Z(n3419) );
  XNOR U3895 ( .A(n3424), .B(n3425), .Z(n3423) );
  ANDN U3896 ( .B(n3414), .A(n3426), .Z(n3424) );
  IV U3897 ( .A(n3427), .Z(n3414) );
  ANDN U3898 ( .B(n3418), .A(n3426), .Z(n3416) );
  IV U3899 ( .A(n3422), .Z(n3426) );
  IV U3900 ( .A(n3415), .Z(n3418) );
  XNOR U3901 ( .A(n3421), .B(n3428), .Z(n3415) );
  XOR U3902 ( .A(n3429), .B(n3425), .Z(n3428) );
  NAND U3903 ( .A(n3417), .B(n3413), .Z(n3425) );
  XNOR U3904 ( .A(n3406), .B(n3427), .Z(n3413) );
  XOR U3905 ( .A(n3430), .B(n3431), .Z(n3427) );
  XOR U3906 ( .A(n3432), .B(n3433), .Z(n3431) );
  XOR U3907 ( .A(n3434), .B(n3435), .Z(n3433) );
  XOR U3908 ( .A(n3181), .B(n3436), .Z(n3430) );
  XNOR U3909 ( .A(n3437), .B(n3438), .Z(n3436) );
  AND U3910 ( .A(n3173), .B(n2150), .Z(n3437) );
  XNOR U3911 ( .A(n3422), .B(n3409), .Z(n3417) );
  XOR U3912 ( .A(n3439), .B(n3440), .Z(n3422) );
  XNOR U3913 ( .A(n3441), .B(n3435), .Z(n3440) );
  XOR U3914 ( .A(n3442), .B(n3443), .Z(n3435) );
  XNOR U3915 ( .A(n3444), .B(n3445), .Z(n3443) );
  NAND U3916 ( .A(n2168), .B(n3177), .Z(n3445) );
  XNOR U3917 ( .A(n3446), .B(n3447), .Z(n3439) );
  ANDN U3918 ( .B(n2161), .A(n3168), .Z(n3446) );
  ANDN U3919 ( .B(n3406), .A(n3409), .Z(n3429) );
  XOR U3920 ( .A(n3409), .B(n3406), .Z(n3421) );
  XNOR U3921 ( .A(n3448), .B(n3449), .Z(n3406) );
  XNOR U3922 ( .A(n3442), .B(n3450), .Z(n3449) );
  XNOR U3923 ( .A(n3173), .B(n3441), .Z(n3450) );
  XNOR U3924 ( .A(n2150), .B(n3451), .Z(n3448) );
  XNOR U3925 ( .A(n3452), .B(n3438), .Z(n3451) );
  OR U3926 ( .A(n3183), .B(n3399), .Z(n3438) );
  XNOR U3927 ( .A(n2150), .B(n3434), .Z(n3399) );
  XNOR U3928 ( .A(n3173), .B(n3181), .Z(n3183) );
  ANDN U3929 ( .B(n3181), .A(n3400), .Z(n3452) );
  IV U3930 ( .A(n3434), .Z(n3400) );
  XOR U3931 ( .A(n3453), .B(n3454), .Z(n3409) );
  XOR U3932 ( .A(n3442), .B(n3432), .Z(n3454) );
  XOR U3933 ( .A(n3455), .B(n3395), .Z(n3432) );
  XOR U3934 ( .A(n3456), .B(n3444), .Z(n3442) );
  NANDN U3935 ( .A(n3185), .B(n3402), .Z(n3444) );
  XOR U3936 ( .A(n3410), .B(n2168), .Z(n3402) );
  XNOR U3937 ( .A(n3395), .B(n3434), .Z(n2168) );
  XOR U3938 ( .A(n3457), .B(n3458), .Z(n3434) );
  XNOR U3939 ( .A(n3459), .B(n3460), .Z(n3458) );
  XOR U3940 ( .A(n2150), .B(n3461), .Z(n3457) );
  XOR U3941 ( .A(n3188), .B(n3177), .Z(n3185) );
  XOR U3942 ( .A(n3455), .B(n3181), .Z(n3177) );
  XOR U3943 ( .A(n3462), .B(n3463), .Z(n3181) );
  XNOR U3944 ( .A(n3168), .B(n3464), .Z(n3463) );
  ANDN U3945 ( .B(n3410), .A(n3188), .Z(n3456) );
  XOR U3946 ( .A(n3168), .B(n3173), .Z(n3188) );
  XOR U3947 ( .A(n3459), .B(n3465), .Z(n3173) );
  XOR U3948 ( .A(n3466), .B(n3467), .Z(n3465) );
  XOR U3949 ( .A(n3468), .B(n3469), .Z(n3459) );
  XNOR U3950 ( .A(n1695), .B(n3370), .Z(n3469) );
  XOR U3951 ( .A(n212), .B(n1697), .Z(n3370) );
  XOR U3952 ( .A(n3470), .B(n220), .Z(n1697) );
  XNOR U3953 ( .A(n3471), .B(n222), .Z(n1695) );
  XNOR U3954 ( .A(n1699), .B(n3472), .Z(n3468) );
  XNOR U3955 ( .A(key[1228]), .B(n3372), .Z(n3472) );
  XNOR U3956 ( .A(n1711), .B(n1682), .Z(n3372) );
  XNOR U3957 ( .A(n3473), .B(n3474), .Z(n1682) );
  XNOR U3958 ( .A(n3475), .B(n3476), .Z(n3474) );
  XNOR U3959 ( .A(n3477), .B(n3478), .Z(n3473) );
  XOR U3960 ( .A(n3479), .B(n3480), .Z(n3478) );
  ANDN U3961 ( .B(n3481), .A(n3482), .Z(n3480) );
  XOR U3962 ( .A(n198), .B(n3483), .Z(n1699) );
  XOR U3963 ( .A(n2150), .B(n2161), .Z(n3410) );
  XOR U3964 ( .A(n3441), .B(n3484), .Z(n3453) );
  XNOR U3965 ( .A(n3485), .B(n3447), .Z(n3484) );
  OR U3966 ( .A(n3396), .B(n3167), .Z(n3447) );
  XOR U3967 ( .A(n3168), .B(n3455), .Z(n3167) );
  XNOR U3968 ( .A(n2161), .B(n3487), .Z(n3396) );
  ANDN U3969 ( .B(n3455), .A(n3395), .Z(n3485) );
  XOR U3970 ( .A(n3486), .B(n3467), .Z(n3395) );
  IV U3971 ( .A(n2155), .Z(n3455) );
  XNOR U3972 ( .A(n3464), .B(n3487), .Z(n2155) );
  XOR U3973 ( .A(n3168), .B(n2161), .Z(n3441) );
  XNOR U3974 ( .A(n3460), .B(n3488), .Z(n2161) );
  XNOR U3975 ( .A(n3467), .B(n3462), .Z(n3488) );
  XOR U3976 ( .A(n3489), .B(n3490), .Z(n3462) );
  XNOR U3977 ( .A(n227), .B(n3345), .Z(n3490) );
  IV U3978 ( .A(n3382), .Z(n3345) );
  XNOR U3979 ( .A(n3491), .B(n3492), .Z(n3382) );
  XOR U3980 ( .A(n3493), .B(n3494), .Z(n3492) );
  XNOR U3981 ( .A(n3495), .B(n3496), .Z(n3491) );
  XOR U3982 ( .A(key[1226]), .B(n222), .Z(n3497) );
  XOR U3983 ( .A(n3498), .B(n3499), .Z(n222) );
  XOR U3984 ( .A(n3500), .B(n220), .Z(n1705) );
  XOR U3985 ( .A(n3501), .B(n3502), .Z(n220) );
  XOR U3986 ( .A(n3503), .B(n3504), .Z(n3460) );
  XOR U3987 ( .A(n177), .B(n3505), .Z(n3504) );
  XNOR U3988 ( .A(n1708), .B(n1667), .Z(n3505) );
  IV U3989 ( .A(n3376), .Z(n1667) );
  XOR U3990 ( .A(n227), .B(n179), .Z(n3376) );
  XOR U3991 ( .A(n3506), .B(n3507), .Z(n179) );
  XOR U3992 ( .A(n3508), .B(n3509), .Z(n3506) );
  XOR U3993 ( .A(n3510), .B(n3511), .Z(n227) );
  XNOR U3994 ( .A(n3512), .B(n3513), .Z(n3510) );
  XOR U3995 ( .A(n3483), .B(n212), .Z(n1708) );
  XNOR U3996 ( .A(n3514), .B(n181), .Z(n212) );
  XNOR U3997 ( .A(n3515), .B(n3516), .Z(n177) );
  XOR U3998 ( .A(n3517), .B(n3518), .Z(n3515) );
  XNOR U3999 ( .A(n3380), .B(n3519), .Z(n3503) );
  XNOR U4000 ( .A(key[1227]), .B(n3464), .Z(n3519) );
  XOR U4001 ( .A(n3520), .B(n3521), .Z(n3464) );
  XOR U4002 ( .A(n1712), .B(n231), .Z(n3521) );
  XOR U4003 ( .A(n3522), .B(n3523), .Z(n231) );
  XOR U4004 ( .A(n224), .B(n1706), .Z(n1712) );
  IV U4005 ( .A(n230), .Z(n1706) );
  XNOR U4006 ( .A(n3525), .B(n3526), .Z(n230) );
  XOR U4007 ( .A(n3346), .B(n3528), .Z(n3520) );
  XNOR U4008 ( .A(key[1225]), .B(n181), .Z(n3528) );
  IV U4009 ( .A(n3500), .Z(n181) );
  XNOR U4010 ( .A(n3529), .B(n3530), .Z(n3500) );
  XNOR U4011 ( .A(n1711), .B(n1696), .Z(n3380) );
  XNOR U4012 ( .A(n3475), .B(n3346), .Z(n1696) );
  XOR U4013 ( .A(n3531), .B(n3532), .Z(n3346) );
  XNOR U4014 ( .A(n3461), .B(n3487), .Z(n3168) );
  XNOR U4015 ( .A(n3486), .B(n3467), .Z(n3487) );
  XOR U4016 ( .A(n3533), .B(n3534), .Z(n3467) );
  XNOR U4017 ( .A(n196), .B(n3354), .Z(n3534) );
  XNOR U4018 ( .A(n1680), .B(n3365), .Z(n3354) );
  XOR U4019 ( .A(n1711), .B(n1688), .Z(n3365) );
  XOR U4020 ( .A(n3535), .B(n3536), .Z(n1688) );
  XNOR U4021 ( .A(n3537), .B(n3476), .Z(n3536) );
  XNOR U4022 ( .A(n3538), .B(n3539), .Z(n3476) );
  XNOR U4023 ( .A(n3540), .B(n3541), .Z(n3539) );
  OR U4024 ( .A(n3542), .B(n3543), .Z(n3541) );
  XNOR U4025 ( .A(n3493), .B(n3494), .Z(n3535) );
  XNOR U4026 ( .A(n191), .B(n194), .Z(n1680) );
  XOR U4027 ( .A(n3508), .B(n3527), .Z(n194) );
  XNOR U4028 ( .A(n3544), .B(n3545), .Z(n3508) );
  XNOR U4029 ( .A(n3546), .B(n3547), .Z(n3545) );
  NOR U4030 ( .A(n3548), .B(n3549), .Z(n3546) );
  IV U4031 ( .A(n3359), .Z(n196) );
  XNOR U4032 ( .A(n3517), .B(n3524), .Z(n3359) );
  XNOR U4033 ( .A(n3550), .B(n3551), .Z(n3517) );
  XNOR U4034 ( .A(n3552), .B(n3553), .Z(n3551) );
  NOR U4035 ( .A(n3554), .B(n3555), .Z(n3552) );
  XNOR U4036 ( .A(n2150), .B(n3556), .Z(n3533) );
  XNOR U4037 ( .A(key[1230]), .B(n1677), .Z(n3556) );
  XOR U4038 ( .A(n3483), .B(n3557), .Z(n1677) );
  XOR U4039 ( .A(n3558), .B(n3559), .Z(n2150) );
  XOR U4040 ( .A(n224), .B(n3379), .Z(n3559) );
  XOR U4041 ( .A(n3537), .B(n3560), .Z(n3379) );
  XNOR U4042 ( .A(n3532), .B(n3494), .Z(n3560) );
  XNOR U4043 ( .A(n3561), .B(n3562), .Z(n3494) );
  XOR U4044 ( .A(n3563), .B(n3564), .Z(n3562) );
  NOR U4045 ( .A(n3565), .B(n3542), .Z(n3563) );
  IV U4046 ( .A(n3493), .Z(n3532) );
  XOR U4047 ( .A(n3566), .B(n3567), .Z(n3493) );
  XOR U4048 ( .A(n3568), .B(n3569), .Z(n3567) );
  ANDN U4049 ( .B(n3570), .A(n3482), .Z(n3568) );
  XOR U4050 ( .A(n3496), .B(n3531), .Z(n3537) );
  XNOR U4051 ( .A(n3571), .B(n3572), .Z(n224) );
  XOR U4052 ( .A(n3573), .B(n3530), .Z(n3572) );
  XOR U4053 ( .A(n203), .B(n3574), .Z(n3558) );
  XNOR U4054 ( .A(key[1224]), .B(n1692), .Z(n3574) );
  IV U4055 ( .A(n3483), .Z(n1692) );
  XNOR U4056 ( .A(n1690), .B(n234), .Z(n203) );
  IV U4057 ( .A(n3353), .Z(n234) );
  XOR U4058 ( .A(n3471), .B(n3498), .Z(n3353) );
  XOR U4059 ( .A(n3470), .B(n3501), .Z(n1690) );
  IV U4060 ( .A(n3466), .Z(n3486) );
  XNOR U4061 ( .A(n3575), .B(n3576), .Z(n3466) );
  XOR U4062 ( .A(n3356), .B(n3369), .Z(n3576) );
  IV U4063 ( .A(n1681), .Z(n3369) );
  XNOR U4064 ( .A(n3577), .B(n3578), .Z(n1681) );
  XOR U4065 ( .A(n3579), .B(n3580), .Z(n3578) );
  XNOR U4066 ( .A(n3471), .B(n3581), .Z(n3577) );
  XOR U4067 ( .A(n3553), .B(n3582), .Z(n3581) );
  ANDN U4068 ( .B(n3583), .A(n3584), .Z(n3582) );
  ANDN U4069 ( .B(n3585), .A(n3586), .Z(n3553) );
  XNOR U4070 ( .A(n3587), .B(n3588), .Z(n3471) );
  XOR U4071 ( .A(n3589), .B(n3590), .Z(n3588) );
  NOR U4072 ( .A(n3591), .B(n3555), .Z(n3589) );
  XOR U4073 ( .A(n3531), .B(n3592), .Z(n3356) );
  XOR U4074 ( .A(n3495), .B(n3496), .Z(n3592) );
  XOR U4075 ( .A(n3477), .B(n3593), .Z(n3496) );
  XNOR U4076 ( .A(n3564), .B(n3594), .Z(n3593) );
  NANDN U4077 ( .A(n3595), .B(n3596), .Z(n3594) );
  OR U4078 ( .A(n3597), .B(n3598), .Z(n3564) );
  XNOR U4079 ( .A(n3561), .B(n3599), .Z(n3495) );
  XNOR U4080 ( .A(n3600), .B(n3479), .Z(n3599) );
  NOR U4081 ( .A(n3601), .B(n3602), .Z(n3479) );
  NOR U4082 ( .A(n3603), .B(n3604), .Z(n3600) );
  XNOR U4083 ( .A(n3477), .B(n3605), .Z(n3561) );
  XNOR U4084 ( .A(n3606), .B(n3607), .Z(n3605) );
  NANDN U4085 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U4086 ( .A(n3610), .B(n3606), .Z(n3477) );
  OR U4087 ( .A(n3611), .B(n3612), .Z(n3606) );
  ANDN U4088 ( .B(n3613), .A(n3614), .Z(n3610) );
  XNOR U4089 ( .A(n191), .B(n3615), .Z(n3575) );
  XNOR U4090 ( .A(key[1229]), .B(n3360), .Z(n3615) );
  XNOR U4091 ( .A(n1683), .B(n198), .Z(n3360) );
  XOR U4092 ( .A(n3616), .B(n3617), .Z(n198) );
  XOR U4093 ( .A(n3618), .B(n3619), .Z(n3617) );
  XNOR U4094 ( .A(n3514), .B(n3620), .Z(n3616) );
  XNOR U4095 ( .A(n3621), .B(n3622), .Z(n3620) );
  ANDN U4096 ( .B(n3623), .A(n3624), .Z(n3621) );
  XOR U4097 ( .A(n3625), .B(n3626), .Z(n1683) );
  XOR U4098 ( .A(n3627), .B(n3628), .Z(n3626) );
  XNOR U4099 ( .A(n3470), .B(n3629), .Z(n3625) );
  XOR U4100 ( .A(n3547), .B(n3630), .Z(n3629) );
  ANDN U4101 ( .B(n3631), .A(n3632), .Z(n3630) );
  ANDN U4102 ( .B(n3633), .A(n3634), .Z(n3547) );
  XNOR U4103 ( .A(n3635), .B(n3636), .Z(n3470) );
  XOR U4104 ( .A(n3637), .B(n3638), .Z(n3636) );
  NOR U4105 ( .A(n3639), .B(n3549), .Z(n3637) );
  XOR U4106 ( .A(n3513), .B(n3640), .Z(n191) );
  XNOR U4107 ( .A(n3512), .B(n3529), .Z(n3640) );
  XNOR U4108 ( .A(n3641), .B(n3642), .Z(n3512) );
  XNOR U4109 ( .A(n3622), .B(n3643), .Z(n3642) );
  OR U4110 ( .A(n3644), .B(n3645), .Z(n3643) );
  NANDN U4111 ( .A(n3646), .B(n3647), .Z(n3622) );
  XOR U4112 ( .A(n3648), .B(n3649), .Z(n3461) );
  XNOR U4113 ( .A(n232), .B(n1689), .Z(n3649) );
  XNOR U4114 ( .A(n3650), .B(n3516), .Z(n1689) );
  XNOR U4115 ( .A(n3499), .B(n3522), .Z(n3516) );
  XNOR U4116 ( .A(n3550), .B(n3651), .Z(n3522) );
  XNOR U4117 ( .A(n3652), .B(n3653), .Z(n3651) );
  NANDN U4118 ( .A(n3654), .B(n3655), .Z(n3653) );
  XNOR U4119 ( .A(n3656), .B(n3657), .Z(n3550) );
  XNOR U4120 ( .A(n3658), .B(n3659), .Z(n3657) );
  NANDN U4121 ( .A(n3660), .B(n3661), .Z(n3659) );
  XNOR U4122 ( .A(n3662), .B(n3663), .Z(n3499) );
  XNOR U4123 ( .A(n3590), .B(n3664), .Z(n3663) );
  NANDN U4124 ( .A(n3665), .B(n3583), .Z(n3664) );
  XNOR U4125 ( .A(n3555), .B(n3583), .Z(n3585) );
  XNOR U4126 ( .A(n3580), .B(n3524), .Z(n3650) );
  XOR U4127 ( .A(n3498), .B(n3518), .Z(n3524) );
  XNOR U4128 ( .A(n3656), .B(n3667), .Z(n3518) );
  XNOR U4129 ( .A(n3652), .B(n3668), .Z(n3667) );
  NANDN U4130 ( .A(n3669), .B(n3670), .Z(n3668) );
  OR U4131 ( .A(n3671), .B(n3672), .Z(n3652) );
  IV U4132 ( .A(n3579), .Z(n3656) );
  XNOR U4133 ( .A(n3673), .B(n3658), .Z(n3579) );
  NANDN U4134 ( .A(n3674), .B(n3675), .Z(n3658) );
  ANDN U4135 ( .B(n3676), .A(n3677), .Z(n3673) );
  XNOR U4136 ( .A(n3662), .B(n3678), .Z(n3498) );
  XOR U4137 ( .A(n3679), .B(n3680), .Z(n3678) );
  ANDN U4138 ( .B(n3670), .A(n3681), .Z(n3679) );
  XNOR U4139 ( .A(n3587), .B(n3682), .Z(n3580) );
  XNOR U4140 ( .A(n3680), .B(n3683), .Z(n3682) );
  NANDN U4141 ( .A(n3684), .B(n3655), .Z(n3683) );
  OR U4142 ( .A(n3671), .B(n3685), .Z(n3680) );
  XNOR U4143 ( .A(n3655), .B(n3670), .Z(n3671) );
  XNOR U4144 ( .A(n3662), .B(n3686), .Z(n3587) );
  XNOR U4145 ( .A(n3687), .B(n3688), .Z(n3686) );
  NANDN U4146 ( .A(n3660), .B(n3689), .Z(n3688) );
  XOR U4147 ( .A(n3690), .B(n3687), .Z(n3662) );
  OR U4148 ( .A(n3674), .B(n3691), .Z(n3687) );
  XOR U4149 ( .A(n3692), .B(n3660), .Z(n3674) );
  XNOR U4150 ( .A(n3670), .B(n3583), .Z(n3660) );
  XOR U4151 ( .A(n3693), .B(n3694), .Z(n3583) );
  NANDN U4152 ( .A(n3695), .B(n3696), .Z(n3694) );
  XOR U4153 ( .A(n3697), .B(n3698), .Z(n3670) );
  NANDN U4154 ( .A(n3695), .B(n3699), .Z(n3698) );
  ANDN U4155 ( .B(n3692), .A(n3700), .Z(n3690) );
  IV U4156 ( .A(n3677), .Z(n3692) );
  XOR U4157 ( .A(n3555), .B(n3655), .Z(n3677) );
  XNOR U4158 ( .A(n3701), .B(n3697), .Z(n3655) );
  NANDN U4159 ( .A(n3702), .B(n3703), .Z(n3697) );
  XOR U4160 ( .A(n3699), .B(n3704), .Z(n3703) );
  ANDN U4161 ( .B(n3704), .A(n3705), .Z(n3701) );
  XOR U4162 ( .A(n3706), .B(n3693), .Z(n3555) );
  NANDN U4163 ( .A(n3702), .B(n3707), .Z(n3693) );
  XOR U4164 ( .A(n3708), .B(n3696), .Z(n3707) );
  XNOR U4165 ( .A(n3709), .B(n3710), .Z(n3695) );
  XOR U4166 ( .A(n3711), .B(n3712), .Z(n3710) );
  XNOR U4167 ( .A(n3713), .B(n3714), .Z(n3709) );
  XNOR U4168 ( .A(n3715), .B(n3716), .Z(n3714) );
  ANDN U4169 ( .B(n3708), .A(n3712), .Z(n3715) );
  ANDN U4170 ( .B(n3708), .A(n3705), .Z(n3706) );
  XNOR U4171 ( .A(n3711), .B(n3717), .Z(n3705) );
  XOR U4172 ( .A(n3718), .B(n3716), .Z(n3717) );
  NAND U4173 ( .A(n3719), .B(n3720), .Z(n3716) );
  XNOR U4174 ( .A(n3713), .B(n3696), .Z(n3720) );
  IV U4175 ( .A(n3708), .Z(n3713) );
  XNOR U4176 ( .A(n3699), .B(n3712), .Z(n3719) );
  IV U4177 ( .A(n3704), .Z(n3712) );
  XOR U4178 ( .A(n3721), .B(n3722), .Z(n3704) );
  XNOR U4179 ( .A(n3723), .B(n3724), .Z(n3722) );
  XNOR U4180 ( .A(n3725), .B(n3726), .Z(n3721) );
  NOR U4181 ( .A(n3554), .B(n3591), .Z(n3725) );
  AND U4182 ( .A(n3696), .B(n3699), .Z(n3718) );
  XNOR U4183 ( .A(n3696), .B(n3699), .Z(n3711) );
  XNOR U4184 ( .A(n3727), .B(n3728), .Z(n3699) );
  XNOR U4185 ( .A(n3729), .B(n3724), .Z(n3728) );
  XOR U4186 ( .A(n3730), .B(n3731), .Z(n3727) );
  XNOR U4187 ( .A(n3732), .B(n3726), .Z(n3731) );
  OR U4188 ( .A(n3586), .B(n3666), .Z(n3726) );
  XNOR U4189 ( .A(n3591), .B(n3665), .Z(n3666) );
  XNOR U4190 ( .A(n3554), .B(n3584), .Z(n3586) );
  ANDN U4191 ( .B(n3733), .A(n3665), .Z(n3732) );
  XNOR U4192 ( .A(n3734), .B(n3735), .Z(n3696) );
  XNOR U4193 ( .A(n3724), .B(n3736), .Z(n3735) );
  XOR U4194 ( .A(n3654), .B(n3730), .Z(n3736) );
  XNOR U4195 ( .A(n3591), .B(n3737), .Z(n3724) );
  XOR U4196 ( .A(n3684), .B(n3738), .Z(n3734) );
  XNOR U4197 ( .A(n3739), .B(n3740), .Z(n3738) );
  ANDN U4198 ( .B(n3741), .A(n3681), .Z(n3739) );
  XNOR U4199 ( .A(n3742), .B(n3743), .Z(n3708) );
  XNOR U4200 ( .A(n3729), .B(n3744), .Z(n3743) );
  XNOR U4201 ( .A(n3669), .B(n3723), .Z(n3744) );
  XOR U4202 ( .A(n3730), .B(n3745), .Z(n3723) );
  XNOR U4203 ( .A(n3746), .B(n3747), .Z(n3745) );
  NAND U4204 ( .A(n3689), .B(n3661), .Z(n3747) );
  XNOR U4205 ( .A(n3748), .B(n3746), .Z(n3730) );
  NANDN U4206 ( .A(n3691), .B(n3675), .Z(n3746) );
  XOR U4207 ( .A(n3676), .B(n3661), .Z(n3675) );
  XNOR U4208 ( .A(n3741), .B(n3584), .Z(n3661) );
  XOR U4209 ( .A(n3700), .B(n3689), .Z(n3691) );
  XNOR U4210 ( .A(n3681), .B(n3749), .Z(n3689) );
  ANDN U4211 ( .B(n3676), .A(n3700), .Z(n3748) );
  XNOR U4212 ( .A(n3684), .B(n3591), .Z(n3700) );
  XOR U4213 ( .A(n3750), .B(n3751), .Z(n3591) );
  XNOR U4214 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U4215 ( .A(n3749), .B(n3733), .Z(n3729) );
  IV U4216 ( .A(n3584), .Z(n3733) );
  XOR U4217 ( .A(n3754), .B(n3755), .Z(n3584) );
  XNOR U4218 ( .A(n3756), .B(n3753), .Z(n3755) );
  IV U4219 ( .A(n3665), .Z(n3749) );
  XOR U4220 ( .A(n3753), .B(n3757), .Z(n3665) );
  XNOR U4221 ( .A(n3758), .B(n3759), .Z(n3742) );
  XNOR U4222 ( .A(n3760), .B(n3740), .Z(n3759) );
  OR U4223 ( .A(n3672), .B(n3685), .Z(n3740) );
  XNOR U4224 ( .A(n3684), .B(n3681), .Z(n3685) );
  IV U4225 ( .A(n3758), .Z(n3681) );
  XOR U4226 ( .A(n3654), .B(n3741), .Z(n3672) );
  IV U4227 ( .A(n3669), .Z(n3741) );
  XOR U4228 ( .A(n3737), .B(n3761), .Z(n3669) );
  XNOR U4229 ( .A(n3756), .B(n3750), .Z(n3761) );
  XOR U4230 ( .A(n3762), .B(n3763), .Z(n3750) );
  XNOR U4231 ( .A(n2779), .B(n3764), .Z(n3763) );
  XNOR U4232 ( .A(key[1074]), .B(n2821), .Z(n3762) );
  IV U4233 ( .A(n3554), .Z(n3737) );
  XOR U4234 ( .A(n3754), .B(n3765), .Z(n3554) );
  XOR U4235 ( .A(n3753), .B(n3766), .Z(n3765) );
  NOR U4236 ( .A(n3654), .B(n3684), .Z(n3760) );
  XOR U4237 ( .A(n3754), .B(n3767), .Z(n3654) );
  XOR U4238 ( .A(n3753), .B(n3768), .Z(n3767) );
  XOR U4239 ( .A(n3769), .B(n3770), .Z(n3753) );
  XOR U4240 ( .A(n2797), .B(n3771), .Z(n3770) );
  XNOR U4241 ( .A(n2792), .B(n3772), .Z(n3769) );
  XOR U4242 ( .A(key[1078]), .B(n3684), .Z(n3772) );
  XNOR U4243 ( .A(n3773), .B(n3774), .Z(n2792) );
  IV U4244 ( .A(n3757), .Z(n3754) );
  XOR U4245 ( .A(n3775), .B(n3776), .Z(n3757) );
  XNOR U4246 ( .A(n2796), .B(n3777), .Z(n3776) );
  XNOR U4247 ( .A(n3778), .B(n3779), .Z(n2796) );
  XNOR U4248 ( .A(key[1077]), .B(n3780), .Z(n3775) );
  XOR U4249 ( .A(n3781), .B(n3782), .Z(n3758) );
  XNOR U4250 ( .A(n3768), .B(n3766), .Z(n3782) );
  XNOR U4251 ( .A(n3783), .B(n3784), .Z(n3766) );
  XNOR U4252 ( .A(n3774), .B(n2805), .Z(n3784) );
  XOR U4253 ( .A(n3785), .B(n3786), .Z(n2805) );
  XNOR U4254 ( .A(n3787), .B(n3788), .Z(n3774) );
  XNOR U4255 ( .A(key[1079]), .B(n3789), .Z(n3783) );
  XNOR U4256 ( .A(n3790), .B(n3791), .Z(n3768) );
  XNOR U4257 ( .A(n2809), .B(n3792), .Z(n3791) );
  XOR U4258 ( .A(n3793), .B(n3794), .Z(n2809) );
  XNOR U4259 ( .A(n2811), .B(n3795), .Z(n3790) );
  XNOR U4260 ( .A(n3787), .B(n3780), .Z(n2811) );
  XNOR U4261 ( .A(n3684), .B(n3752), .Z(n3781) );
  XOR U4262 ( .A(n3797), .B(n3798), .Z(n3752) );
  XNOR U4263 ( .A(n3799), .B(n3800), .Z(n3798) );
  XNOR U4264 ( .A(n3756), .B(n2826), .Z(n3800) );
  XOR U4265 ( .A(n3787), .B(n3796), .Z(n2826) );
  XOR U4266 ( .A(n3801), .B(n3802), .Z(n3756) );
  XOR U4267 ( .A(n2823), .B(n3803), .Z(n3802) );
  XOR U4268 ( .A(key[1073]), .B(n2835), .Z(n3801) );
  XNOR U4269 ( .A(n2780), .B(n3804), .Z(n3797) );
  XNOR U4270 ( .A(key[1075]), .B(n3805), .Z(n3804) );
  XNOR U4271 ( .A(n3806), .B(n3807), .Z(n3684) );
  XOR U4272 ( .A(n3808), .B(n2806), .Z(n3807) );
  IV U4273 ( .A(n3809), .Z(n2806) );
  XNOR U4274 ( .A(key[1072]), .B(n3810), .Z(n3806) );
  XOR U4275 ( .A(n3483), .B(n1711), .Z(n232) );
  XOR U4276 ( .A(n3531), .B(n3475), .Z(n1711) );
  XNOR U4277 ( .A(n3538), .B(n3811), .Z(n3475) );
  XNOR U4278 ( .A(n3569), .B(n3812), .Z(n3811) );
  OR U4279 ( .A(n3604), .B(n3813), .Z(n3812) );
  OR U4280 ( .A(n3814), .B(n3601), .Z(n3569) );
  XOR U4281 ( .A(n3604), .B(n3815), .Z(n3601) );
  XNOR U4282 ( .A(n3566), .B(n3816), .Z(n3538) );
  XNOR U4283 ( .A(n3817), .B(n3818), .Z(n3816) );
  NAND U4284 ( .A(n3609), .B(n3819), .Z(n3818) );
  XNOR U4285 ( .A(n3566), .B(n3820), .Z(n3531) );
  XOR U4286 ( .A(n3821), .B(n3540), .Z(n3820) );
  OR U4287 ( .A(n3822), .B(n3597), .Z(n3540) );
  XNOR U4288 ( .A(n3542), .B(n3595), .Z(n3597) );
  NOR U4289 ( .A(n3823), .B(n3595), .Z(n3821) );
  XOR U4290 ( .A(n3824), .B(n3817), .Z(n3566) );
  OR U4291 ( .A(n3611), .B(n3825), .Z(n3817) );
  XNOR U4292 ( .A(n3613), .B(n3609), .Z(n3611) );
  XOR U4293 ( .A(n3595), .B(n3482), .Z(n3609) );
  IV U4294 ( .A(n3815), .Z(n3482) );
  XOR U4295 ( .A(n3826), .B(n3827), .Z(n3815) );
  NANDN U4296 ( .A(n3828), .B(n3829), .Z(n3827) );
  XNOR U4297 ( .A(n3830), .B(n3831), .Z(n3595) );
  OR U4298 ( .A(n3828), .B(n3832), .Z(n3831) );
  XOR U4299 ( .A(n3542), .B(n3604), .Z(n3613) );
  XNOR U4300 ( .A(n3826), .B(n3834), .Z(n3604) );
  NANDN U4301 ( .A(n3835), .B(n3836), .Z(n3834) );
  NANDN U4302 ( .A(n3837), .B(n3838), .Z(n3826) );
  OR U4303 ( .A(n3840), .B(n3837), .Z(n3830) );
  XOR U4304 ( .A(n3841), .B(n3828), .Z(n3837) );
  XNOR U4305 ( .A(n3842), .B(n3843), .Z(n3828) );
  XOR U4306 ( .A(n3844), .B(n3836), .Z(n3843) );
  XNOR U4307 ( .A(n3845), .B(n3846), .Z(n3842) );
  XNOR U4308 ( .A(n3847), .B(n3848), .Z(n3846) );
  ANDN U4309 ( .B(n3836), .A(n3849), .Z(n3847) );
  IV U4310 ( .A(n3850), .Z(n3836) );
  ANDN U4311 ( .B(n3841), .A(n3849), .Z(n3839) );
  IV U4312 ( .A(n3835), .Z(n3841) );
  XNOR U4313 ( .A(n3844), .B(n3851), .Z(n3835) );
  XNOR U4314 ( .A(n3848), .B(n3852), .Z(n3851) );
  NANDN U4315 ( .A(n3832), .B(n3829), .Z(n3852) );
  NANDN U4316 ( .A(n3840), .B(n3838), .Z(n3848) );
  XNOR U4317 ( .A(n3829), .B(n3850), .Z(n3838) );
  XOR U4318 ( .A(n3853), .B(n3854), .Z(n3850) );
  XOR U4319 ( .A(n3855), .B(n3856), .Z(n3854) );
  XOR U4320 ( .A(n3857), .B(n3858), .Z(n3856) );
  XOR U4321 ( .A(n3596), .B(n3859), .Z(n3853) );
  XNOR U4322 ( .A(n3860), .B(n3861), .Z(n3859) );
  ANDN U4323 ( .B(n3862), .A(n3543), .Z(n3860) );
  XNOR U4324 ( .A(n3849), .B(n3832), .Z(n3840) );
  IV U4325 ( .A(n3845), .Z(n3849) );
  XOR U4326 ( .A(n3863), .B(n3864), .Z(n3845) );
  XNOR U4327 ( .A(n3865), .B(n3858), .Z(n3864) );
  XOR U4328 ( .A(n3866), .B(n3867), .Z(n3858) );
  XNOR U4329 ( .A(n3868), .B(n3869), .Z(n3867) );
  NANDN U4330 ( .A(n3608), .B(n3819), .Z(n3869) );
  XNOR U4331 ( .A(n3870), .B(n3871), .Z(n3863) );
  NOR U4332 ( .A(n3603), .B(n3813), .Z(n3870) );
  XOR U4333 ( .A(n3832), .B(n3829), .Z(n3844) );
  XNOR U4334 ( .A(n3872), .B(n3873), .Z(n3829) );
  XNOR U4335 ( .A(n3866), .B(n3874), .Z(n3873) );
  XNOR U4336 ( .A(n3862), .B(n3865), .Z(n3874) );
  XNOR U4337 ( .A(n3875), .B(n3876), .Z(n3872) );
  XNOR U4338 ( .A(n3877), .B(n3861), .Z(n3876) );
  OR U4339 ( .A(n3598), .B(n3822), .Z(n3861) );
  XNOR U4340 ( .A(n3875), .B(n3857), .Z(n3822) );
  XNOR U4341 ( .A(n3862), .B(n3596), .Z(n3598) );
  ANDN U4342 ( .B(n3596), .A(n3823), .Z(n3877) );
  IV U4343 ( .A(n3857), .Z(n3823) );
  XOR U4344 ( .A(n3878), .B(n3879), .Z(n3832) );
  XOR U4345 ( .A(n3866), .B(n3855), .Z(n3879) );
  XNOR U4346 ( .A(n3481), .B(n3570), .Z(n3855) );
  XOR U4347 ( .A(n3880), .B(n3868), .Z(n3866) );
  OR U4348 ( .A(n3825), .B(n3612), .Z(n3868) );
  XOR U4349 ( .A(n3881), .B(n3608), .Z(n3612) );
  XNOR U4350 ( .A(n3596), .B(n3481), .Z(n3608) );
  XOR U4351 ( .A(n3882), .B(n3883), .Z(n3596) );
  XOR U4352 ( .A(n3603), .B(n3884), .Z(n3883) );
  XNOR U4353 ( .A(n3833), .B(n3819), .Z(n3825) );
  XOR U4354 ( .A(n3570), .B(n3857), .Z(n3819) );
  XOR U4355 ( .A(n3885), .B(n3886), .Z(n3857) );
  XNOR U4356 ( .A(n3887), .B(n3888), .Z(n3886) );
  XOR U4357 ( .A(n3889), .B(n3875), .Z(n3885) );
  ANDN U4358 ( .B(n3833), .A(n3614), .Z(n3880) );
  IV U4359 ( .A(n3881), .Z(n3614) );
  XNOR U4360 ( .A(n3862), .B(n3603), .Z(n3881) );
  IV U4361 ( .A(n3565), .Z(n3862) );
  XNOR U4362 ( .A(n3890), .B(n3891), .Z(n3565) );
  XOR U4363 ( .A(n3892), .B(n3889), .Z(n3891) );
  XOR U4364 ( .A(n3893), .B(n3894), .Z(n3889) );
  XOR U4365 ( .A(n3895), .B(n2669), .Z(n3894) );
  XNOR U4366 ( .A(n3896), .B(n2666), .Z(n2669) );
  XNOR U4367 ( .A(key[1036]), .B(n3897), .Z(n3893) );
  XOR U4368 ( .A(n3865), .B(n3898), .Z(n3878) );
  XNOR U4369 ( .A(n3899), .B(n3871), .Z(n3898) );
  OR U4370 ( .A(n3602), .B(n3814), .Z(n3871) );
  XOR U4371 ( .A(n3813), .B(n3570), .Z(n3814) );
  XOR U4372 ( .A(n3603), .B(n3481), .Z(n3602) );
  AND U4373 ( .A(n3570), .B(n3481), .Z(n3899) );
  XOR U4374 ( .A(n3882), .B(n3900), .Z(n3481) );
  XOR U4375 ( .A(n3892), .B(n3890), .Z(n3570) );
  XNOR U4376 ( .A(n3887), .B(n3900), .Z(n3603) );
  XNOR U4377 ( .A(n3901), .B(n3902), .Z(n3892) );
  XOR U4378 ( .A(n3903), .B(n3904), .Z(n3902) );
  XNOR U4379 ( .A(n3905), .B(n3906), .Z(n3901) );
  XNOR U4380 ( .A(key[1037]), .B(n3907), .Z(n3906) );
  XOR U4381 ( .A(n3908), .B(n3909), .Z(n3887) );
  XNOR U4382 ( .A(n3910), .B(n3911), .Z(n3909) );
  XNOR U4383 ( .A(key[1039]), .B(n3912), .Z(n3908) );
  XOR U4384 ( .A(n3543), .B(n3813), .Z(n3833) );
  XOR U4385 ( .A(n3888), .B(n3913), .Z(n3813) );
  XOR U4386 ( .A(n3890), .B(n3884), .Z(n3913) );
  XNOR U4387 ( .A(n3914), .B(n3915), .Z(n3884) );
  XOR U4388 ( .A(n3916), .B(n2681), .Z(n3915) );
  XNOR U4389 ( .A(n3917), .B(n3918), .Z(n3914) );
  XOR U4390 ( .A(key[1034]), .B(n3919), .Z(n3918) );
  XOR U4391 ( .A(n3920), .B(n3921), .Z(n3890) );
  XNOR U4392 ( .A(n2654), .B(n3922), .Z(n3921) );
  XOR U4393 ( .A(n3923), .B(n3924), .Z(n2654) );
  XNOR U4394 ( .A(n3875), .B(n3925), .Z(n3920) );
  XOR U4395 ( .A(key[1038]), .B(n3926), .Z(n3925) );
  XOR U4396 ( .A(n3927), .B(n3928), .Z(n3888) );
  XNOR U4397 ( .A(n2682), .B(n3929), .Z(n3928) );
  XOR U4398 ( .A(n3930), .B(n3931), .Z(n3929) );
  XNOR U4399 ( .A(n3932), .B(n2666), .Z(n2682) );
  XNOR U4400 ( .A(n3933), .B(n3934), .Z(n3927) );
  XNOR U4401 ( .A(key[1035]), .B(n3882), .Z(n3934) );
  XOR U4402 ( .A(n3935), .B(n3936), .Z(n3882) );
  XOR U4403 ( .A(n2688), .B(n3937), .Z(n3936) );
  XOR U4404 ( .A(n3938), .B(n3939), .Z(n3935) );
  XOR U4405 ( .A(key[1033]), .B(n3940), .Z(n3939) );
  IV U4406 ( .A(n3875), .Z(n3543) );
  XOR U4407 ( .A(n3941), .B(n3942), .Z(n3875) );
  XNOR U4408 ( .A(n3943), .B(n3944), .Z(n3942) );
  XNOR U4409 ( .A(key[1032]), .B(n2666), .Z(n3945) );
  XOR U4410 ( .A(n3514), .B(n3529), .Z(n3483) );
  XNOR U4411 ( .A(n3946), .B(n3947), .Z(n3514) );
  XOR U4412 ( .A(n3948), .B(n3949), .Z(n3947) );
  NOR U4413 ( .A(n3950), .B(n3644), .Z(n3948) );
  XNOR U4414 ( .A(key[1231]), .B(n3366), .Z(n3648) );
  XOR U4415 ( .A(n3557), .B(n1691), .Z(n3366) );
  XNOR U4416 ( .A(n3951), .B(n3507), .Z(n1691) );
  XNOR U4417 ( .A(n3502), .B(n3525), .Z(n3507) );
  XNOR U4418 ( .A(n3544), .B(n3952), .Z(n3525) );
  XNOR U4419 ( .A(n3953), .B(n3954), .Z(n3952) );
  NANDN U4420 ( .A(n3955), .B(n3956), .Z(n3954) );
  XNOR U4421 ( .A(n3957), .B(n3958), .Z(n3544) );
  XNOR U4422 ( .A(n3959), .B(n3960), .Z(n3958) );
  NANDN U4423 ( .A(n3961), .B(n3962), .Z(n3960) );
  XNOR U4424 ( .A(n3963), .B(n3964), .Z(n3502) );
  XNOR U4425 ( .A(n3638), .B(n3965), .Z(n3964) );
  NANDN U4426 ( .A(n3966), .B(n3631), .Z(n3965) );
  XNOR U4427 ( .A(n3549), .B(n3631), .Z(n3633) );
  XNOR U4428 ( .A(n3628), .B(n3527), .Z(n3951) );
  XOR U4429 ( .A(n3501), .B(n3509), .Z(n3527) );
  XNOR U4430 ( .A(n3957), .B(n3968), .Z(n3509) );
  XNOR U4431 ( .A(n3953), .B(n3969), .Z(n3968) );
  NANDN U4432 ( .A(n3970), .B(n3971), .Z(n3969) );
  OR U4433 ( .A(n3972), .B(n3973), .Z(n3953) );
  IV U4434 ( .A(n3627), .Z(n3957) );
  XNOR U4435 ( .A(n3974), .B(n3959), .Z(n3627) );
  NANDN U4436 ( .A(n3975), .B(n3976), .Z(n3959) );
  ANDN U4437 ( .B(n3977), .A(n3978), .Z(n3974) );
  XNOR U4438 ( .A(n3963), .B(n3979), .Z(n3501) );
  XOR U4439 ( .A(n3980), .B(n3981), .Z(n3979) );
  ANDN U4440 ( .B(n3971), .A(n3982), .Z(n3980) );
  XNOR U4441 ( .A(n3635), .B(n3983), .Z(n3628) );
  XNOR U4442 ( .A(n3981), .B(n3984), .Z(n3983) );
  NANDN U4443 ( .A(n3985), .B(n3956), .Z(n3984) );
  OR U4444 ( .A(n3972), .B(n3986), .Z(n3981) );
  XNOR U4445 ( .A(n3956), .B(n3971), .Z(n3972) );
  XNOR U4446 ( .A(n3963), .B(n3987), .Z(n3635) );
  XNOR U4447 ( .A(n3988), .B(n3989), .Z(n3987) );
  NANDN U4448 ( .A(n3961), .B(n3990), .Z(n3989) );
  XOR U4449 ( .A(n3991), .B(n3988), .Z(n3963) );
  OR U4450 ( .A(n3975), .B(n3992), .Z(n3988) );
  XOR U4451 ( .A(n3993), .B(n3961), .Z(n3975) );
  XNOR U4452 ( .A(n3971), .B(n3631), .Z(n3961) );
  XOR U4453 ( .A(n3994), .B(n3995), .Z(n3631) );
  NANDN U4454 ( .A(n3996), .B(n3997), .Z(n3995) );
  XOR U4455 ( .A(n3998), .B(n3999), .Z(n3971) );
  NANDN U4456 ( .A(n3996), .B(n4000), .Z(n3999) );
  ANDN U4457 ( .B(n3993), .A(n4001), .Z(n3991) );
  IV U4458 ( .A(n3978), .Z(n3993) );
  XOR U4459 ( .A(n3549), .B(n3956), .Z(n3978) );
  XNOR U4460 ( .A(n4002), .B(n3998), .Z(n3956) );
  NANDN U4461 ( .A(n4003), .B(n4004), .Z(n3998) );
  XOR U4462 ( .A(n4000), .B(n4005), .Z(n4004) );
  ANDN U4463 ( .B(n4005), .A(n4006), .Z(n4002) );
  XOR U4464 ( .A(n4007), .B(n3994), .Z(n3549) );
  NANDN U4465 ( .A(n4003), .B(n4008), .Z(n3994) );
  XOR U4466 ( .A(n4009), .B(n3997), .Z(n4008) );
  XNOR U4467 ( .A(n4010), .B(n4011), .Z(n3996) );
  XOR U4468 ( .A(n4012), .B(n4013), .Z(n4011) );
  XNOR U4469 ( .A(n4014), .B(n4015), .Z(n4010) );
  XNOR U4470 ( .A(n4016), .B(n4017), .Z(n4015) );
  ANDN U4471 ( .B(n4009), .A(n4013), .Z(n4016) );
  ANDN U4472 ( .B(n4009), .A(n4006), .Z(n4007) );
  XNOR U4473 ( .A(n4012), .B(n4018), .Z(n4006) );
  XOR U4474 ( .A(n4019), .B(n4017), .Z(n4018) );
  NAND U4475 ( .A(n4020), .B(n4021), .Z(n4017) );
  XNOR U4476 ( .A(n4014), .B(n3997), .Z(n4021) );
  IV U4477 ( .A(n4009), .Z(n4014) );
  XNOR U4478 ( .A(n4000), .B(n4013), .Z(n4020) );
  IV U4479 ( .A(n4005), .Z(n4013) );
  XOR U4480 ( .A(n4022), .B(n4023), .Z(n4005) );
  XNOR U4481 ( .A(n4024), .B(n4025), .Z(n4023) );
  XNOR U4482 ( .A(n4026), .B(n4027), .Z(n4022) );
  NOR U4483 ( .A(n3548), .B(n3639), .Z(n4026) );
  AND U4484 ( .A(n3997), .B(n4000), .Z(n4019) );
  XNOR U4485 ( .A(n3997), .B(n4000), .Z(n4012) );
  XNOR U4486 ( .A(n4028), .B(n4029), .Z(n4000) );
  XNOR U4487 ( .A(n4030), .B(n4025), .Z(n4029) );
  XOR U4488 ( .A(n4031), .B(n4032), .Z(n4028) );
  XNOR U4489 ( .A(n4033), .B(n4027), .Z(n4032) );
  OR U4490 ( .A(n3634), .B(n3967), .Z(n4027) );
  XNOR U4491 ( .A(n3639), .B(n3966), .Z(n3967) );
  XNOR U4492 ( .A(n3548), .B(n3632), .Z(n3634) );
  ANDN U4493 ( .B(n4034), .A(n3966), .Z(n4033) );
  XNOR U4494 ( .A(n4035), .B(n4036), .Z(n3997) );
  XNOR U4495 ( .A(n4025), .B(n4037), .Z(n4036) );
  XOR U4496 ( .A(n3955), .B(n4031), .Z(n4037) );
  XNOR U4497 ( .A(n3639), .B(n4038), .Z(n4025) );
  XOR U4498 ( .A(n3985), .B(n4039), .Z(n4035) );
  XNOR U4499 ( .A(n4040), .B(n4041), .Z(n4039) );
  ANDN U4500 ( .B(n4042), .A(n3982), .Z(n4040) );
  XNOR U4501 ( .A(n4043), .B(n4044), .Z(n4009) );
  XNOR U4502 ( .A(n4030), .B(n4045), .Z(n4044) );
  XNOR U4503 ( .A(n3970), .B(n4024), .Z(n4045) );
  XOR U4504 ( .A(n4031), .B(n4046), .Z(n4024) );
  XNOR U4505 ( .A(n4047), .B(n4048), .Z(n4046) );
  NAND U4506 ( .A(n3990), .B(n3962), .Z(n4048) );
  XNOR U4507 ( .A(n4049), .B(n4047), .Z(n4031) );
  NANDN U4508 ( .A(n3992), .B(n3976), .Z(n4047) );
  XOR U4509 ( .A(n3977), .B(n3962), .Z(n3976) );
  XNOR U4510 ( .A(n4042), .B(n3632), .Z(n3962) );
  XOR U4511 ( .A(n4001), .B(n3990), .Z(n3992) );
  XNOR U4512 ( .A(n3982), .B(n4050), .Z(n3990) );
  ANDN U4513 ( .B(n3977), .A(n4001), .Z(n4049) );
  XNOR U4514 ( .A(n3985), .B(n3639), .Z(n4001) );
  XOR U4515 ( .A(n4051), .B(n4052), .Z(n3639) );
  XNOR U4516 ( .A(n4053), .B(n4054), .Z(n4052) );
  XOR U4517 ( .A(n4050), .B(n4034), .Z(n4030) );
  IV U4518 ( .A(n3632), .Z(n4034) );
  XOR U4519 ( .A(n4055), .B(n4056), .Z(n3632) );
  XNOR U4520 ( .A(n4057), .B(n4054), .Z(n4056) );
  IV U4521 ( .A(n3966), .Z(n4050) );
  XOR U4522 ( .A(n4054), .B(n4058), .Z(n3966) );
  XNOR U4523 ( .A(n4059), .B(n4060), .Z(n4043) );
  XNOR U4524 ( .A(n4061), .B(n4041), .Z(n4060) );
  OR U4525 ( .A(n3973), .B(n3986), .Z(n4041) );
  XNOR U4526 ( .A(n3985), .B(n3982), .Z(n3986) );
  IV U4527 ( .A(n4059), .Z(n3982) );
  XOR U4528 ( .A(n3955), .B(n4042), .Z(n3973) );
  IV U4529 ( .A(n3970), .Z(n4042) );
  XOR U4530 ( .A(n4038), .B(n4062), .Z(n3970) );
  XNOR U4531 ( .A(n4057), .B(n4051), .Z(n4062) );
  XOR U4532 ( .A(n4063), .B(n4064), .Z(n4051) );
  XNOR U4533 ( .A(n4065), .B(n4066), .Z(n4064) );
  XNOR U4534 ( .A(n4067), .B(n4068), .Z(n4063) );
  XNOR U4535 ( .A(key[1114]), .B(n4069), .Z(n4068) );
  IV U4536 ( .A(n3548), .Z(n4038) );
  XOR U4537 ( .A(n4055), .B(n4070), .Z(n3548) );
  XOR U4538 ( .A(n4054), .B(n4071), .Z(n4070) );
  NOR U4539 ( .A(n3955), .B(n3985), .Z(n4061) );
  XOR U4540 ( .A(n4055), .B(n4072), .Z(n3955) );
  XOR U4541 ( .A(n4054), .B(n4073), .Z(n4072) );
  XOR U4542 ( .A(n4074), .B(n4075), .Z(n4054) );
  XNOR U4543 ( .A(n3125), .B(n4076), .Z(n4075) );
  XOR U4544 ( .A(n4077), .B(n4078), .Z(n3125) );
  XNOR U4545 ( .A(n4079), .B(n4080), .Z(n4074) );
  XOR U4546 ( .A(key[1118]), .B(n3985), .Z(n4080) );
  IV U4547 ( .A(n4058), .Z(n4055) );
  XOR U4548 ( .A(n4081), .B(n4082), .Z(n4058) );
  XOR U4549 ( .A(n4083), .B(n4084), .Z(n4082) );
  XNOR U4550 ( .A(n4085), .B(n4086), .Z(n4081) );
  XOR U4551 ( .A(key[1117]), .B(n4087), .Z(n4086) );
  XOR U4552 ( .A(n4088), .B(n4089), .Z(n4059) );
  XNOR U4553 ( .A(n4073), .B(n4071), .Z(n4089) );
  XNOR U4554 ( .A(n4090), .B(n4091), .Z(n4071) );
  XNOR U4555 ( .A(n4092), .B(n4093), .Z(n4091) );
  XNOR U4556 ( .A(key[1119]), .B(n4094), .Z(n4090) );
  XNOR U4557 ( .A(n4095), .B(n4096), .Z(n4073) );
  XOR U4558 ( .A(n4097), .B(n4098), .Z(n4096) );
  XNOR U4559 ( .A(n4099), .B(n4100), .Z(n4095) );
  XNOR U4560 ( .A(key[1116]), .B(n3142), .Z(n4100) );
  XOR U4561 ( .A(n3137), .B(n4101), .Z(n3142) );
  XNOR U4562 ( .A(n3985), .B(n4053), .Z(n4088) );
  XOR U4563 ( .A(n4102), .B(n4103), .Z(n4053) );
  XNOR U4564 ( .A(n4104), .B(n4105), .Z(n4103) );
  XNOR U4565 ( .A(n4057), .B(n4106), .Z(n4105) );
  XOR U4566 ( .A(n4107), .B(n4108), .Z(n4057) );
  XOR U4567 ( .A(n4109), .B(n3159), .Z(n4108) );
  XNOR U4568 ( .A(n4113), .B(n4114), .Z(n4102) );
  XNOR U4569 ( .A(key[1115]), .B(n3155), .Z(n4114) );
  XOR U4570 ( .A(n3137), .B(n4115), .Z(n3155) );
  XNOR U4571 ( .A(n4116), .B(n4117), .Z(n3985) );
  XNOR U4572 ( .A(n4118), .B(n4119), .Z(n4117) );
  XNOR U4573 ( .A(n3160), .B(n4120), .Z(n4116) );
  XNOR U4574 ( .A(key[1112]), .B(n4077), .Z(n4120) );
  IV U4575 ( .A(n3137), .Z(n4077) );
  IV U4576 ( .A(n205), .Z(n3557) );
  XNOR U4577 ( .A(n4121), .B(n3511), .Z(n205) );
  XOR U4578 ( .A(n3530), .B(n3571), .Z(n3511) );
  XNOR U4579 ( .A(n3641), .B(n4122), .Z(n3571) );
  XNOR U4580 ( .A(n4123), .B(n4124), .Z(n4122) );
  OR U4581 ( .A(n4125), .B(n4126), .Z(n4124) );
  XNOR U4582 ( .A(n4127), .B(n4128), .Z(n3641) );
  XNOR U4583 ( .A(n4129), .B(n4130), .Z(n4128) );
  NANDN U4584 ( .A(n4131), .B(n4132), .Z(n4130) );
  XOR U4585 ( .A(n4133), .B(n4134), .Z(n3530) );
  XNOR U4586 ( .A(n3949), .B(n4135), .Z(n4134) );
  NAND U4587 ( .A(n4136), .B(n3623), .Z(n4135) );
  NANDN U4588 ( .A(n4137), .B(n3647), .Z(n3949) );
  XNOR U4589 ( .A(n3644), .B(n3623), .Z(n3647) );
  XOR U4590 ( .A(n3619), .B(n3573), .Z(n4121) );
  XOR U4591 ( .A(n3529), .B(n3513), .Z(n3573) );
  XOR U4592 ( .A(n4127), .B(n4138), .Z(n3513) );
  XOR U4593 ( .A(n4139), .B(n4123), .Z(n4138) );
  OR U4594 ( .A(n4140), .B(n4141), .Z(n4123) );
  AND U4595 ( .A(n4142), .B(n4143), .Z(n4139) );
  IV U4596 ( .A(n3618), .Z(n4127) );
  XNOR U4597 ( .A(n4144), .B(n4129), .Z(n3618) );
  NANDN U4598 ( .A(n4145), .B(n4146), .Z(n4129) );
  AND U4599 ( .A(n4147), .B(n4148), .Z(n4144) );
  XNOR U4600 ( .A(n4133), .B(n4149), .Z(n3529) );
  XOR U4601 ( .A(n4150), .B(n4151), .Z(n4149) );
  ANDN U4602 ( .B(n4143), .A(n4152), .Z(n4150) );
  XNOR U4603 ( .A(n3946), .B(n4153), .Z(n3619) );
  XNOR U4604 ( .A(n4151), .B(n4154), .Z(n4153) );
  OR U4605 ( .A(n4125), .B(n4155), .Z(n4154) );
  OR U4606 ( .A(n4156), .B(n4140), .Z(n4151) );
  XOR U4607 ( .A(n4125), .B(n4143), .Z(n4140) );
  XNOR U4608 ( .A(n4133), .B(n4157), .Z(n3946) );
  XNOR U4609 ( .A(n4158), .B(n4159), .Z(n4157) );
  NANDN U4610 ( .A(n4131), .B(n4160), .Z(n4159) );
  XOR U4611 ( .A(n4161), .B(n4158), .Z(n4133) );
  OR U4612 ( .A(n4145), .B(n4162), .Z(n4158) );
  XOR U4613 ( .A(n4147), .B(n4131), .Z(n4145) );
  XNOR U4614 ( .A(n4143), .B(n3623), .Z(n4131) );
  XOR U4615 ( .A(n4163), .B(n4164), .Z(n3623) );
  NANDN U4616 ( .A(n4165), .B(n4166), .Z(n4164) );
  XOR U4617 ( .A(n4167), .B(n4168), .Z(n4143) );
  OR U4618 ( .A(n4165), .B(n4169), .Z(n4168) );
  ANDN U4619 ( .B(n4147), .A(n4170), .Z(n4161) );
  XOR U4620 ( .A(n4125), .B(n3644), .Z(n4147) );
  XOR U4621 ( .A(n4171), .B(n4163), .Z(n3644) );
  NANDN U4622 ( .A(n4172), .B(n4173), .Z(n4163) );
  ANDN U4623 ( .B(n4174), .A(n4175), .Z(n4171) );
  NANDN U4624 ( .A(n4172), .B(n4177), .Z(n4167) );
  XOR U4625 ( .A(n4178), .B(n4165), .Z(n4172) );
  XNOR U4626 ( .A(n4179), .B(n4180), .Z(n4165) );
  XOR U4627 ( .A(n4181), .B(n4174), .Z(n4180) );
  XNOR U4628 ( .A(n4182), .B(n4183), .Z(n4179) );
  XNOR U4629 ( .A(n4184), .B(n4185), .Z(n4183) );
  ANDN U4630 ( .B(n4174), .A(n4186), .Z(n4184) );
  IV U4631 ( .A(n4187), .Z(n4174) );
  ANDN U4632 ( .B(n4178), .A(n4186), .Z(n4176) );
  IV U4633 ( .A(n4182), .Z(n4186) );
  IV U4634 ( .A(n4175), .Z(n4178) );
  XNOR U4635 ( .A(n4181), .B(n4188), .Z(n4175) );
  XOR U4636 ( .A(n4189), .B(n4185), .Z(n4188) );
  NAND U4637 ( .A(n4177), .B(n4173), .Z(n4185) );
  XNOR U4638 ( .A(n4166), .B(n4187), .Z(n4173) );
  XOR U4639 ( .A(n4190), .B(n4191), .Z(n4187) );
  XOR U4640 ( .A(n4192), .B(n4193), .Z(n4191) );
  XNOR U4641 ( .A(n4142), .B(n4194), .Z(n4193) );
  XNOR U4642 ( .A(n4195), .B(n4196), .Z(n4190) );
  XNOR U4643 ( .A(n4197), .B(n4198), .Z(n4196) );
  ANDN U4644 ( .B(n4199), .A(n4155), .Z(n4197) );
  XNOR U4645 ( .A(n4182), .B(n4169), .Z(n4177) );
  XOR U4646 ( .A(n4200), .B(n4201), .Z(n4182) );
  XNOR U4647 ( .A(n4202), .B(n4194), .Z(n4201) );
  XOR U4648 ( .A(n4203), .B(n4204), .Z(n4194) );
  XNOR U4649 ( .A(n4205), .B(n4206), .Z(n4204) );
  NAND U4650 ( .A(n4160), .B(n4132), .Z(n4206) );
  XNOR U4651 ( .A(n4207), .B(n4208), .Z(n4200) );
  ANDN U4652 ( .B(n4209), .A(n3950), .Z(n4207) );
  ANDN U4653 ( .B(n4166), .A(n4169), .Z(n4189) );
  XOR U4654 ( .A(n4169), .B(n4166), .Z(n4181) );
  XNOR U4655 ( .A(n4210), .B(n4211), .Z(n4166) );
  XNOR U4656 ( .A(n4203), .B(n4212), .Z(n4211) );
  XOR U4657 ( .A(n4202), .B(n4126), .Z(n4212) );
  XOR U4658 ( .A(n4155), .B(n4213), .Z(n4210) );
  XNOR U4659 ( .A(n4214), .B(n4198), .Z(n4213) );
  OR U4660 ( .A(n4141), .B(n4156), .Z(n4198) );
  XNOR U4661 ( .A(n4155), .B(n4152), .Z(n4156) );
  XOR U4662 ( .A(n4126), .B(n4142), .Z(n4141) );
  ANDN U4663 ( .B(n4142), .A(n4152), .Z(n4214) );
  XOR U4664 ( .A(n4215), .B(n4216), .Z(n4169) );
  XOR U4665 ( .A(n4203), .B(n4192), .Z(n4216) );
  XOR U4666 ( .A(n4136), .B(n3624), .Z(n4192) );
  XOR U4667 ( .A(n4217), .B(n4205), .Z(n4203) );
  NANDN U4668 ( .A(n4162), .B(n4146), .Z(n4205) );
  XOR U4669 ( .A(n4148), .B(n4132), .Z(n4146) );
  XNOR U4670 ( .A(n4209), .B(n4218), .Z(n4142) );
  XOR U4671 ( .A(n4219), .B(n4220), .Z(n4218) );
  XOR U4672 ( .A(n4170), .B(n4160), .Z(n4162) );
  XNOR U4673 ( .A(n4152), .B(n4136), .Z(n4160) );
  IV U4674 ( .A(n4195), .Z(n4152) );
  XOR U4675 ( .A(n4221), .B(n4222), .Z(n4195) );
  XOR U4676 ( .A(n4223), .B(n4224), .Z(n4222) );
  XNOR U4677 ( .A(n4155), .B(n4225), .Z(n4221) );
  ANDN U4678 ( .B(n4148), .A(n4170), .Z(n4217) );
  XNOR U4679 ( .A(n4155), .B(n3950), .Z(n4170) );
  XOR U4680 ( .A(n4209), .B(n4199), .Z(n4148) );
  IV U4681 ( .A(n4126), .Z(n4199) );
  XOR U4682 ( .A(n4226), .B(n4227), .Z(n4126) );
  XOR U4683 ( .A(n4228), .B(n4224), .Z(n4227) );
  XNOR U4684 ( .A(n4229), .B(n4230), .Z(n4224) );
  XNOR U4685 ( .A(n4231), .B(n2970), .Z(n4230) );
  XNOR U4686 ( .A(n4232), .B(n4233), .Z(n2970) );
  XNOR U4687 ( .A(n2972), .B(n4234), .Z(n4229) );
  XOR U4688 ( .A(key[1124]), .B(n4235), .Z(n4234) );
  XOR U4689 ( .A(n4236), .B(n4237), .Z(n2972) );
  IV U4690 ( .A(n3645), .Z(n4209) );
  XOR U4691 ( .A(n4202), .B(n4238), .Z(n4215) );
  XNOR U4692 ( .A(n4239), .B(n4208), .Z(n4238) );
  OR U4693 ( .A(n3646), .B(n4137), .Z(n4208) );
  XNOR U4694 ( .A(n4240), .B(n4136), .Z(n4137) );
  XNOR U4695 ( .A(n3645), .B(n3624), .Z(n3646) );
  ANDN U4696 ( .B(n4136), .A(n3624), .Z(n4239) );
  XOR U4697 ( .A(n4226), .B(n4241), .Z(n3624) );
  XNOR U4698 ( .A(n4242), .B(n4228), .Z(n4241) );
  XOR U4699 ( .A(n4228), .B(n4226), .Z(n4136) );
  XNOR U4700 ( .A(n3950), .B(n3645), .Z(n4202) );
  XOR U4701 ( .A(n4226), .B(n4243), .Z(n3645) );
  XNOR U4702 ( .A(n4228), .B(n4223), .Z(n4243) );
  XOR U4703 ( .A(n4244), .B(n4245), .Z(n4223) );
  XNOR U4704 ( .A(n4246), .B(n2987), .Z(n4245) );
  XNOR U4705 ( .A(n4247), .B(n4248), .Z(n2987) );
  XOR U4706 ( .A(key[1127]), .B(n4249), .Z(n4244) );
  XNOR U4707 ( .A(n4250), .B(n4251), .Z(n4226) );
  XNOR U4708 ( .A(n2980), .B(n4252), .Z(n4251) );
  XNOR U4709 ( .A(n4253), .B(n4254), .Z(n2980) );
  XOR U4710 ( .A(key[1125]), .B(n4237), .Z(n4250) );
  IV U4711 ( .A(n4240), .Z(n3950) );
  XNOR U4712 ( .A(n4219), .B(n4225), .Z(n4255) );
  XOR U4713 ( .A(n4256), .B(n4257), .Z(n4225) );
  XOR U4714 ( .A(n3006), .B(n4258), .Z(n4257) );
  XOR U4715 ( .A(n4259), .B(n4220), .Z(n4258) );
  IV U4716 ( .A(n4242), .Z(n4220) );
  XOR U4717 ( .A(n4260), .B(n4261), .Z(n4242) );
  XNOR U4718 ( .A(n4262), .B(n3011), .Z(n4261) );
  XOR U4719 ( .A(key[1121]), .B(n3024), .Z(n4260) );
  XNOR U4720 ( .A(n3015), .B(n4263), .Z(n4256) );
  XNOR U4721 ( .A(key[1123]), .B(n2996), .Z(n4263) );
  XOR U4722 ( .A(n4236), .B(n4235), .Z(n3015) );
  XOR U4723 ( .A(n4264), .B(n4265), .Z(n4219) );
  XOR U4724 ( .A(n4266), .B(n2994), .Z(n4265) );
  XNOR U4725 ( .A(key[1122]), .B(n3012), .Z(n4264) );
  XOR U4726 ( .A(n4267), .B(n4268), .Z(n4228) );
  XOR U4727 ( .A(n4246), .B(n4269), .Z(n3002) );
  XOR U4728 ( .A(n4236), .B(n4270), .Z(n4246) );
  XNOR U4729 ( .A(n4271), .B(n4272), .Z(n4267) );
  XOR U4730 ( .A(key[1126]), .B(n4155), .Z(n4272) );
  XNOR U4731 ( .A(n4273), .B(n4274), .Z(n4155) );
  XOR U4732 ( .A(n2988), .B(n4275), .Z(n4274) );
  IV U4733 ( .A(n4276), .Z(n2988) );
  XNOR U4734 ( .A(key[1120]), .B(n4277), .Z(n4273) );
  XOR U4735 ( .A(n4278), .B(n4279), .Z(out[109]) );
  XNOR U4736 ( .A(n4280), .B(n4281), .Z(n4279) );
  XOR U4737 ( .A(n3387), .B(n4282), .Z(n4281) );
  XNOR U4738 ( .A(n4284), .B(n4285), .Z(n4283) );
  NANDN U4739 ( .A(n4286), .B(n4287), .Z(n4285) );
  XOR U4740 ( .A(n4289), .B(n4290), .Z(n4278) );
  XOR U4741 ( .A(key[1261]), .B(n4291), .Z(n4290) );
  ANDN U4742 ( .B(n4292), .A(n4293), .Z(n4289) );
  XNOR U4743 ( .A(n4294), .B(n4295), .Z(out[108]) );
  XNOR U4744 ( .A(key[1260]), .B(n4296), .Z(n4295) );
  XOR U4745 ( .A(n4297), .B(n4298), .Z(out[107]) );
  XNOR U4746 ( .A(n4299), .B(n3390), .Z(n4298) );
  XNOR U4747 ( .A(n4300), .B(n4301), .Z(n3390) );
  XNOR U4748 ( .A(n4302), .B(n4291), .Z(n4301) );
  ANDN U4749 ( .B(n4303), .A(n4304), .Z(n4291) );
  NOR U4750 ( .A(n4305), .B(n4306), .Z(n4302) );
  XNOR U4751 ( .A(n4307), .B(n4308), .Z(n4297) );
  XOR U4752 ( .A(key[1259]), .B(n4309), .Z(n4308) );
  XOR U4753 ( .A(key[1258]), .B(n4294), .Z(out[106]) );
  XNOR U4754 ( .A(n3389), .B(n4310), .Z(n4294) );
  IV U4755 ( .A(n4309), .Z(n3389) );
  XOR U4756 ( .A(n4311), .B(n3386), .Z(out[105]) );
  XNOR U4757 ( .A(n4300), .B(n4312), .Z(n4299) );
  XNOR U4758 ( .A(n4313), .B(n4314), .Z(n4312) );
  NANDN U4759 ( .A(n4315), .B(n4287), .Z(n4314) );
  XNOR U4760 ( .A(n4282), .B(n4316), .Z(n4300) );
  XNOR U4761 ( .A(n4317), .B(n4318), .Z(n4316) );
  NANDN U4762 ( .A(n4319), .B(n4320), .Z(n4318) );
  XOR U4763 ( .A(n4310), .B(n4307), .Z(n3392) );
  XNOR U4764 ( .A(n4282), .B(n4321), .Z(n4307) );
  XNOR U4765 ( .A(n4313), .B(n4322), .Z(n4321) );
  NANDN U4766 ( .A(n4323), .B(n4324), .Z(n4322) );
  OR U4767 ( .A(n4325), .B(n4326), .Z(n4313) );
  XOR U4768 ( .A(n4327), .B(n4317), .Z(n4282) );
  NANDN U4769 ( .A(n4328), .B(n4329), .Z(n4317) );
  ANDN U4770 ( .B(n4330), .A(n4331), .Z(n4327) );
  XOR U4771 ( .A(key[1257]), .B(n4309), .Z(n4311) );
  XOR U4772 ( .A(n4332), .B(n4333), .Z(n4309) );
  XNOR U4773 ( .A(n4334), .B(n4335), .Z(n4333) );
  NANDN U4774 ( .A(n4336), .B(n4292), .Z(n4335) );
  XNOR U4775 ( .A(n4280), .B(n4337), .Z(out[104]) );
  XOR U4776 ( .A(key[1256]), .B(n4310), .Z(n4337) );
  XNOR U4777 ( .A(n4332), .B(n4338), .Z(n4310) );
  XOR U4778 ( .A(n4339), .B(n4284), .Z(n4338) );
  OR U4779 ( .A(n4340), .B(n4325), .Z(n4284) );
  XNOR U4780 ( .A(n4287), .B(n4324), .Z(n4325) );
  ANDN U4781 ( .B(n4341), .A(n4342), .Z(n4339) );
  IV U4782 ( .A(n4296), .Z(n4280) );
  XOR U4783 ( .A(n4288), .B(n4343), .Z(n4296) );
  XOR U4784 ( .A(n4344), .B(n4334), .Z(n4343) );
  XNOR U4785 ( .A(n4306), .B(n4292), .Z(n4303) );
  NOR U4786 ( .A(n4346), .B(n4306), .Z(n4344) );
  XNOR U4787 ( .A(n4332), .B(n4347), .Z(n4288) );
  XNOR U4788 ( .A(n4348), .B(n4349), .Z(n4347) );
  NANDN U4789 ( .A(n4319), .B(n4350), .Z(n4349) );
  XOR U4790 ( .A(n4351), .B(n4348), .Z(n4332) );
  OR U4791 ( .A(n4328), .B(n4352), .Z(n4348) );
  XOR U4792 ( .A(n4353), .B(n4319), .Z(n4328) );
  XNOR U4793 ( .A(n4324), .B(n4292), .Z(n4319) );
  XOR U4794 ( .A(n4354), .B(n4355), .Z(n4292) );
  NANDN U4795 ( .A(n4356), .B(n4357), .Z(n4355) );
  IV U4796 ( .A(n4342), .Z(n4324) );
  XNOR U4797 ( .A(n4358), .B(n4359), .Z(n4342) );
  NANDN U4798 ( .A(n4356), .B(n4360), .Z(n4359) );
  ANDN U4799 ( .B(n4353), .A(n4361), .Z(n4351) );
  IV U4800 ( .A(n4331), .Z(n4353) );
  XOR U4801 ( .A(n4306), .B(n4287), .Z(n4331) );
  XNOR U4802 ( .A(n4362), .B(n4358), .Z(n4287) );
  NANDN U4803 ( .A(n4363), .B(n4364), .Z(n4358) );
  XOR U4804 ( .A(n4360), .B(n4365), .Z(n4364) );
  ANDN U4805 ( .B(n4365), .A(n4366), .Z(n4362) );
  XOR U4806 ( .A(n4367), .B(n4354), .Z(n4306) );
  NANDN U4807 ( .A(n4363), .B(n4368), .Z(n4354) );
  XOR U4808 ( .A(n4369), .B(n4357), .Z(n4368) );
  XNOR U4809 ( .A(n4370), .B(n4371), .Z(n4356) );
  XOR U4810 ( .A(n4372), .B(n4373), .Z(n4371) );
  XNOR U4811 ( .A(n4374), .B(n4375), .Z(n4370) );
  XNOR U4812 ( .A(n4376), .B(n4377), .Z(n4375) );
  ANDN U4813 ( .B(n4369), .A(n4373), .Z(n4376) );
  ANDN U4814 ( .B(n4369), .A(n4366), .Z(n4367) );
  XNOR U4815 ( .A(n4372), .B(n4378), .Z(n4366) );
  XOR U4816 ( .A(n4379), .B(n4377), .Z(n4378) );
  NAND U4817 ( .A(n4380), .B(n4381), .Z(n4377) );
  XNOR U4818 ( .A(n4374), .B(n4357), .Z(n4381) );
  IV U4819 ( .A(n4369), .Z(n4374) );
  XNOR U4820 ( .A(n4360), .B(n4373), .Z(n4380) );
  IV U4821 ( .A(n4365), .Z(n4373) );
  XOR U4822 ( .A(n4382), .B(n4383), .Z(n4365) );
  XNOR U4823 ( .A(n4384), .B(n4385), .Z(n4383) );
  XNOR U4824 ( .A(n4386), .B(n4387), .Z(n4382) );
  NOR U4825 ( .A(n4305), .B(n4346), .Z(n4386) );
  AND U4826 ( .A(n4357), .B(n4360), .Z(n4379) );
  XNOR U4827 ( .A(n4357), .B(n4360), .Z(n4372) );
  XNOR U4828 ( .A(n4388), .B(n4389), .Z(n4360) );
  XNOR U4829 ( .A(n4390), .B(n4385), .Z(n4389) );
  XOR U4830 ( .A(n4391), .B(n4392), .Z(n4388) );
  XNOR U4831 ( .A(n4393), .B(n4387), .Z(n4392) );
  OR U4832 ( .A(n4304), .B(n4345), .Z(n4387) );
  XNOR U4833 ( .A(n4346), .B(n4336), .Z(n4345) );
  XNOR U4834 ( .A(n4305), .B(n4293), .Z(n4304) );
  ANDN U4835 ( .B(n4394), .A(n4336), .Z(n4393) );
  XNOR U4836 ( .A(n4395), .B(n4396), .Z(n4357) );
  XNOR U4837 ( .A(n4385), .B(n4397), .Z(n4396) );
  XOR U4838 ( .A(n4315), .B(n4391), .Z(n4397) );
  XNOR U4839 ( .A(n4346), .B(n4398), .Z(n4385) );
  XNOR U4840 ( .A(n4399), .B(n4400), .Z(n4395) );
  XNOR U4841 ( .A(n4401), .B(n4402), .Z(n4400) );
  ANDN U4842 ( .B(n4341), .A(n4323), .Z(n4401) );
  XNOR U4843 ( .A(n4403), .B(n4404), .Z(n4369) );
  XNOR U4844 ( .A(n4390), .B(n4405), .Z(n4404) );
  XNOR U4845 ( .A(n4323), .B(n4384), .Z(n4405) );
  XOR U4846 ( .A(n4391), .B(n4406), .Z(n4384) );
  XNOR U4847 ( .A(n4407), .B(n4408), .Z(n4406) );
  NAND U4848 ( .A(n4350), .B(n4320), .Z(n4408) );
  XNOR U4849 ( .A(n4409), .B(n4407), .Z(n4391) );
  NANDN U4850 ( .A(n4352), .B(n4329), .Z(n4407) );
  XOR U4851 ( .A(n4330), .B(n4320), .Z(n4329) );
  XNOR U4852 ( .A(n4410), .B(n4293), .Z(n4320) );
  XOR U4853 ( .A(n4361), .B(n4350), .Z(n4352) );
  XOR U4854 ( .A(n4341), .B(n4411), .Z(n4350) );
  ANDN U4855 ( .B(n4330), .A(n4361), .Z(n4409) );
  XOR U4856 ( .A(n4399), .B(n4346), .Z(n4361) );
  XOR U4857 ( .A(n4412), .B(n4413), .Z(n4346) );
  XNOR U4858 ( .A(n4414), .B(n4415), .Z(n4413) );
  XOR U4859 ( .A(n4416), .B(n4398), .Z(n4330) );
  XOR U4860 ( .A(n4411), .B(n4394), .Z(n4390) );
  IV U4861 ( .A(n4293), .Z(n4394) );
  XOR U4862 ( .A(n4417), .B(n4418), .Z(n4293) );
  XNOR U4863 ( .A(n4419), .B(n4415), .Z(n4418) );
  IV U4864 ( .A(n4336), .Z(n4411) );
  XOR U4865 ( .A(n4415), .B(n4420), .Z(n4336) );
  XNOR U4866 ( .A(n4341), .B(n4421), .Z(n4403) );
  XNOR U4867 ( .A(n4422), .B(n4402), .Z(n4421) );
  OR U4868 ( .A(n4326), .B(n4340), .Z(n4402) );
  XNOR U4869 ( .A(n4399), .B(n4341), .Z(n4340) );
  XOR U4870 ( .A(n4315), .B(n4410), .Z(n4326) );
  IV U4871 ( .A(n4323), .Z(n4410) );
  XOR U4872 ( .A(n4398), .B(n4423), .Z(n4323) );
  XNOR U4873 ( .A(n4419), .B(n4412), .Z(n4423) );
  XOR U4874 ( .A(n4424), .B(n4425), .Z(n4412) );
  XOR U4875 ( .A(n1071), .B(n389), .Z(n4425) );
  XNOR U4876 ( .A(n431), .B(n4426), .Z(n4424) );
  XNOR U4877 ( .A(key[1194]), .B(n1076), .Z(n4426) );
  IV U4878 ( .A(n4305), .Z(n4398) );
  XOR U4879 ( .A(n4417), .B(n4427), .Z(n4305) );
  XOR U4880 ( .A(n4415), .B(n4428), .Z(n4427) );
  ANDN U4881 ( .B(n4416), .A(n4286), .Z(n4422) );
  IV U4882 ( .A(n4315), .Z(n4416) );
  XOR U4883 ( .A(n4417), .B(n4429), .Z(n4315) );
  XOR U4884 ( .A(n4415), .B(n4430), .Z(n4429) );
  XOR U4885 ( .A(n4431), .B(n4432), .Z(n4415) );
  XOR U4886 ( .A(n4433), .B(n4286), .Z(n4432) );
  IV U4887 ( .A(n4399), .Z(n4286) );
  XOR U4888 ( .A(n4434), .B(n4435), .Z(n4431) );
  XNOR U4889 ( .A(key[1198]), .B(n400), .Z(n4435) );
  XNOR U4890 ( .A(n4436), .B(n411), .Z(n400) );
  XNOR U4891 ( .A(n4437), .B(n4438), .Z(n411) );
  IV U4892 ( .A(n4420), .Z(n4417) );
  XOR U4893 ( .A(n4439), .B(n4440), .Z(n4420) );
  XOR U4894 ( .A(n1063), .B(n404), .Z(n4440) );
  XNOR U4895 ( .A(n4441), .B(n1048), .Z(n404) );
  XNOR U4896 ( .A(n398), .B(n4442), .Z(n4439) );
  XNOR U4897 ( .A(key[1197]), .B(n1042), .Z(n4442) );
  XOR U4898 ( .A(n4443), .B(n4444), .Z(n4341) );
  XNOR U4899 ( .A(n4430), .B(n4428), .Z(n4444) );
  XNOR U4900 ( .A(n4445), .B(n4446), .Z(n4428) );
  XOR U4901 ( .A(n1043), .B(n412), .Z(n4446) );
  XOR U4902 ( .A(key[1199]), .B(n437), .Z(n4445) );
  IV U4903 ( .A(n1081), .Z(n437) );
  XOR U4904 ( .A(n4448), .B(n4437), .Z(n1081) );
  XNOR U4905 ( .A(n4449), .B(n4450), .Z(n4430) );
  XNOR U4906 ( .A(n416), .B(n4451), .Z(n4450) );
  XNOR U4907 ( .A(n4452), .B(n1061), .Z(n416) );
  XNOR U4908 ( .A(n418), .B(n4453), .Z(n4449) );
  XOR U4909 ( .A(key[1196]), .B(n1077), .Z(n4453) );
  XNOR U4910 ( .A(n4437), .B(n406), .Z(n418) );
  XOR U4911 ( .A(n4399), .B(n4414), .Z(n4443) );
  XOR U4912 ( .A(n4454), .B(n4455), .Z(n4414) );
  XNOR U4913 ( .A(n4419), .B(n4456), .Z(n4455) );
  XNOR U4914 ( .A(n1031), .B(n4457), .Z(n4456) );
  XOR U4915 ( .A(n4458), .B(n4459), .Z(n4419) );
  XNOR U4916 ( .A(n391), .B(n1030), .Z(n4459) );
  XNOR U4917 ( .A(n428), .B(n4460), .Z(n4458) );
  XOR U4918 ( .A(key[1193]), .B(n4461), .Z(n4460) );
  XNOR U4919 ( .A(n425), .B(n4462), .Z(n4454) );
  XOR U4920 ( .A(key[1195]), .B(n4463), .Z(n4462) );
  XOR U4921 ( .A(n4437), .B(n420), .Z(n425) );
  XOR U4922 ( .A(n4464), .B(n4465), .Z(n4399) );
  XOR U4923 ( .A(n1073), .B(n1055), .Z(n4465) );
  XOR U4924 ( .A(n4448), .B(n4466), .Z(n4464) );
  XOR U4925 ( .A(key[1192]), .B(n430), .Z(n4466) );
  XOR U4926 ( .A(n4467), .B(n4468), .Z(out[103]) );
  XNOR U4927 ( .A(n16), .B(n4469), .Z(n4468) );
  IV U4928 ( .A(n4470), .Z(n16) );
  XNOR U4929 ( .A(n8), .B(n4471), .Z(n4467) );
  XOR U4930 ( .A(key[1255]), .B(n4472), .Z(n4471) );
  XNOR U4931 ( .A(n4473), .B(n4474), .Z(n8) );
  XNOR U4932 ( .A(n4475), .B(n4476), .Z(n4474) );
  NANDN U4933 ( .A(n4477), .B(n4478), .Z(n4476) );
  XOR U4934 ( .A(n4470), .B(n4479), .Z(out[102]) );
  XNOR U4935 ( .A(key[1254]), .B(n10), .Z(n4479) );
  XNOR U4936 ( .A(n4481), .B(n4482), .Z(n4480) );
  OR U4937 ( .A(n4483), .B(n4484), .Z(n4482) );
  XNOR U4938 ( .A(n4485), .B(n4486), .Z(n4473) );
  XNOR U4939 ( .A(n4487), .B(n4488), .Z(n4486) );
  NAND U4940 ( .A(n4489), .B(n4490), .Z(n4488) );
  XNOR U4941 ( .A(n9), .B(n19), .Z(n4470) );
  XNOR U4942 ( .A(n4485), .B(n4491), .Z(n9) );
  XNOR U4943 ( .A(n4475), .B(n4492), .Z(n4491) );
  NANDN U4944 ( .A(n4493), .B(n4494), .Z(n4492) );
  OR U4945 ( .A(n4495), .B(n4496), .Z(n4475) );
  XOR U4946 ( .A(n4497), .B(n4498), .Z(out[101]) );
  XNOR U4947 ( .A(n4469), .B(n4499), .Z(n4498) );
  XOR U4948 ( .A(n4485), .B(n17), .Z(n4499) );
  XOR U4949 ( .A(n4500), .B(n4487), .Z(n4485) );
  NANDN U4950 ( .A(n4501), .B(n4502), .Z(n4487) );
  ANDN U4951 ( .B(n4503), .A(n4504), .Z(n4500) );
  XNOR U4952 ( .A(n4505), .B(n4506), .Z(n4469) );
  XNOR U4953 ( .A(n4507), .B(n4508), .Z(n4506) );
  NANDN U4954 ( .A(n4509), .B(n4478), .Z(n4508) );
  XOR U4955 ( .A(n4510), .B(n4511), .Z(n4497) );
  XNOR U4956 ( .A(key[1253]), .B(n4481), .Z(n4511) );
  NANDN U4957 ( .A(n4512), .B(n4513), .Z(n4481) );
  ANDN U4958 ( .B(n4514), .A(n4515), .Z(n4510) );
  XOR U4959 ( .A(n17), .B(n4516), .Z(out[100]) );
  XNOR U4960 ( .A(key[1252]), .B(n13), .Z(n4516) );
  XOR U4961 ( .A(n4472), .B(n19), .Z(n13) );
  XOR U4962 ( .A(n4517), .B(n4518), .Z(n19) );
  XOR U4963 ( .A(n4519), .B(n4507), .Z(n4518) );
  OR U4964 ( .A(n4495), .B(n4520), .Z(n4507) );
  XNOR U4965 ( .A(n4478), .B(n4494), .Z(n4495) );
  ANDN U4966 ( .B(n4494), .A(n4521), .Z(n4519) );
  IV U4967 ( .A(n12), .Z(n4472) );
  XNOR U4968 ( .A(n4517), .B(n4522), .Z(n12) );
  XNOR U4969 ( .A(n4523), .B(n4524), .Z(n4522) );
  NAND U4970 ( .A(n4514), .B(n4525), .Z(n4524) );
  XOR U4971 ( .A(n4505), .B(n4526), .Z(n17) );
  XOR U4972 ( .A(n4527), .B(n4523), .Z(n4526) );
  NANDN U4973 ( .A(n4528), .B(n4513), .Z(n4523) );
  XNOR U4974 ( .A(n4483), .B(n4514), .Z(n4513) );
  NOR U4975 ( .A(n4529), .B(n4483), .Z(n4527) );
  XNOR U4976 ( .A(n4517), .B(n4530), .Z(n4505) );
  XNOR U4977 ( .A(n4531), .B(n4532), .Z(n4530) );
  NAND U4978 ( .A(n4490), .B(n4533), .Z(n4532) );
  XOR U4979 ( .A(n4534), .B(n4531), .Z(n4517) );
  OR U4980 ( .A(n4501), .B(n4535), .Z(n4531) );
  XOR U4981 ( .A(n4504), .B(n4490), .Z(n4501) );
  XOR U4982 ( .A(n4494), .B(n4514), .Z(n4490) );
  XOR U4983 ( .A(n4536), .B(n4537), .Z(n4514) );
  NANDN U4984 ( .A(n4538), .B(n4539), .Z(n4537) );
  XOR U4985 ( .A(n4540), .B(n4541), .Z(n4494) );
  NANDN U4986 ( .A(n4538), .B(n4542), .Z(n4541) );
  NOR U4987 ( .A(n4504), .B(n4543), .Z(n4534) );
  XOR U4988 ( .A(n4483), .B(n4478), .Z(n4504) );
  XNOR U4989 ( .A(n4544), .B(n4540), .Z(n4478) );
  NANDN U4990 ( .A(n4545), .B(n4546), .Z(n4540) );
  XOR U4991 ( .A(n4542), .B(n4547), .Z(n4546) );
  ANDN U4992 ( .B(n4547), .A(n4548), .Z(n4544) );
  XOR U4993 ( .A(n4549), .B(n4536), .Z(n4483) );
  NANDN U4994 ( .A(n4545), .B(n4550), .Z(n4536) );
  XOR U4995 ( .A(n4551), .B(n4539), .Z(n4550) );
  XNOR U4996 ( .A(n4552), .B(n4553), .Z(n4538) );
  XOR U4997 ( .A(n4554), .B(n4555), .Z(n4553) );
  XNOR U4998 ( .A(n4556), .B(n4557), .Z(n4552) );
  XNOR U4999 ( .A(n4558), .B(n4559), .Z(n4557) );
  ANDN U5000 ( .B(n4551), .A(n4555), .Z(n4558) );
  ANDN U5001 ( .B(n4551), .A(n4548), .Z(n4549) );
  XNOR U5002 ( .A(n4554), .B(n4560), .Z(n4548) );
  XOR U5003 ( .A(n4561), .B(n4559), .Z(n4560) );
  NAND U5004 ( .A(n4562), .B(n4563), .Z(n4559) );
  XNOR U5005 ( .A(n4556), .B(n4539), .Z(n4563) );
  IV U5006 ( .A(n4551), .Z(n4556) );
  XNOR U5007 ( .A(n4542), .B(n4555), .Z(n4562) );
  IV U5008 ( .A(n4547), .Z(n4555) );
  XOR U5009 ( .A(n4564), .B(n4565), .Z(n4547) );
  XNOR U5010 ( .A(n4566), .B(n4567), .Z(n4565) );
  XNOR U5011 ( .A(n4568), .B(n4569), .Z(n4564) );
  ANDN U5012 ( .B(n4570), .A(n4529), .Z(n4568) );
  AND U5013 ( .A(n4539), .B(n4542), .Z(n4561) );
  XNOR U5014 ( .A(n4539), .B(n4542), .Z(n4554) );
  XNOR U5015 ( .A(n4571), .B(n4572), .Z(n4542) );
  XOR U5016 ( .A(n4573), .B(n4567), .Z(n4572) );
  XNOR U5017 ( .A(n4574), .B(n4575), .Z(n4571) );
  XNOR U5018 ( .A(n4576), .B(n4569), .Z(n4575) );
  OR U5019 ( .A(n4512), .B(n4528), .Z(n4569) );
  XNOR U5020 ( .A(n4577), .B(n4525), .Z(n4528) );
  XNOR U5021 ( .A(n4515), .B(n4484), .Z(n4512) );
  ANDN U5022 ( .B(n4525), .A(n4515), .Z(n4576) );
  XNOR U5023 ( .A(n4578), .B(n4579), .Z(n4539) );
  XNOR U5024 ( .A(n4567), .B(n4580), .Z(n4579) );
  XOR U5025 ( .A(n4477), .B(n4573), .Z(n4580) );
  XNOR U5026 ( .A(n4577), .B(n4484), .Z(n4567) );
  XOR U5027 ( .A(n4509), .B(n4581), .Z(n4578) );
  XNOR U5028 ( .A(n4582), .B(n4583), .Z(n4581) );
  XNOR U5029 ( .A(n4584), .B(n4585), .Z(n4551) );
  XNOR U5030 ( .A(n4566), .B(n4586), .Z(n4585) );
  XNOR U5031 ( .A(n4574), .B(n4493), .Z(n4586) );
  XOR U5032 ( .A(n4525), .B(n4587), .Z(n4574) );
  XOR U5033 ( .A(n4573), .B(n4588), .Z(n4566) );
  XNOR U5034 ( .A(n4589), .B(n4590), .Z(n4588) );
  NAND U5035 ( .A(n4533), .B(n4489), .Z(n4590) );
  XNOR U5036 ( .A(n4591), .B(n4589), .Z(n4573) );
  NANDN U5037 ( .A(n4535), .B(n4502), .Z(n4589) );
  XOR U5038 ( .A(n4503), .B(n4489), .Z(n4502) );
  XNOR U5039 ( .A(n4587), .B(n4493), .Z(n4489) );
  IV U5040 ( .A(n4515), .Z(n4587) );
  XOR U5041 ( .A(n4592), .B(n4593), .Z(n4515) );
  XOR U5042 ( .A(n4594), .B(n4595), .Z(n4593) );
  XOR U5043 ( .A(n4543), .B(n4533), .Z(n4535) );
  XOR U5044 ( .A(n4525), .B(n4596), .Z(n4533) );
  ANDN U5045 ( .B(n4503), .A(n4543), .Z(n4591) );
  XOR U5046 ( .A(n4509), .B(n4577), .Z(n4543) );
  IV U5047 ( .A(n4529), .Z(n4577) );
  XOR U5048 ( .A(n4597), .B(n4598), .Z(n4529) );
  XOR U5049 ( .A(n4599), .B(n4594), .Z(n4598) );
  XOR U5050 ( .A(n4600), .B(n4570), .Z(n4503) );
  XNOR U5051 ( .A(n4596), .B(n4601), .Z(n4584) );
  XNOR U5052 ( .A(n4602), .B(n4583), .Z(n4601) );
  OR U5053 ( .A(n4496), .B(n4520), .Z(n4583) );
  XNOR U5054 ( .A(n4509), .B(n4521), .Z(n4520) );
  IV U5055 ( .A(n4596), .Z(n4521) );
  XNOR U5056 ( .A(n4477), .B(n4493), .Z(n4496) );
  XOR U5057 ( .A(n4570), .B(n4603), .Z(n4493) );
  XNOR U5058 ( .A(n4599), .B(n4595), .Z(n4603) );
  XOR U5059 ( .A(n4604), .B(n4605), .Z(n4599) );
  XOR U5060 ( .A(n645), .B(n1283), .Z(n4605) );
  IV U5061 ( .A(n1871), .Z(n1283) );
  XNOR U5062 ( .A(n640), .B(n650), .Z(n1871) );
  XOR U5063 ( .A(n1873), .B(n652), .Z(n645) );
  XOR U5064 ( .A(n4606), .B(n4607), .Z(n652) );
  XOR U5065 ( .A(n4608), .B(n4609), .Z(n4607) );
  XNOR U5066 ( .A(n4610), .B(n4611), .Z(n4606) );
  XNOR U5067 ( .A(key[1154]), .B(n1907), .Z(n4604) );
  IV U5068 ( .A(n4484), .Z(n4570) );
  XNOR U5069 ( .A(n4612), .B(n4525), .Z(n4484) );
  NOR U5070 ( .A(n4477), .B(n4509), .Z(n4602) );
  IV U5071 ( .A(n4600), .Z(n4477) );
  XOR U5072 ( .A(n4613), .B(n4525), .Z(n4600) );
  XNOR U5073 ( .A(n4594), .B(n4592), .Z(n4525) );
  XNOR U5074 ( .A(n4614), .B(n4615), .Z(n4592) );
  XOR U5075 ( .A(n1257), .B(n1252), .Z(n4615) );
  XNOR U5076 ( .A(n1888), .B(n612), .Z(n1252) );
  XOR U5077 ( .A(n4616), .B(n4609), .Z(n612) );
  XOR U5078 ( .A(n4617), .B(n4618), .Z(n4609) );
  XOR U5079 ( .A(n4619), .B(n4620), .Z(n4618) );
  NOR U5080 ( .A(n4621), .B(n4622), .Z(n4619) );
  XNOR U5081 ( .A(key[1157]), .B(n1886), .Z(n4614) );
  XNOR U5082 ( .A(n1256), .B(n1898), .Z(n1886) );
  IV U5083 ( .A(n614), .Z(n1898) );
  XOR U5084 ( .A(n4623), .B(n4624), .Z(n614) );
  XNOR U5085 ( .A(n4625), .B(n4626), .Z(n4624) );
  XNOR U5086 ( .A(n4627), .B(n4628), .Z(n4623) );
  XOR U5087 ( .A(n4629), .B(n4630), .Z(n4628) );
  ANDN U5088 ( .B(n4631), .A(n4632), .Z(n4630) );
  XNOR U5089 ( .A(n4633), .B(n4634), .Z(n1256) );
  XNOR U5090 ( .A(n4635), .B(n4636), .Z(n4634) );
  XNOR U5091 ( .A(n4637), .B(n4638), .Z(n4633) );
  XOR U5092 ( .A(n4639), .B(n4640), .Z(n4638) );
  ANDN U5093 ( .B(n4641), .A(n4642), .Z(n4640) );
  XNOR U5094 ( .A(n4643), .B(n4644), .Z(n4594) );
  XNOR U5095 ( .A(n1883), .B(n628), .Z(n4644) );
  XNOR U5096 ( .A(n4645), .B(n1265), .Z(n628) );
  XNOR U5097 ( .A(n4646), .B(n4647), .Z(n1265) );
  XNOR U5098 ( .A(n4616), .B(n4648), .Z(n4647) );
  XOR U5099 ( .A(n4610), .B(n4649), .Z(n4646) );
  XNOR U5100 ( .A(n4650), .B(n1259), .Z(n1883) );
  XNOR U5101 ( .A(n630), .B(n616), .Z(n1259) );
  XOR U5102 ( .A(n4651), .B(n4652), .Z(n616) );
  XOR U5103 ( .A(n4653), .B(n4654), .Z(n630) );
  XOR U5104 ( .A(n1888), .B(n4655), .Z(n4643) );
  XOR U5105 ( .A(key[1158]), .B(n4509), .Z(n4655) );
  XNOR U5106 ( .A(n4656), .B(n4657), .Z(n1888) );
  XOR U5107 ( .A(n4658), .B(n4659), .Z(n4596) );
  XNOR U5108 ( .A(n4613), .B(n4612), .Z(n4659) );
  XOR U5109 ( .A(n4660), .B(n4661), .Z(n4612) );
  XNOR U5110 ( .A(n623), .B(n1893), .Z(n4661) );
  XNOR U5111 ( .A(n1881), .B(n1267), .Z(n1893) );
  XNOR U5112 ( .A(n4662), .B(n4663), .Z(n1267) );
  XNOR U5113 ( .A(n4664), .B(n4636), .Z(n4663) );
  XNOR U5114 ( .A(n4665), .B(n4666), .Z(n4636) );
  XNOR U5115 ( .A(n4667), .B(n4668), .Z(n4666) );
  OR U5116 ( .A(n4669), .B(n4670), .Z(n4668) );
  XOR U5117 ( .A(n4671), .B(n4651), .Z(n4662) );
  IV U5118 ( .A(n609), .Z(n1881) );
  XOR U5119 ( .A(n4672), .B(n4673), .Z(n609) );
  XOR U5120 ( .A(n4674), .B(n4626), .Z(n4673) );
  XNOR U5121 ( .A(n4675), .B(n4676), .Z(n4626) );
  XNOR U5122 ( .A(n4677), .B(n4678), .Z(n4676) );
  OR U5123 ( .A(n4679), .B(n4680), .Z(n4678) );
  XNOR U5124 ( .A(n4681), .B(n4653), .Z(n4672) );
  XNOR U5125 ( .A(key[1159]), .B(n4650), .Z(n4660) );
  XNOR U5126 ( .A(n1288), .B(n1264), .Z(n4650) );
  XOR U5127 ( .A(n4682), .B(n4683), .Z(n1264) );
  XOR U5128 ( .A(n4684), .B(n4685), .Z(n4683) );
  XNOR U5129 ( .A(n4656), .B(n4686), .Z(n4682) );
  XOR U5130 ( .A(n4687), .B(n4688), .Z(n4613) );
  XOR U5131 ( .A(n599), .B(n1897), .Z(n4688) );
  XOR U5132 ( .A(n1276), .B(n597), .Z(n1897) );
  XOR U5133 ( .A(n4627), .B(n650), .Z(n597) );
  XNOR U5134 ( .A(n4689), .B(n4690), .Z(n650) );
  XNOR U5135 ( .A(n4637), .B(n640), .Z(n1276) );
  XOR U5136 ( .A(n4691), .B(n4671), .Z(n640) );
  XOR U5137 ( .A(n623), .B(n1258), .Z(n599) );
  XNOR U5138 ( .A(n4692), .B(n4693), .Z(n1258) );
  XNOR U5139 ( .A(n4694), .B(n4648), .Z(n4693) );
  XNOR U5140 ( .A(n4695), .B(n4696), .Z(n4648) );
  XNOR U5141 ( .A(n4697), .B(n4698), .Z(n4696) );
  NANDN U5142 ( .A(n4699), .B(n4700), .Z(n4698) );
  XNOR U5143 ( .A(n4701), .B(n4702), .Z(n4692) );
  XNOR U5144 ( .A(n4620), .B(n4703), .Z(n4702) );
  ANDN U5145 ( .B(n4704), .A(n4705), .Z(n4703) );
  OR U5146 ( .A(n4706), .B(n4707), .Z(n4620) );
  XNOR U5147 ( .A(n1899), .B(n4708), .Z(n4687) );
  XNOR U5148 ( .A(key[1156]), .B(n1274), .Z(n4708) );
  XNOR U5149 ( .A(n1288), .B(n1257), .Z(n1899) );
  XOR U5150 ( .A(n4709), .B(n4710), .Z(n1257) );
  XNOR U5151 ( .A(n4711), .B(n4685), .Z(n4710) );
  XNOR U5152 ( .A(n4712), .B(n4713), .Z(n4685) );
  XOR U5153 ( .A(n4714), .B(n4715), .Z(n4713) );
  NANDN U5154 ( .A(n4716), .B(n4717), .Z(n4715) );
  XNOR U5155 ( .A(n4718), .B(n4719), .Z(n4709) );
  XNOR U5156 ( .A(n4720), .B(n4721), .Z(n4719) );
  ANDN U5157 ( .B(n4722), .A(n4723), .Z(n4721) );
  XNOR U5158 ( .A(n4509), .B(n4597), .Z(n4658) );
  XOR U5159 ( .A(n4724), .B(n4725), .Z(n4597) );
  XNOR U5160 ( .A(n1904), .B(n4726), .Z(n4725) );
  XOR U5161 ( .A(n4595), .B(n1243), .Z(n4726) );
  XOR U5162 ( .A(n1870), .B(n649), .Z(n1243) );
  XNOR U5163 ( .A(n4727), .B(n4728), .Z(n649) );
  XNOR U5164 ( .A(n4729), .B(n4730), .Z(n4652) );
  XNOR U5165 ( .A(n4731), .B(n4639), .Z(n4730) );
  ANDN U5166 ( .B(n4732), .A(n4733), .Z(n4639) );
  ANDN U5167 ( .B(n4734), .A(n4735), .Z(n4731) );
  XNOR U5168 ( .A(n4671), .B(n4736), .Z(n4727) );
  IV U5169 ( .A(n635), .Z(n1870) );
  XOR U5170 ( .A(n4737), .B(n4738), .Z(n635) );
  XOR U5171 ( .A(n4654), .B(n4674), .Z(n4738) );
  XNOR U5172 ( .A(n4739), .B(n4740), .Z(n4654) );
  XNOR U5173 ( .A(n4741), .B(n4629), .Z(n4740) );
  ANDN U5174 ( .B(n4742), .A(n4743), .Z(n4629) );
  ANDN U5175 ( .B(n4744), .A(n4745), .Z(n4741) );
  XOR U5176 ( .A(n4681), .B(n4746), .Z(n4737) );
  XOR U5177 ( .A(n4747), .B(n4748), .Z(n4595) );
  XNOR U5178 ( .A(n648), .B(n1287), .Z(n4748) );
  XOR U5179 ( .A(n624), .B(n639), .Z(n1287) );
  XNOR U5180 ( .A(n4674), .B(n4749), .Z(n639) );
  XOR U5181 ( .A(n4681), .B(n4653), .Z(n4749) );
  XOR U5182 ( .A(n4689), .B(n4746), .Z(n4653) );
  XNOR U5183 ( .A(n4625), .B(n4750), .Z(n4746) );
  XNOR U5184 ( .A(n4751), .B(n4752), .Z(n4750) );
  NANDN U5185 ( .A(n4753), .B(n4754), .Z(n4752) );
  IV U5186 ( .A(n4690), .Z(n4681) );
  XOR U5187 ( .A(n4755), .B(n4756), .Z(n4690) );
  XOR U5188 ( .A(n4757), .B(n4758), .Z(n4756) );
  NAND U5189 ( .A(n4759), .B(n4631), .Z(n4758) );
  XOR U5190 ( .A(n4739), .B(n4760), .Z(n4674) );
  XNOR U5191 ( .A(n4751), .B(n4761), .Z(n4760) );
  OR U5192 ( .A(n4679), .B(n4762), .Z(n4761) );
  OR U5193 ( .A(n4763), .B(n4764), .Z(n4751) );
  XNOR U5194 ( .A(n4625), .B(n4765), .Z(n4739) );
  XNOR U5195 ( .A(n4766), .B(n4767), .Z(n4765) );
  NANDN U5196 ( .A(n4768), .B(n4769), .Z(n4767) );
  XOR U5197 ( .A(n4770), .B(n4766), .Z(n4625) );
  NANDN U5198 ( .A(n4771), .B(n4772), .Z(n4766) );
  ANDN U5199 ( .B(n4773), .A(n4774), .Z(n4770) );
  XNOR U5200 ( .A(n4664), .B(n4775), .Z(n624) );
  XNOR U5201 ( .A(n4671), .B(n4651), .Z(n4775) );
  XOR U5202 ( .A(n4691), .B(n4736), .Z(n4651) );
  XNOR U5203 ( .A(n4635), .B(n4776), .Z(n4736) );
  XNOR U5204 ( .A(n4777), .B(n4778), .Z(n4776) );
  NANDN U5205 ( .A(n4779), .B(n4780), .Z(n4778) );
  XOR U5206 ( .A(n4781), .B(n4782), .Z(n4671) );
  XOR U5207 ( .A(n4783), .B(n4784), .Z(n4782) );
  NAND U5208 ( .A(n4785), .B(n4641), .Z(n4784) );
  XNOR U5209 ( .A(n4729), .B(n4786), .Z(n4664) );
  XNOR U5210 ( .A(n4777), .B(n4787), .Z(n4786) );
  OR U5211 ( .A(n4669), .B(n4788), .Z(n4787) );
  OR U5212 ( .A(n4789), .B(n4790), .Z(n4777) );
  XNOR U5213 ( .A(n4635), .B(n4791), .Z(n4729) );
  XNOR U5214 ( .A(n4792), .B(n4793), .Z(n4791) );
  NANDN U5215 ( .A(n4794), .B(n4795), .Z(n4793) );
  XOR U5216 ( .A(n4796), .B(n4792), .Z(n4635) );
  NANDN U5217 ( .A(n4797), .B(n4798), .Z(n4792) );
  ANDN U5218 ( .B(n4799), .A(n4800), .Z(n4796) );
  IV U5219 ( .A(n1242), .Z(n648) );
  XNOR U5220 ( .A(n1907), .B(n638), .Z(n1242) );
  XNOR U5221 ( .A(key[1153]), .B(n4801), .Z(n4747) );
  XNOR U5222 ( .A(n1288), .B(n1274), .Z(n1904) );
  XNOR U5223 ( .A(n4711), .B(n1907), .Z(n1274) );
  XOR U5224 ( .A(n4802), .B(n4803), .Z(n1907) );
  XNOR U5225 ( .A(n643), .B(n4804), .Z(n4724) );
  XNOR U5226 ( .A(key[1155]), .B(n1873), .Z(n4804) );
  XOR U5227 ( .A(n4805), .B(n4806), .Z(n1873) );
  XNOR U5228 ( .A(n4807), .B(n4657), .Z(n4806) );
  XNOR U5229 ( .A(n4808), .B(n4809), .Z(n4657) );
  XOR U5230 ( .A(n4810), .B(n4720), .Z(n4809) );
  OR U5231 ( .A(n4811), .B(n4812), .Z(n4720) );
  NOR U5232 ( .A(n4813), .B(n4814), .Z(n4810) );
  XOR U5233 ( .A(n4815), .B(n4686), .Z(n4805) );
  XOR U5234 ( .A(n4645), .B(n1275), .Z(n643) );
  XOR U5235 ( .A(n4694), .B(n638), .Z(n1275) );
  XOR U5236 ( .A(n4611), .B(n4816), .Z(n638) );
  IV U5237 ( .A(n623), .Z(n4645) );
  XOR U5238 ( .A(n4816), .B(n4694), .Z(n623) );
  XNOR U5239 ( .A(n4695), .B(n4817), .Z(n4694) );
  XOR U5240 ( .A(n4818), .B(n4819), .Z(n4817) );
  ANDN U5241 ( .B(n4820), .A(n4622), .Z(n4818) );
  XNOR U5242 ( .A(n4821), .B(n4822), .Z(n4695) );
  XNOR U5243 ( .A(n4823), .B(n4824), .Z(n4822) );
  NAND U5244 ( .A(n4825), .B(n4826), .Z(n4824) );
  XNOR U5245 ( .A(n4827), .B(n4828), .Z(n4509) );
  XOR U5246 ( .A(n642), .B(n1894), .Z(n4828) );
  IV U5247 ( .A(n625), .Z(n1894) );
  XOR U5248 ( .A(n1880), .B(n1288), .Z(n625) );
  XNOR U5249 ( .A(n4712), .B(n4829), .Z(n4711) );
  XOR U5250 ( .A(n4830), .B(n4831), .Z(n4829) );
  NOR U5251 ( .A(n4832), .B(n4814), .Z(n4830) );
  XNOR U5252 ( .A(n4833), .B(n4834), .Z(n4712) );
  XNOR U5253 ( .A(n4835), .B(n4836), .Z(n4834) );
  NANDN U5254 ( .A(n4837), .B(n4838), .Z(n4836) );
  XOR U5255 ( .A(n4689), .B(n4627), .Z(n1880) );
  XNOR U5256 ( .A(n4675), .B(n4839), .Z(n4627) );
  XNOR U5257 ( .A(n4840), .B(n4757), .Z(n4839) );
  XOR U5258 ( .A(n4744), .B(n4631), .Z(n4742) );
  ANDN U5259 ( .B(n4744), .A(n4842), .Z(n4840) );
  XNOR U5260 ( .A(n4755), .B(n4843), .Z(n4675) );
  XNOR U5261 ( .A(n4844), .B(n4845), .Z(n4843) );
  NANDN U5262 ( .A(n4768), .B(n4846), .Z(n4845) );
  XNOR U5263 ( .A(n4755), .B(n4847), .Z(n4689) );
  XOR U5264 ( .A(n4848), .B(n4677), .Z(n4847) );
  OR U5265 ( .A(n4849), .B(n4763), .Z(n4677) );
  XNOR U5266 ( .A(n4679), .B(n4753), .Z(n4763) );
  NOR U5267 ( .A(n4850), .B(n4753), .Z(n4848) );
  XOR U5268 ( .A(n4851), .B(n4844), .Z(n4755) );
  OR U5269 ( .A(n4771), .B(n4852), .Z(n4844) );
  XOR U5270 ( .A(n4853), .B(n4768), .Z(n4771) );
  XOR U5271 ( .A(n4753), .B(n4631), .Z(n4768) );
  XOR U5272 ( .A(n4854), .B(n4855), .Z(n4631) );
  NANDN U5273 ( .A(n4856), .B(n4857), .Z(n4855) );
  XNOR U5274 ( .A(n4858), .B(n4859), .Z(n4753) );
  OR U5275 ( .A(n4856), .B(n4860), .Z(n4859) );
  ANDN U5276 ( .B(n4853), .A(n4861), .Z(n4851) );
  IV U5277 ( .A(n4774), .Z(n4853) );
  XOR U5278 ( .A(n4679), .B(n4744), .Z(n4774) );
  XNOR U5279 ( .A(n4862), .B(n4854), .Z(n4744) );
  NANDN U5280 ( .A(n4863), .B(n4864), .Z(n4854) );
  ANDN U5281 ( .B(n4865), .A(n4866), .Z(n4862) );
  NANDN U5282 ( .A(n4863), .B(n4868), .Z(n4858) );
  XOR U5283 ( .A(n4869), .B(n4856), .Z(n4863) );
  XNOR U5284 ( .A(n4870), .B(n4871), .Z(n4856) );
  XOR U5285 ( .A(n4872), .B(n4865), .Z(n4871) );
  XNOR U5286 ( .A(n4873), .B(n4874), .Z(n4870) );
  XNOR U5287 ( .A(n4875), .B(n4876), .Z(n4874) );
  ANDN U5288 ( .B(n4865), .A(n4877), .Z(n4875) );
  IV U5289 ( .A(n4878), .Z(n4865) );
  ANDN U5290 ( .B(n4869), .A(n4877), .Z(n4867) );
  IV U5291 ( .A(n4873), .Z(n4877) );
  IV U5292 ( .A(n4866), .Z(n4869) );
  XNOR U5293 ( .A(n4872), .B(n4879), .Z(n4866) );
  XOR U5294 ( .A(n4880), .B(n4876), .Z(n4879) );
  NAND U5295 ( .A(n4868), .B(n4864), .Z(n4876) );
  XNOR U5296 ( .A(n4857), .B(n4878), .Z(n4864) );
  XOR U5297 ( .A(n4881), .B(n4882), .Z(n4878) );
  XOR U5298 ( .A(n4883), .B(n4884), .Z(n4882) );
  XNOR U5299 ( .A(n4754), .B(n4885), .Z(n4884) );
  XNOR U5300 ( .A(n4886), .B(n4887), .Z(n4881) );
  XNOR U5301 ( .A(n4888), .B(n4889), .Z(n4887) );
  ANDN U5302 ( .B(n4890), .A(n4680), .Z(n4888) );
  XNOR U5303 ( .A(n4873), .B(n4860), .Z(n4868) );
  XOR U5304 ( .A(n4891), .B(n4892), .Z(n4873) );
  XNOR U5305 ( .A(n4893), .B(n4885), .Z(n4892) );
  XOR U5306 ( .A(n4894), .B(n4895), .Z(n4885) );
  XNOR U5307 ( .A(n4896), .B(n4897), .Z(n4895) );
  NAND U5308 ( .A(n4846), .B(n4769), .Z(n4897) );
  XNOR U5309 ( .A(n4898), .B(n4899), .Z(n4891) );
  ANDN U5310 ( .B(n4900), .A(n4842), .Z(n4898) );
  ANDN U5311 ( .B(n4857), .A(n4860), .Z(n4880) );
  XOR U5312 ( .A(n4860), .B(n4857), .Z(n4872) );
  XNOR U5313 ( .A(n4901), .B(n4902), .Z(n4857) );
  XNOR U5314 ( .A(n4894), .B(n4903), .Z(n4902) );
  XOR U5315 ( .A(n4893), .B(n4762), .Z(n4903) );
  XOR U5316 ( .A(n4680), .B(n4904), .Z(n4901) );
  XNOR U5317 ( .A(n4905), .B(n4889), .Z(n4904) );
  OR U5318 ( .A(n4764), .B(n4849), .Z(n4889) );
  XNOR U5319 ( .A(n4680), .B(n4850), .Z(n4849) );
  XOR U5320 ( .A(n4762), .B(n4754), .Z(n4764) );
  ANDN U5321 ( .B(n4754), .A(n4850), .Z(n4905) );
  XOR U5322 ( .A(n4906), .B(n4907), .Z(n4860) );
  XOR U5323 ( .A(n4894), .B(n4883), .Z(n4907) );
  XOR U5324 ( .A(n4759), .B(n4632), .Z(n4883) );
  XOR U5325 ( .A(n4908), .B(n4896), .Z(n4894) );
  NANDN U5326 ( .A(n4852), .B(n4772), .Z(n4896) );
  XOR U5327 ( .A(n4773), .B(n4769), .Z(n4772) );
  XNOR U5328 ( .A(n4900), .B(n4909), .Z(n4754) );
  XNOR U5329 ( .A(n4910), .B(n4911), .Z(n4909) );
  XOR U5330 ( .A(n4861), .B(n4846), .Z(n4852) );
  XNOR U5331 ( .A(n4850), .B(n4759), .Z(n4846) );
  IV U5332 ( .A(n4886), .Z(n4850) );
  XOR U5333 ( .A(n4912), .B(n4913), .Z(n4886) );
  XOR U5334 ( .A(n4914), .B(n4915), .Z(n4913) );
  XNOR U5335 ( .A(n4680), .B(n4916), .Z(n4912) );
  ANDN U5336 ( .B(n4773), .A(n4861), .Z(n4908) );
  XNOR U5337 ( .A(n4680), .B(n4842), .Z(n4861) );
  XOR U5338 ( .A(n4900), .B(n4890), .Z(n4773) );
  IV U5339 ( .A(n4762), .Z(n4890) );
  XOR U5340 ( .A(n4917), .B(n4918), .Z(n4762) );
  XOR U5341 ( .A(n4919), .B(n4915), .Z(n4918) );
  XNOR U5342 ( .A(n4920), .B(n4921), .Z(n4915) );
  XNOR U5343 ( .A(n4922), .B(n2971), .Z(n4921) );
  XOR U5344 ( .A(n3022), .B(n4253), .Z(n2971) );
  XNOR U5345 ( .A(n4923), .B(n4924), .Z(n4920) );
  XOR U5346 ( .A(key[1140]), .B(n4232), .Z(n4924) );
  IV U5347 ( .A(n4745), .Z(n4900) );
  XOR U5348 ( .A(n4893), .B(n4925), .Z(n4906) );
  XNOR U5349 ( .A(n4926), .B(n4899), .Z(n4925) );
  OR U5350 ( .A(n4743), .B(n4841), .Z(n4899) );
  XNOR U5351 ( .A(n4927), .B(n4759), .Z(n4841) );
  XNOR U5352 ( .A(n4745), .B(n4632), .Z(n4743) );
  ANDN U5353 ( .B(n4759), .A(n4632), .Z(n4926) );
  XOR U5354 ( .A(n4917), .B(n4928), .Z(n4632) );
  XOR U5355 ( .A(n4910), .B(n4929), .Z(n4928) );
  XOR U5356 ( .A(n4919), .B(n4917), .Z(n4759) );
  XNOR U5357 ( .A(n4842), .B(n4745), .Z(n4893) );
  XOR U5358 ( .A(n4917), .B(n4930), .Z(n4745) );
  XNOR U5359 ( .A(n4919), .B(n4914), .Z(n4930) );
  XOR U5360 ( .A(n4931), .B(n4932), .Z(n4914) );
  XOR U5361 ( .A(n4933), .B(n4934), .Z(n4932) );
  XNOR U5362 ( .A(key[1143]), .B(n4935), .Z(n4931) );
  XNOR U5363 ( .A(n4936), .B(n4937), .Z(n4917) );
  XOR U5364 ( .A(n4938), .B(n4939), .Z(n4937) );
  XNOR U5365 ( .A(key[1141]), .B(n4269), .Z(n4936) );
  XNOR U5366 ( .A(n2983), .B(n4940), .Z(n4269) );
  IV U5367 ( .A(n4927), .Z(n4842) );
  XNOR U5368 ( .A(n4911), .B(n4941), .Z(n4927) );
  XOR U5369 ( .A(n4916), .B(n4929), .Z(n4941) );
  IV U5370 ( .A(n4919), .Z(n4929) );
  XOR U5371 ( .A(n4942), .B(n4943), .Z(n4919) );
  XOR U5372 ( .A(n4944), .B(n2999), .Z(n4943) );
  XNOR U5373 ( .A(n3022), .B(n4248), .Z(n2999) );
  XOR U5374 ( .A(n4680), .B(n4945), .Z(n4942) );
  XNOR U5375 ( .A(key[1142]), .B(n4940), .Z(n4945) );
  XNOR U5376 ( .A(n4946), .B(n4947), .Z(n4680) );
  XOR U5377 ( .A(n3011), .B(n3021), .Z(n4947) );
  IV U5378 ( .A(n4948), .Z(n3021) );
  XOR U5379 ( .A(n4949), .B(n3020), .Z(n3011) );
  XOR U5380 ( .A(key[1136]), .B(n4950), .Z(n4946) );
  XOR U5381 ( .A(n4951), .B(n4952), .Z(n4916) );
  XNOR U5382 ( .A(n3007), .B(n4953), .Z(n4952) );
  XOR U5383 ( .A(n4910), .B(n4954), .Z(n4953) );
  XOR U5384 ( .A(n4955), .B(n4956), .Z(n4910) );
  XOR U5385 ( .A(n2994), .B(n4949), .Z(n4956) );
  XOR U5386 ( .A(n4957), .B(n3010), .Z(n2994) );
  XNOR U5387 ( .A(key[1137]), .B(n4277), .Z(n4955) );
  XNOR U5388 ( .A(n3022), .B(n4233), .Z(n3007) );
  XNOR U5389 ( .A(n4958), .B(n4959), .Z(n4951) );
  XNOR U5390 ( .A(key[1139]), .B(n4266), .Z(n4959) );
  IV U5391 ( .A(n4960), .Z(n4266) );
  XOR U5392 ( .A(n4961), .B(n4962), .Z(n4911) );
  XOR U5393 ( .A(n4262), .B(n3006), .Z(n4962) );
  IV U5394 ( .A(n4963), .Z(n4262) );
  XOR U5395 ( .A(key[1138]), .B(n4957), .Z(n4961) );
  XNOR U5396 ( .A(n1913), .B(n627), .Z(n642) );
  XOR U5397 ( .A(n4616), .B(n4964), .Z(n627) );
  XNOR U5398 ( .A(n4610), .B(n4649), .Z(n4964) );
  IV U5399 ( .A(n4611), .Z(n4649) );
  XOR U5400 ( .A(n4821), .B(n4965), .Z(n4611) );
  XNOR U5401 ( .A(n4819), .B(n4966), .Z(n4965) );
  NANDN U5402 ( .A(n4967), .B(n4704), .Z(n4966) );
  OR U5403 ( .A(n4968), .B(n4706), .Z(n4819) );
  XOR U5404 ( .A(n4622), .B(n4704), .Z(n4706) );
  XNOR U5405 ( .A(n4617), .B(n4969), .Z(n4610) );
  XNOR U5406 ( .A(n4970), .B(n4971), .Z(n4969) );
  NAND U5407 ( .A(n4972), .B(n4700), .Z(n4971) );
  XNOR U5408 ( .A(n4701), .B(n4973), .Z(n4617) );
  XNOR U5409 ( .A(n4974), .B(n4975), .Z(n4973) );
  NANDN U5410 ( .A(n4976), .B(n4825), .Z(n4975) );
  XOR U5411 ( .A(n4816), .B(n4608), .Z(n4616) );
  XNOR U5412 ( .A(n4701), .B(n4977), .Z(n4608) );
  XNOR U5413 ( .A(n4970), .B(n4978), .Z(n4977) );
  NANDN U5414 ( .A(n4979), .B(n4980), .Z(n4978) );
  OR U5415 ( .A(n4981), .B(n4982), .Z(n4970) );
  XOR U5416 ( .A(n4983), .B(n4974), .Z(n4701) );
  OR U5417 ( .A(n4984), .B(n4985), .Z(n4974) );
  ANDN U5418 ( .B(n4986), .A(n4987), .Z(n4983) );
  XOR U5419 ( .A(n4821), .B(n4988), .Z(n4816) );
  XOR U5420 ( .A(n4989), .B(n4697), .Z(n4988) );
  OR U5421 ( .A(n4990), .B(n4981), .Z(n4697) );
  XNOR U5422 ( .A(n4700), .B(n4980), .Z(n4981) );
  ANDN U5423 ( .B(n4980), .A(n4991), .Z(n4989) );
  XOR U5424 ( .A(n4992), .B(n4823), .Z(n4821) );
  OR U5425 ( .A(n4984), .B(n4993), .Z(n4823) );
  XNOR U5426 ( .A(n4986), .B(n4825), .Z(n4984) );
  XOR U5427 ( .A(n4704), .B(n4980), .Z(n4825) );
  XOR U5428 ( .A(n4994), .B(n4995), .Z(n4980) );
  NANDN U5429 ( .A(n4996), .B(n4997), .Z(n4995) );
  XOR U5430 ( .A(n4998), .B(n4999), .Z(n4704) );
  NANDN U5431 ( .A(n4996), .B(n5000), .Z(n4999) );
  AND U5432 ( .A(n5001), .B(n4986), .Z(n4992) );
  XNOR U5433 ( .A(n4622), .B(n4700), .Z(n4986) );
  XNOR U5434 ( .A(n5002), .B(n4994), .Z(n4700) );
  NANDN U5435 ( .A(n5003), .B(n5004), .Z(n4994) );
  XOR U5436 ( .A(n4997), .B(n5005), .Z(n5004) );
  ANDN U5437 ( .B(n5005), .A(n5006), .Z(n5002) );
  NANDN U5438 ( .A(n5003), .B(n5008), .Z(n4998) );
  XOR U5439 ( .A(n5009), .B(n5000), .Z(n5008) );
  XNOR U5440 ( .A(n5010), .B(n5011), .Z(n4996) );
  XOR U5441 ( .A(n5012), .B(n5013), .Z(n5011) );
  XNOR U5442 ( .A(n5014), .B(n5015), .Z(n5010) );
  XNOR U5443 ( .A(n5016), .B(n5017), .Z(n5015) );
  ANDN U5444 ( .B(n5009), .A(n5013), .Z(n5016) );
  ANDN U5445 ( .B(n5009), .A(n5006), .Z(n5007) );
  XNOR U5446 ( .A(n5012), .B(n5018), .Z(n5006) );
  XOR U5447 ( .A(n5019), .B(n5017), .Z(n5018) );
  NAND U5448 ( .A(n5020), .B(n5021), .Z(n5017) );
  XNOR U5449 ( .A(n5014), .B(n5000), .Z(n5021) );
  IV U5450 ( .A(n5009), .Z(n5014) );
  XNOR U5451 ( .A(n4997), .B(n5013), .Z(n5020) );
  IV U5452 ( .A(n5005), .Z(n5013) );
  XOR U5453 ( .A(n5022), .B(n5023), .Z(n5005) );
  XNOR U5454 ( .A(n5024), .B(n5025), .Z(n5023) );
  XNOR U5455 ( .A(n5026), .B(n5027), .Z(n5022) );
  ANDN U5456 ( .B(n4820), .A(n4621), .Z(n5026) );
  AND U5457 ( .A(n5000), .B(n4997), .Z(n5019) );
  XNOR U5458 ( .A(n5000), .B(n4997), .Z(n5012) );
  XNOR U5459 ( .A(n5028), .B(n5029), .Z(n4997) );
  XOR U5460 ( .A(n5030), .B(n5025), .Z(n5029) );
  XNOR U5461 ( .A(n5031), .B(n5032), .Z(n5028) );
  XNOR U5462 ( .A(n5033), .B(n5027), .Z(n5032) );
  OR U5463 ( .A(n4707), .B(n4968), .Z(n5027) );
  XNOR U5464 ( .A(n5034), .B(n4820), .Z(n4968) );
  XNOR U5465 ( .A(n4621), .B(n4705), .Z(n4707) );
  ANDN U5466 ( .B(n5035), .A(n4967), .Z(n5033) );
  XNOR U5467 ( .A(n5036), .B(n5037), .Z(n5000) );
  XNOR U5468 ( .A(n5025), .B(n5038), .Z(n5037) );
  XNOR U5469 ( .A(n4972), .B(n5030), .Z(n5038) );
  XNOR U5470 ( .A(n4621), .B(n4820), .Z(n5025) );
  XOR U5471 ( .A(n4699), .B(n5039), .Z(n5036) );
  XNOR U5472 ( .A(n5040), .B(n5041), .Z(n5039) );
  ANDN U5473 ( .B(n5042), .A(n4991), .Z(n5040) );
  XNOR U5474 ( .A(n5043), .B(n5044), .Z(n5009) );
  XNOR U5475 ( .A(n5024), .B(n5045), .Z(n5044) );
  XNOR U5476 ( .A(n5031), .B(n5046), .Z(n5045) );
  XNOR U5477 ( .A(n4705), .B(n5034), .Z(n5031) );
  XOR U5478 ( .A(n5030), .B(n5047), .Z(n5024) );
  XNOR U5479 ( .A(n5048), .B(n5049), .Z(n5047) );
  NANDN U5480 ( .A(n4976), .B(n4826), .Z(n5049) );
  XNOR U5481 ( .A(n5050), .B(n5048), .Z(n5030) );
  OR U5482 ( .A(n4993), .B(n4985), .Z(n5048) );
  XOR U5483 ( .A(n5051), .B(n4976), .Z(n4985) );
  XNOR U5484 ( .A(n5035), .B(n5042), .Z(n4976) );
  IV U5485 ( .A(n4705), .Z(n5035) );
  XOR U5486 ( .A(n5052), .B(n5053), .Z(n4705) );
  XNOR U5487 ( .A(n5001), .B(n4826), .Z(n4993) );
  XNOR U5488 ( .A(n4967), .B(n5046), .Z(n4826) );
  IV U5489 ( .A(n5034), .Z(n4967) );
  XOR U5490 ( .A(n5054), .B(n5055), .Z(n5034) );
  ANDN U5491 ( .B(n5001), .A(n4987), .Z(n5050) );
  IV U5492 ( .A(n5051), .Z(n4987) );
  XNOR U5493 ( .A(n4979), .B(n5056), .Z(n5043) );
  XNOR U5494 ( .A(n5057), .B(n5041), .Z(n5056) );
  OR U5495 ( .A(n4982), .B(n4990), .Z(n5041) );
  XNOR U5496 ( .A(n4699), .B(n4991), .Z(n4990) );
  IV U5497 ( .A(n5046), .Z(n4991) );
  XOR U5498 ( .A(n5058), .B(n5059), .Z(n5046) );
  XNOR U5499 ( .A(n5060), .B(n5061), .Z(n5059) );
  XNOR U5500 ( .A(n5062), .B(n4699), .Z(n5058) );
  XNOR U5501 ( .A(n4972), .B(n5042), .Z(n4982) );
  IV U5502 ( .A(n4979), .Z(n5042) );
  ANDN U5503 ( .B(n4972), .A(n4699), .Z(n5057) );
  XOR U5504 ( .A(n5060), .B(n5053), .Z(n4972) );
  XNOR U5505 ( .A(n5054), .B(n5063), .Z(n5053) );
  XOR U5506 ( .A(n5064), .B(n5065), .Z(n5060) );
  XNOR U5507 ( .A(n2810), .B(n5066), .Z(n5064) );
  XOR U5508 ( .A(key[1060]), .B(n5067), .Z(n5066) );
  XOR U5509 ( .A(n5068), .B(n3778), .Z(n2810) );
  XNOR U5510 ( .A(n5069), .B(n5070), .Z(n4979) );
  XOR U5511 ( .A(n4621), .B(n5052), .Z(n5070) );
  XOR U5512 ( .A(n5063), .B(n5071), .Z(n4621) );
  XOR U5513 ( .A(n5062), .B(n5054), .Z(n5071) );
  XNOR U5514 ( .A(n5072), .B(n5073), .Z(n5054) );
  XNOR U5515 ( .A(n3779), .B(n5074), .Z(n5073) );
  XNOR U5516 ( .A(key[1061]), .B(n3773), .Z(n5072) );
  XNOR U5517 ( .A(n2799), .B(n5075), .Z(n3773) );
  XOR U5518 ( .A(n5076), .B(n5077), .Z(n5062) );
  XNOR U5519 ( .A(n5078), .B(n5079), .Z(n5077) );
  XNOR U5520 ( .A(key[1063]), .B(n5068), .Z(n5076) );
  IV U5521 ( .A(n2833), .Z(n5068) );
  IV U5522 ( .A(n5055), .Z(n5063) );
  XNOR U5523 ( .A(n4699), .B(n4820), .Z(n5001) );
  XNOR U5524 ( .A(n5061), .B(n5080), .Z(n4820) );
  XNOR U5525 ( .A(n5055), .B(n5069), .Z(n5080) );
  XOR U5526 ( .A(n5081), .B(n5082), .Z(n5069) );
  XNOR U5527 ( .A(n3803), .B(n5083), .Z(n5082) );
  XNOR U5528 ( .A(key[1058]), .B(n3805), .Z(n5081) );
  IV U5529 ( .A(n2828), .Z(n3805) );
  XOR U5530 ( .A(n2782), .B(n5084), .Z(n2828) );
  XOR U5531 ( .A(n5085), .B(n5086), .Z(n5055) );
  XNOR U5532 ( .A(n2789), .B(n5087), .Z(n5086) );
  XNOR U5533 ( .A(n2833), .B(n3786), .Z(n2789) );
  XOR U5534 ( .A(n4699), .B(n5088), .Z(n5085) );
  XNOR U5535 ( .A(key[1062]), .B(n5075), .Z(n5088) );
  XOR U5536 ( .A(n5089), .B(n5090), .Z(n5061) );
  XNOR U5537 ( .A(n2818), .B(n5091), .Z(n5090) );
  XNOR U5538 ( .A(n5052), .B(n5092), .Z(n5091) );
  XNOR U5539 ( .A(n5093), .B(n5094), .Z(n5052) );
  XNOR U5540 ( .A(n5095), .B(n2779), .Z(n5094) );
  XNOR U5541 ( .A(n5096), .B(n2822), .Z(n2779) );
  XNOR U5542 ( .A(key[1057]), .B(n3808), .Z(n5093) );
  XNOR U5543 ( .A(n2833), .B(n3794), .Z(n2818) );
  XNOR U5544 ( .A(n3764), .B(n5097), .Z(n5089) );
  XNOR U5545 ( .A(key[1059]), .B(n5084), .Z(n5097) );
  IV U5546 ( .A(n5098), .Z(n3764) );
  XNOR U5547 ( .A(n5099), .B(n5100), .Z(n4699) );
  XOR U5548 ( .A(n2823), .B(n2832), .Z(n5100) );
  XNOR U5549 ( .A(n5101), .B(n2831), .Z(n2823) );
  XNOR U5550 ( .A(key[1056]), .B(n3787), .Z(n5099) );
  IV U5551 ( .A(n4801), .Z(n1913) );
  XOR U5552 ( .A(n4684), .B(n5102), .Z(n4801) );
  XNOR U5553 ( .A(n4656), .B(n4803), .Z(n5102) );
  IV U5554 ( .A(n4686), .Z(n4803) );
  XNOR U5555 ( .A(n4833), .B(n5103), .Z(n4686) );
  XNOR U5556 ( .A(n4831), .B(n5104), .Z(n5103) );
  NAND U5557 ( .A(n4722), .B(n5105), .Z(n5104) );
  OR U5558 ( .A(n5106), .B(n4811), .Z(n4831) );
  XOR U5559 ( .A(n4814), .B(n4722), .Z(n4811) );
  XOR U5560 ( .A(n4802), .B(n4815), .Z(n4656) );
  XNOR U5561 ( .A(n4718), .B(n5107), .Z(n4815) );
  XNOR U5562 ( .A(n5108), .B(n5109), .Z(n5107) );
  NANDN U5563 ( .A(n5110), .B(n5111), .Z(n5109) );
  XNOR U5564 ( .A(n4833), .B(n5112), .Z(n4802) );
  XNOR U5565 ( .A(n5113), .B(n4714), .Z(n5112) );
  NOR U5566 ( .A(n5114), .B(n5115), .Z(n4714) );
  ANDN U5567 ( .B(n5111), .A(n5116), .Z(n5113) );
  XOR U5568 ( .A(n5117), .B(n4835), .Z(n4833) );
  OR U5569 ( .A(n5118), .B(n5119), .Z(n4835) );
  ANDN U5570 ( .B(n5120), .A(n5121), .Z(n5117) );
  IV U5571 ( .A(n4807), .Z(n4684) );
  XNOR U5572 ( .A(n5108), .B(n5123), .Z(n5122) );
  NANDN U5573 ( .A(n5124), .B(n4717), .Z(n5123) );
  OR U5574 ( .A(n5125), .B(n5114), .Z(n5108) );
  XNOR U5575 ( .A(n4717), .B(n5111), .Z(n5114) );
  XNOR U5576 ( .A(n4718), .B(n5126), .Z(n4808) );
  XNOR U5577 ( .A(n5127), .B(n5128), .Z(n5126) );
  NANDN U5578 ( .A(n4837), .B(n5129), .Z(n5128) );
  XOR U5579 ( .A(n5130), .B(n5127), .Z(n4718) );
  NANDN U5580 ( .A(n5118), .B(n5131), .Z(n5127) );
  XOR U5581 ( .A(n5120), .B(n4837), .Z(n5118) );
  XNOR U5582 ( .A(n4722), .B(n5111), .Z(n4837) );
  XOR U5583 ( .A(n5132), .B(n5133), .Z(n5111) );
  NANDN U5584 ( .A(n5134), .B(n5135), .Z(n5133) );
  XOR U5585 ( .A(n5136), .B(n5137), .Z(n4722) );
  NANDN U5586 ( .A(n5134), .B(n5138), .Z(n5137) );
  AND U5587 ( .A(n5139), .B(n5120), .Z(n5130) );
  XNOR U5588 ( .A(n4814), .B(n4717), .Z(n5120) );
  XNOR U5589 ( .A(n5140), .B(n5132), .Z(n4717) );
  NANDN U5590 ( .A(n5141), .B(n5142), .Z(n5132) );
  XOR U5591 ( .A(n5135), .B(n5143), .Z(n5142) );
  ANDN U5592 ( .B(n5143), .A(n5144), .Z(n5140) );
  NANDN U5593 ( .A(n5141), .B(n5146), .Z(n5136) );
  XOR U5594 ( .A(n5147), .B(n5138), .Z(n5146) );
  XNOR U5595 ( .A(n5148), .B(n5149), .Z(n5134) );
  XOR U5596 ( .A(n5150), .B(n5151), .Z(n5149) );
  XNOR U5597 ( .A(n5152), .B(n5153), .Z(n5148) );
  XNOR U5598 ( .A(n5154), .B(n5155), .Z(n5153) );
  ANDN U5599 ( .B(n5147), .A(n5151), .Z(n5154) );
  ANDN U5600 ( .B(n5147), .A(n5144), .Z(n5145) );
  XNOR U5601 ( .A(n5150), .B(n5156), .Z(n5144) );
  XOR U5602 ( .A(n5157), .B(n5155), .Z(n5156) );
  NAND U5603 ( .A(n5158), .B(n5159), .Z(n5155) );
  XNOR U5604 ( .A(n5152), .B(n5138), .Z(n5159) );
  IV U5605 ( .A(n5147), .Z(n5152) );
  XNOR U5606 ( .A(n5135), .B(n5151), .Z(n5158) );
  IV U5607 ( .A(n5143), .Z(n5151) );
  XOR U5608 ( .A(n5160), .B(n5161), .Z(n5143) );
  XNOR U5609 ( .A(n5162), .B(n5163), .Z(n5161) );
  XNOR U5610 ( .A(n5164), .B(n5165), .Z(n5160) );
  ANDN U5611 ( .B(n5166), .A(n4832), .Z(n5164) );
  AND U5612 ( .A(n5138), .B(n5135), .Z(n5157) );
  XNOR U5613 ( .A(n5138), .B(n5135), .Z(n5150) );
  XNOR U5614 ( .A(n5167), .B(n5168), .Z(n5135) );
  XOR U5615 ( .A(n5169), .B(n5163), .Z(n5168) );
  XNOR U5616 ( .A(n5170), .B(n5171), .Z(n5167) );
  XNOR U5617 ( .A(n5172), .B(n5165), .Z(n5171) );
  OR U5618 ( .A(n4812), .B(n5106), .Z(n5165) );
  XNOR U5619 ( .A(n5173), .B(n5105), .Z(n5106) );
  XNOR U5620 ( .A(n4723), .B(n4813), .Z(n4812) );
  ANDN U5621 ( .B(n5105), .A(n4723), .Z(n5172) );
  XNOR U5622 ( .A(n5174), .B(n5175), .Z(n5138) );
  XNOR U5623 ( .A(n5163), .B(n5176), .Z(n5175) );
  XOR U5624 ( .A(n5124), .B(n5169), .Z(n5176) );
  XNOR U5625 ( .A(n5173), .B(n4813), .Z(n5163) );
  XOR U5626 ( .A(n4716), .B(n5177), .Z(n5174) );
  XNOR U5627 ( .A(n5178), .B(n5179), .Z(n5177) );
  XNOR U5628 ( .A(n5180), .B(n5181), .Z(n5147) );
  XNOR U5629 ( .A(n5162), .B(n5182), .Z(n5181) );
  XNOR U5630 ( .A(n5170), .B(n5110), .Z(n5182) );
  XOR U5631 ( .A(n5105), .B(n5183), .Z(n5170) );
  XOR U5632 ( .A(n5169), .B(n5184), .Z(n5162) );
  XNOR U5633 ( .A(n5185), .B(n5186), .Z(n5184) );
  NAND U5634 ( .A(n4838), .B(n5129), .Z(n5186) );
  XNOR U5635 ( .A(n5187), .B(n5185), .Z(n5169) );
  NANDN U5636 ( .A(n5119), .B(n5131), .Z(n5185) );
  XOR U5637 ( .A(n5139), .B(n5129), .Z(n5131) );
  XNOR U5638 ( .A(n5183), .B(n5110), .Z(n5129) );
  IV U5639 ( .A(n4723), .Z(n5183) );
  XOR U5640 ( .A(n5188), .B(n5189), .Z(n4723) );
  XOR U5641 ( .A(n5190), .B(n5191), .Z(n5189) );
  XOR U5642 ( .A(n5121), .B(n4838), .Z(n5119) );
  XOR U5643 ( .A(n5105), .B(n5192), .Z(n4838) );
  ANDN U5644 ( .B(n5139), .A(n5121), .Z(n5187) );
  XOR U5645 ( .A(n4716), .B(n5173), .Z(n5121) );
  IV U5646 ( .A(n4832), .Z(n5173) );
  XOR U5647 ( .A(n5193), .B(n5194), .Z(n4832) );
  XOR U5648 ( .A(n5195), .B(n5190), .Z(n5194) );
  XNOR U5649 ( .A(n5192), .B(n5196), .Z(n5180) );
  XNOR U5650 ( .A(n5197), .B(n5179), .Z(n5196) );
  OR U5651 ( .A(n5125), .B(n5115), .Z(n5179) );
  XNOR U5652 ( .A(n4716), .B(n5116), .Z(n5115) );
  IV U5653 ( .A(n5192), .Z(n5116) );
  XNOR U5654 ( .A(n5124), .B(n5110), .Z(n5125) );
  XOR U5655 ( .A(n5166), .B(n5198), .Z(n5110) );
  XNOR U5656 ( .A(n5195), .B(n5191), .Z(n5198) );
  XOR U5657 ( .A(n5199), .B(n5200), .Z(n5195) );
  XNOR U5658 ( .A(n3931), .B(n2643), .Z(n5200) );
  IV U5659 ( .A(n5201), .Z(n2643) );
  XNOR U5660 ( .A(n2684), .B(n5202), .Z(n5199) );
  XOR U5661 ( .A(key[1050]), .B(n3940), .Z(n5202) );
  NOR U5662 ( .A(n5124), .B(n4716), .Z(n5197) );
  IV U5663 ( .A(n5203), .Z(n5124) );
  XOR U5664 ( .A(n5204), .B(n5205), .Z(n5192) );
  XNOR U5665 ( .A(n5206), .B(n5207), .Z(n5205) );
  XNOR U5666 ( .A(n4716), .B(n5193), .Z(n5204) );
  XOR U5667 ( .A(n5208), .B(n5209), .Z(n5193) );
  XNOR U5668 ( .A(n2676), .B(n5210), .Z(n5209) );
  XOR U5669 ( .A(n2675), .B(n5211), .Z(n5210) );
  XOR U5670 ( .A(n5212), .B(n5213), .Z(n2676) );
  XNOR U5671 ( .A(n5191), .B(n5214), .Z(n5208) );
  XNOR U5672 ( .A(key[1051]), .B(n3917), .Z(n5214) );
  XOR U5673 ( .A(n5215), .B(n5216), .Z(n5191) );
  XOR U5674 ( .A(n3943), .B(n2680), .Z(n5216) );
  XOR U5675 ( .A(n3919), .B(n5217), .Z(n5215) );
  XOR U5676 ( .A(key[1049]), .B(n2644), .Z(n5217) );
  XOR U5677 ( .A(n5203), .B(n5166), .Z(n5139) );
  IV U5678 ( .A(n4813), .Z(n5166) );
  XNOR U5679 ( .A(n5207), .B(n5105), .Z(n4813) );
  XOR U5680 ( .A(n5218), .B(n5219), .Z(n5207) );
  XNOR U5681 ( .A(n5220), .B(n2665), .Z(n5219) );
  XNOR U5682 ( .A(n5221), .B(n3911), .Z(n2665) );
  XOR U5683 ( .A(key[1055]), .B(n2687), .Z(n5218) );
  XOR U5684 ( .A(n5222), .B(n5213), .Z(n2687) );
  XOR U5685 ( .A(n5206), .B(n5105), .Z(n5203) );
  XNOR U5686 ( .A(n5190), .B(n5188), .Z(n5105) );
  XNOR U5687 ( .A(n5223), .B(n5224), .Z(n5188) );
  XNOR U5688 ( .A(n5225), .B(n2658), .Z(n5224) );
  XNOR U5689 ( .A(n3904), .B(n5226), .Z(n2658) );
  XOR U5690 ( .A(n3926), .B(n5227), .Z(n5223) );
  XNOR U5691 ( .A(key[1053]), .B(n3896), .Z(n5227) );
  XNOR U5692 ( .A(n5228), .B(n5229), .Z(n5190) );
  XOR U5693 ( .A(n5230), .B(n2651), .Z(n5229) );
  XOR U5694 ( .A(n5231), .B(n2664), .Z(n2651) );
  XNOR U5695 ( .A(n5213), .B(n5232), .Z(n2664) );
  XOR U5696 ( .A(n4716), .B(n5233), .Z(n5228) );
  XNOR U5697 ( .A(key[1054]), .B(n3905), .Z(n5233) );
  XNOR U5698 ( .A(n5234), .B(n5235), .Z(n4716) );
  XOR U5699 ( .A(n5236), .B(n3937), .Z(n5235) );
  XOR U5700 ( .A(n3910), .B(n5237), .Z(n5234) );
  XNOR U5701 ( .A(key[1048]), .B(n5238), .Z(n5237) );
  XOR U5702 ( .A(n5239), .B(n2668), .Z(n5206) );
  XOR U5703 ( .A(n5240), .B(n5241), .Z(n2668) );
  XOR U5704 ( .A(n3895), .B(n5242), .Z(n5241) );
  XOR U5705 ( .A(n2659), .B(n5213), .Z(n5240) );
  XNOR U5706 ( .A(n5243), .B(n5244), .Z(n5239) );
  XNOR U5707 ( .A(key[1052]), .B(n3932), .Z(n5244) );
  XNOR U5708 ( .A(key[1152]), .B(n1266), .Z(n4827) );
  XNOR U5709 ( .A(n4665), .B(n5245), .Z(n4637) );
  XNOR U5710 ( .A(n5246), .B(n4783), .Z(n5245) );
  XOR U5711 ( .A(n4734), .B(n4641), .Z(n4732) );
  ANDN U5712 ( .B(n4734), .A(n5248), .Z(n5246) );
  XNOR U5713 ( .A(n4781), .B(n5249), .Z(n4665) );
  XNOR U5714 ( .A(n5250), .B(n5251), .Z(n5249) );
  NANDN U5715 ( .A(n4794), .B(n5252), .Z(n5251) );
  XNOR U5716 ( .A(n4781), .B(n5253), .Z(n4691) );
  XOR U5717 ( .A(n5254), .B(n4667), .Z(n5253) );
  OR U5718 ( .A(n5255), .B(n4789), .Z(n4667) );
  XNOR U5719 ( .A(n4669), .B(n4779), .Z(n4789) );
  NOR U5720 ( .A(n5256), .B(n4779), .Z(n5254) );
  XOR U5721 ( .A(n5257), .B(n5250), .Z(n4781) );
  OR U5722 ( .A(n4797), .B(n5258), .Z(n5250) );
  XOR U5723 ( .A(n5259), .B(n4794), .Z(n4797) );
  XOR U5724 ( .A(n4779), .B(n4641), .Z(n4794) );
  XOR U5725 ( .A(n5260), .B(n5261), .Z(n4641) );
  NANDN U5726 ( .A(n5262), .B(n5263), .Z(n5261) );
  XNOR U5727 ( .A(n5264), .B(n5265), .Z(n4779) );
  OR U5728 ( .A(n5262), .B(n5266), .Z(n5265) );
  ANDN U5729 ( .B(n5259), .A(n5267), .Z(n5257) );
  IV U5730 ( .A(n4800), .Z(n5259) );
  XOR U5731 ( .A(n4669), .B(n4734), .Z(n4800) );
  XNOR U5732 ( .A(n5268), .B(n5260), .Z(n4734) );
  NANDN U5733 ( .A(n5269), .B(n5270), .Z(n5260) );
  ANDN U5734 ( .B(n5271), .A(n5272), .Z(n5268) );
  NANDN U5735 ( .A(n5269), .B(n5274), .Z(n5264) );
  XOR U5736 ( .A(n5275), .B(n5262), .Z(n5269) );
  XNOR U5737 ( .A(n5276), .B(n5277), .Z(n5262) );
  XOR U5738 ( .A(n5278), .B(n5271), .Z(n5277) );
  XNOR U5739 ( .A(n5279), .B(n5280), .Z(n5276) );
  XNOR U5740 ( .A(n5281), .B(n5282), .Z(n5280) );
  ANDN U5741 ( .B(n5271), .A(n5283), .Z(n5281) );
  IV U5742 ( .A(n5284), .Z(n5271) );
  ANDN U5743 ( .B(n5275), .A(n5283), .Z(n5273) );
  IV U5744 ( .A(n5279), .Z(n5283) );
  IV U5745 ( .A(n5272), .Z(n5275) );
  XNOR U5746 ( .A(n5278), .B(n5285), .Z(n5272) );
  XOR U5747 ( .A(n5286), .B(n5282), .Z(n5285) );
  NAND U5748 ( .A(n5274), .B(n5270), .Z(n5282) );
  XNOR U5749 ( .A(n5263), .B(n5284), .Z(n5270) );
  XOR U5750 ( .A(n5287), .B(n5288), .Z(n5284) );
  XOR U5751 ( .A(n5289), .B(n5290), .Z(n5288) );
  XNOR U5752 ( .A(n4780), .B(n5291), .Z(n5290) );
  XNOR U5753 ( .A(n5292), .B(n5293), .Z(n5287) );
  XNOR U5754 ( .A(n5294), .B(n5295), .Z(n5293) );
  ANDN U5755 ( .B(n5296), .A(n4670), .Z(n5294) );
  XNOR U5756 ( .A(n5279), .B(n5266), .Z(n5274) );
  XOR U5757 ( .A(n5297), .B(n5298), .Z(n5279) );
  XNOR U5758 ( .A(n5299), .B(n5291), .Z(n5298) );
  XOR U5759 ( .A(n5300), .B(n5301), .Z(n5291) );
  XNOR U5760 ( .A(n5302), .B(n5303), .Z(n5301) );
  NAND U5761 ( .A(n5252), .B(n4795), .Z(n5303) );
  XNOR U5762 ( .A(n5304), .B(n5305), .Z(n5297) );
  ANDN U5763 ( .B(n5306), .A(n5248), .Z(n5304) );
  ANDN U5764 ( .B(n5263), .A(n5266), .Z(n5286) );
  XOR U5765 ( .A(n5266), .B(n5263), .Z(n5278) );
  XNOR U5766 ( .A(n5307), .B(n5308), .Z(n5263) );
  XNOR U5767 ( .A(n5300), .B(n5309), .Z(n5308) );
  XOR U5768 ( .A(n5299), .B(n4788), .Z(n5309) );
  XOR U5769 ( .A(n4670), .B(n5310), .Z(n5307) );
  XNOR U5770 ( .A(n5311), .B(n5295), .Z(n5310) );
  OR U5771 ( .A(n4790), .B(n5255), .Z(n5295) );
  XNOR U5772 ( .A(n4670), .B(n5256), .Z(n5255) );
  XOR U5773 ( .A(n4788), .B(n4780), .Z(n4790) );
  ANDN U5774 ( .B(n4780), .A(n5256), .Z(n5311) );
  XOR U5775 ( .A(n5312), .B(n5313), .Z(n5266) );
  XOR U5776 ( .A(n5300), .B(n5289), .Z(n5313) );
  XOR U5777 ( .A(n4785), .B(n4642), .Z(n5289) );
  XOR U5778 ( .A(n5314), .B(n5302), .Z(n5300) );
  NANDN U5779 ( .A(n5258), .B(n4798), .Z(n5302) );
  XOR U5780 ( .A(n4799), .B(n4795), .Z(n4798) );
  XNOR U5781 ( .A(n5306), .B(n5315), .Z(n4780) );
  XNOR U5782 ( .A(n5316), .B(n5317), .Z(n5315) );
  XOR U5783 ( .A(n5267), .B(n5252), .Z(n5258) );
  XNOR U5784 ( .A(n5256), .B(n4785), .Z(n5252) );
  IV U5785 ( .A(n5292), .Z(n5256) );
  XOR U5786 ( .A(n5318), .B(n5319), .Z(n5292) );
  XOR U5787 ( .A(n5320), .B(n5321), .Z(n5319) );
  XNOR U5788 ( .A(n4670), .B(n5322), .Z(n5318) );
  ANDN U5789 ( .B(n4799), .A(n5267), .Z(n5314) );
  XNOR U5790 ( .A(n4670), .B(n5248), .Z(n5267) );
  XOR U5791 ( .A(n5306), .B(n5296), .Z(n4799) );
  IV U5792 ( .A(n4788), .Z(n5296) );
  XOR U5793 ( .A(n5323), .B(n5324), .Z(n4788) );
  XOR U5794 ( .A(n5325), .B(n5321), .Z(n5324) );
  XNOR U5795 ( .A(n5326), .B(n3139), .Z(n5321) );
  XOR U5796 ( .A(n5327), .B(n5328), .Z(n3139) );
  XOR U5797 ( .A(n5329), .B(n4097), .Z(n5328) );
  XOR U5798 ( .A(n5330), .B(n3128), .Z(n5327) );
  XNOR U5799 ( .A(n5331), .B(n5332), .Z(n5326) );
  XNOR U5800 ( .A(key[1100]), .B(n4115), .Z(n5332) );
  IV U5801 ( .A(n4735), .Z(n5306) );
  XOR U5802 ( .A(n5299), .B(n5333), .Z(n5312) );
  XNOR U5803 ( .A(n5334), .B(n5305), .Z(n5333) );
  OR U5804 ( .A(n4733), .B(n5247), .Z(n5305) );
  XNOR U5805 ( .A(n5335), .B(n4785), .Z(n5247) );
  XNOR U5806 ( .A(n4735), .B(n4642), .Z(n4733) );
  ANDN U5807 ( .B(n4785), .A(n4642), .Z(n5334) );
  XOR U5808 ( .A(n5323), .B(n5336), .Z(n4642) );
  XOR U5809 ( .A(n5316), .B(n5337), .Z(n5336) );
  XOR U5810 ( .A(n5325), .B(n5323), .Z(n4785) );
  XNOR U5811 ( .A(n5248), .B(n4735), .Z(n5299) );
  XOR U5812 ( .A(n5323), .B(n5338), .Z(n4735) );
  XNOR U5813 ( .A(n5325), .B(n5320), .Z(n5338) );
  XOR U5814 ( .A(n5339), .B(n5340), .Z(n5320) );
  XNOR U5815 ( .A(n4078), .B(n3136), .Z(n5340) );
  XNOR U5816 ( .A(n5341), .B(n4093), .Z(n3136) );
  XNOR U5817 ( .A(key[1103]), .B(n3160), .Z(n5339) );
  XOR U5818 ( .A(n5342), .B(n5330), .Z(n3160) );
  XNOR U5819 ( .A(n5343), .B(n5344), .Z(n5323) );
  XOR U5820 ( .A(n4101), .B(n3129), .Z(n5344) );
  XNOR U5821 ( .A(n5345), .B(n4083), .Z(n3129) );
  XNOR U5822 ( .A(n3123), .B(n5346), .Z(n5343) );
  XNOR U5823 ( .A(key[1101]), .B(n4079), .Z(n5346) );
  IV U5824 ( .A(n5335), .Z(n5248) );
  XNOR U5825 ( .A(n5317), .B(n5347), .Z(n5335) );
  XOR U5826 ( .A(n5322), .B(n5337), .Z(n5347) );
  IV U5827 ( .A(n5325), .Z(n5337) );
  XOR U5828 ( .A(n5348), .B(n5349), .Z(n5325) );
  XNOR U5829 ( .A(n5350), .B(n3122), .Z(n5349) );
  XNOR U5830 ( .A(n5351), .B(n3135), .Z(n3122) );
  XOR U5831 ( .A(n5330), .B(n5352), .Z(n3135) );
  XOR U5832 ( .A(n4670), .B(n5353), .Z(n5348) );
  XOR U5833 ( .A(key[1102]), .B(n4087), .Z(n5353) );
  XNOR U5834 ( .A(n5354), .B(n5355), .Z(n4670) );
  XOR U5835 ( .A(n5356), .B(n4092), .Z(n5355) );
  XOR U5836 ( .A(n4109), .B(n5357), .Z(n5354) );
  XNOR U5837 ( .A(key[1096]), .B(n5358), .Z(n5357) );
  XOR U5838 ( .A(n5359), .B(n5360), .Z(n5322) );
  XNOR U5839 ( .A(n3147), .B(n5361), .Z(n5360) );
  XNOR U5840 ( .A(n5316), .B(n3146), .Z(n5361) );
  XOR U5841 ( .A(n5330), .B(n3140), .Z(n3146) );
  XOR U5842 ( .A(n5362), .B(n5363), .Z(n5316) );
  XNOR U5843 ( .A(n4065), .B(n3151), .Z(n5363) );
  XOR U5844 ( .A(n3113), .B(n5364), .Z(n5362) );
  XNOR U5845 ( .A(key[1097]), .B(n4118), .Z(n5364) );
  XNOR U5846 ( .A(n5365), .B(n5366), .Z(n5359) );
  XNOR U5847 ( .A(key[1099]), .B(n4069), .Z(n5366) );
  XOR U5848 ( .A(n5367), .B(n5368), .Z(n5317) );
  XOR U5849 ( .A(n4104), .B(n3114), .Z(n5368) );
  XNOR U5850 ( .A(n3153), .B(n5369), .Z(n5367) );
  XOR U5851 ( .A(key[1098]), .B(n4111), .Z(n5369) );
  XNOR U5852 ( .A(n887), .B(n5370), .Z(out[0]) );
  XOR U5853 ( .A(key[1152]), .B(n1721), .Z(n5370) );
  XNOR U5854 ( .A(n1962), .B(n5371), .Z(n1721) );
  XOR U5855 ( .A(n5372), .B(n891), .Z(n5371) );
  OR U5856 ( .A(n5373), .B(n1955), .Z(n891) );
  XNOR U5857 ( .A(n894), .B(n1954), .Z(n1955) );
  ANDN U5858 ( .B(n1954), .A(n5374), .Z(n5372) );
  IV U5859 ( .A(n1127), .Z(n887) );
  XOR U5860 ( .A(n895), .B(n5375), .Z(n1127) );
  XOR U5861 ( .A(n5376), .B(n1964), .Z(n5375) );
  XNOR U5862 ( .A(n1507), .B(n899), .Z(n1504) );
  NOR U5863 ( .A(n5378), .B(n1507), .Z(n5376) );
  XNOR U5864 ( .A(n1962), .B(n5379), .Z(n895) );
  XNOR U5865 ( .A(n5380), .B(n5381), .Z(n5379) );
  NANDN U5866 ( .A(n1949), .B(n5382), .Z(n5381) );
  XOR U5867 ( .A(n5383), .B(n5380), .Z(n1962) );
  OR U5868 ( .A(n1958), .B(n5384), .Z(n5380) );
  XOR U5869 ( .A(n5385), .B(n1949), .Z(n1958) );
  XNOR U5870 ( .A(n1954), .B(n899), .Z(n1949) );
  XOR U5871 ( .A(n5386), .B(n5387), .Z(n899) );
  NANDN U5872 ( .A(n5388), .B(n5389), .Z(n5387) );
  XOR U5873 ( .A(n5390), .B(n5391), .Z(n1954) );
  NANDN U5874 ( .A(n5388), .B(n5392), .Z(n5391) );
  ANDN U5875 ( .B(n5385), .A(n5393), .Z(n5383) );
  IV U5876 ( .A(n1961), .Z(n5385) );
  XOR U5877 ( .A(n1507), .B(n894), .Z(n1961) );
  XNOR U5878 ( .A(n5394), .B(n5390), .Z(n894) );
  NANDN U5879 ( .A(n5395), .B(n5396), .Z(n5390) );
  XOR U5880 ( .A(n5392), .B(n5397), .Z(n5396) );
  ANDN U5881 ( .B(n5397), .A(n5398), .Z(n5394) );
  XOR U5882 ( .A(n5399), .B(n5386), .Z(n1507) );
  NANDN U5883 ( .A(n5395), .B(n5400), .Z(n5386) );
  XOR U5884 ( .A(n5401), .B(n5389), .Z(n5400) );
  XNOR U5885 ( .A(n5402), .B(n5403), .Z(n5388) );
  XOR U5886 ( .A(n5404), .B(n5405), .Z(n5403) );
  XNOR U5887 ( .A(n5406), .B(n5407), .Z(n5402) );
  XNOR U5888 ( .A(n5408), .B(n5409), .Z(n5407) );
  ANDN U5889 ( .B(n5401), .A(n5405), .Z(n5408) );
  ANDN U5890 ( .B(n5401), .A(n5398), .Z(n5399) );
  XNOR U5891 ( .A(n5404), .B(n5410), .Z(n5398) );
  XOR U5892 ( .A(n5411), .B(n5409), .Z(n5410) );
  NAND U5893 ( .A(n5412), .B(n5413), .Z(n5409) );
  XNOR U5894 ( .A(n5406), .B(n5389), .Z(n5413) );
  IV U5895 ( .A(n5401), .Z(n5406) );
  XNOR U5896 ( .A(n5392), .B(n5405), .Z(n5412) );
  IV U5897 ( .A(n5397), .Z(n5405) );
  XOR U5898 ( .A(n5414), .B(n5415), .Z(n5397) );
  XNOR U5899 ( .A(n5416), .B(n5417), .Z(n5415) );
  XNOR U5900 ( .A(n5418), .B(n5419), .Z(n5414) );
  NOR U5901 ( .A(n1506), .B(n5378), .Z(n5418) );
  AND U5902 ( .A(n5389), .B(n5392), .Z(n5411) );
  XNOR U5903 ( .A(n5389), .B(n5392), .Z(n5404) );
  XNOR U5904 ( .A(n5420), .B(n5421), .Z(n5392) );
  XNOR U5905 ( .A(n5422), .B(n5417), .Z(n5421) );
  XOR U5906 ( .A(n5423), .B(n5424), .Z(n5420) );
  XNOR U5907 ( .A(n5425), .B(n5419), .Z(n5424) );
  OR U5908 ( .A(n1505), .B(n5377), .Z(n5419) );
  XNOR U5909 ( .A(n5378), .B(n1966), .Z(n5377) );
  XNOR U5910 ( .A(n1506), .B(n900), .Z(n1505) );
  ANDN U5911 ( .B(n5426), .A(n1966), .Z(n5425) );
  XNOR U5912 ( .A(n5427), .B(n5428), .Z(n5389) );
  XNOR U5913 ( .A(n5417), .B(n5429), .Z(n5428) );
  XOR U5914 ( .A(n1945), .B(n5423), .Z(n5429) );
  XNOR U5915 ( .A(n5378), .B(n5430), .Z(n5417) );
  XOR U5916 ( .A(n893), .B(n5431), .Z(n5427) );
  XNOR U5917 ( .A(n5432), .B(n5433), .Z(n5431) );
  ANDN U5918 ( .B(n5434), .A(n5374), .Z(n5432) );
  XNOR U5919 ( .A(n5435), .B(n5436), .Z(n5401) );
  XNOR U5920 ( .A(n5422), .B(n5437), .Z(n5436) );
  XNOR U5921 ( .A(n1953), .B(n5416), .Z(n5437) );
  XOR U5922 ( .A(n5423), .B(n5438), .Z(n5416) );
  XNOR U5923 ( .A(n5439), .B(n5440), .Z(n5438) );
  NAND U5924 ( .A(n5382), .B(n1950), .Z(n5440) );
  XNOR U5925 ( .A(n5441), .B(n5439), .Z(n5423) );
  NANDN U5926 ( .A(n5384), .B(n1959), .Z(n5439) );
  XOR U5927 ( .A(n1960), .B(n1950), .Z(n1959) );
  XNOR U5928 ( .A(n5434), .B(n900), .Z(n1950) );
  XOR U5929 ( .A(n5393), .B(n5382), .Z(n5384) );
  XNOR U5930 ( .A(n5374), .B(n5442), .Z(n5382) );
  ANDN U5931 ( .B(n1960), .A(n5393), .Z(n5441) );
  XNOR U5932 ( .A(n893), .B(n5378), .Z(n5393) );
  XOR U5933 ( .A(n5443), .B(n5444), .Z(n5378) );
  XNOR U5934 ( .A(n5445), .B(n5446), .Z(n5444) );
  XOR U5935 ( .A(n5442), .B(n5426), .Z(n5422) );
  IV U5936 ( .A(n900), .Z(n5426) );
  XOR U5937 ( .A(n5447), .B(n5448), .Z(n900) );
  XNOR U5938 ( .A(n5449), .B(n5446), .Z(n5448) );
  IV U5939 ( .A(n1966), .Z(n5442) );
  XOR U5940 ( .A(n5446), .B(n5450), .Z(n1966) );
  XNOR U5941 ( .A(n5451), .B(n5452), .Z(n5435) );
  XNOR U5942 ( .A(n5453), .B(n5433), .Z(n5452) );
  OR U5943 ( .A(n1956), .B(n5373), .Z(n5433) );
  XNOR U5944 ( .A(n893), .B(n5374), .Z(n5373) );
  IV U5945 ( .A(n5451), .Z(n5374) );
  XOR U5946 ( .A(n1945), .B(n5434), .Z(n1956) );
  IV U5947 ( .A(n1953), .Z(n5434) );
  XOR U5948 ( .A(n5430), .B(n5454), .Z(n1953) );
  XNOR U5949 ( .A(n5449), .B(n5443), .Z(n5454) );
  XOR U5950 ( .A(n5455), .B(n5456), .Z(n5443) );
  XNOR U5951 ( .A(n429), .B(n1072), .Z(n5456) );
  XNOR U5952 ( .A(n391), .B(n1071), .Z(n429) );
  XNOR U5953 ( .A(key[1186]), .B(n433), .Z(n5455) );
  IV U5954 ( .A(n4463), .Z(n433) );
  XOR U5955 ( .A(n1033), .B(n1076), .Z(n4463) );
  XOR U5956 ( .A(n5457), .B(n5458), .Z(n1076) );
  XNOR U5957 ( .A(n5459), .B(n5460), .Z(n5457) );
  IV U5958 ( .A(n1506), .Z(n5430) );
  XOR U5959 ( .A(n5447), .B(n5461), .Z(n1506) );
  XOR U5960 ( .A(n5446), .B(n5462), .Z(n5461) );
  NOR U5961 ( .A(n1945), .B(n893), .Z(n5453) );
  XOR U5962 ( .A(n5447), .B(n5463), .Z(n1945) );
  XOR U5963 ( .A(n5446), .B(n5464), .Z(n5463) );
  XOR U5964 ( .A(n5465), .B(n5466), .Z(n5446) );
  XNOR U5965 ( .A(n4433), .B(n1040), .Z(n5466) );
  XNOR U5966 ( .A(n405), .B(n5467), .Z(n1040) );
  XOR U5967 ( .A(n398), .B(n4434), .Z(n405) );
  IV U5968 ( .A(n1046), .Z(n4434) );
  XOR U5969 ( .A(n5468), .B(n5469), .Z(n1046) );
  XNOR U5970 ( .A(n5470), .B(n5471), .Z(n398) );
  XNOR U5971 ( .A(n5472), .B(n1057), .Z(n4433) );
  XOR U5972 ( .A(n5473), .B(n5474), .Z(n1057) );
  XOR U5973 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U5974 ( .A(n5477), .B(n5478), .Z(n5473) );
  XOR U5975 ( .A(n893), .B(n5479), .Z(n5465) );
  XNOR U5976 ( .A(key[1190]), .B(n1050), .Z(n5479) );
  IV U5977 ( .A(n5450), .Z(n5447) );
  XOR U5978 ( .A(n5480), .B(n5481), .Z(n5450) );
  XNOR U5979 ( .A(n4441), .B(n1047), .Z(n5481) );
  XNOR U5980 ( .A(n406), .B(n1063), .Z(n1047) );
  XNOR U5981 ( .A(n5482), .B(n5483), .Z(n1063) );
  XOR U5982 ( .A(n5484), .B(n5485), .Z(n5483) );
  XNOR U5983 ( .A(n5486), .B(n5487), .Z(n5482) );
  XNOR U5984 ( .A(n5488), .B(n5489), .Z(n5487) );
  ANDN U5985 ( .B(n5490), .A(n5491), .Z(n5489) );
  XOR U5986 ( .A(n5492), .B(n5493), .Z(n406) );
  XNOR U5987 ( .A(n5494), .B(n5495), .Z(n5493) );
  XNOR U5988 ( .A(n5496), .B(n5497), .Z(n5492) );
  XOR U5989 ( .A(n5498), .B(n5499), .Z(n5497) );
  ANDN U5990 ( .B(n5500), .A(n5501), .Z(n5499) );
  XNOR U5991 ( .A(key[1189]), .B(n4436), .Z(n5480) );
  XNOR U5992 ( .A(n1042), .B(n1050), .Z(n4436) );
  XNOR U5993 ( .A(n5502), .B(n5503), .Z(n1050) );
  XNOR U5994 ( .A(n5460), .B(n5504), .Z(n1042) );
  XNOR U5995 ( .A(n5505), .B(n5506), .Z(n5460) );
  XNOR U5996 ( .A(n5507), .B(n5508), .Z(n5506) );
  ANDN U5997 ( .B(n5509), .A(n5510), .Z(n5507) );
  XOR U5998 ( .A(n5511), .B(n5512), .Z(n5451) );
  XNOR U5999 ( .A(n5464), .B(n5462), .Z(n5512) );
  XNOR U6000 ( .A(n5513), .B(n5514), .Z(n5462) );
  XOR U6001 ( .A(n5467), .B(n1056), .Z(n5514) );
  XNOR U6002 ( .A(n4438), .B(n1043), .Z(n1056) );
  XNOR U6003 ( .A(n5515), .B(n5516), .Z(n1043) );
  XNOR U6004 ( .A(n5468), .B(n5485), .Z(n5516) );
  XNOR U6005 ( .A(n5517), .B(n5518), .Z(n5485) );
  XNOR U6006 ( .A(n5519), .B(n5520), .Z(n5518) );
  OR U6007 ( .A(n5521), .B(n5522), .Z(n5520) );
  XOR U6008 ( .A(n5523), .B(n5524), .Z(n5515) );
  XOR U6009 ( .A(n5525), .B(n5526), .Z(n4438) );
  XNOR U6010 ( .A(n5470), .B(n5495), .Z(n5526) );
  XNOR U6011 ( .A(n5527), .B(n5528), .Z(n5495) );
  XNOR U6012 ( .A(n5529), .B(n5530), .Z(n5528) );
  OR U6013 ( .A(n5531), .B(n5532), .Z(n5530) );
  XNOR U6014 ( .A(n5533), .B(n4447), .Z(n5467) );
  XNOR U6015 ( .A(n5534), .B(n5535), .Z(n4447) );
  XOR U6016 ( .A(n5536), .B(n5537), .Z(n5535) );
  XOR U6017 ( .A(n5538), .B(n5539), .Z(n5534) );
  XNOR U6018 ( .A(key[1191]), .B(n5472), .Z(n5513) );
  XNOR U6019 ( .A(n5540), .B(n1059), .Z(n5464) );
  XOR U6020 ( .A(n5541), .B(n5542), .Z(n1059) );
  XOR U6021 ( .A(n420), .B(n1077), .Z(n5542) );
  XOR U6022 ( .A(n1071), .B(n5484), .Z(n1077) );
  XOR U6023 ( .A(n5523), .B(n5543), .Z(n1071) );
  XOR U6024 ( .A(n5494), .B(n391), .Z(n420) );
  XNOR U6025 ( .A(n5544), .B(n5545), .Z(n391) );
  XOR U6026 ( .A(n438), .B(n4441), .Z(n5541) );
  XNOR U6027 ( .A(n5546), .B(n5547), .Z(n4441) );
  XNOR U6028 ( .A(n5548), .B(n5537), .Z(n5547) );
  XNOR U6029 ( .A(n5549), .B(n5550), .Z(n5537) );
  XNOR U6030 ( .A(n5551), .B(n5552), .Z(n5550) );
  NANDN U6031 ( .A(n5553), .B(n5554), .Z(n5552) );
  XNOR U6032 ( .A(n5555), .B(n5556), .Z(n5546) );
  XOR U6033 ( .A(n5557), .B(n5558), .Z(n5556) );
  ANDN U6034 ( .B(n5559), .A(n5560), .Z(n5558) );
  XNOR U6035 ( .A(n4451), .B(n5561), .Z(n5540) );
  XOR U6036 ( .A(key[1188]), .B(n4452), .Z(n5561) );
  XNOR U6037 ( .A(n4448), .B(n1048), .Z(n4451) );
  XNOR U6038 ( .A(n5562), .B(n5563), .Z(n1048) );
  XNOR U6039 ( .A(n5564), .B(n5476), .Z(n5563) );
  XNOR U6040 ( .A(n5565), .B(n5566), .Z(n5476) );
  XNOR U6041 ( .A(n5567), .B(n5568), .Z(n5566) );
  NANDN U6042 ( .A(n5569), .B(n5570), .Z(n5568) );
  XNOR U6043 ( .A(n5571), .B(n5572), .Z(n5562) );
  XOR U6044 ( .A(n5508), .B(n5573), .Z(n5572) );
  ANDN U6045 ( .B(n5574), .A(n5575), .Z(n5573) );
  ANDN U6046 ( .B(n5576), .A(n5577), .Z(n5508) );
  XNOR U6047 ( .A(n893), .B(n5445), .Z(n5511) );
  XOR U6048 ( .A(n5578), .B(n5579), .Z(n5445) );
  XNOR U6049 ( .A(n1068), .B(n5580), .Z(n5579) );
  XOR U6050 ( .A(n5449), .B(n4457), .Z(n5580) );
  XNOR U6051 ( .A(n5472), .B(n1061), .Z(n4457) );
  XOR U6052 ( .A(n5571), .B(n1030), .Z(n1061) );
  IV U6053 ( .A(n4448), .Z(n5472) );
  XOR U6054 ( .A(n5571), .B(n5581), .Z(n4448) );
  XNOR U6055 ( .A(n5565), .B(n5582), .Z(n5571) );
  XNOR U6056 ( .A(n5583), .B(n5584), .Z(n5582) );
  ANDN U6057 ( .B(n5585), .A(n5510), .Z(n5583) );
  IV U6058 ( .A(n5586), .Z(n5510) );
  XNOR U6059 ( .A(n5587), .B(n5588), .Z(n5565) );
  XNOR U6060 ( .A(n5589), .B(n5590), .Z(n5588) );
  NANDN U6061 ( .A(n5591), .B(n5592), .Z(n5590) );
  XOR U6062 ( .A(n5593), .B(n5594), .Z(n5449) );
  XNOR U6063 ( .A(n5595), .B(n389), .Z(n5594) );
  XNOR U6064 ( .A(n5596), .B(n1030), .Z(n389) );
  XOR U6065 ( .A(n5581), .B(n5477), .Z(n1030) );
  XNOR U6066 ( .A(key[1185]), .B(n436), .Z(n5593) );
  XNOR U6067 ( .A(n4461), .B(n430), .Z(n436) );
  XOR U6068 ( .A(n5470), .B(n5597), .Z(n430) );
  XOR U6069 ( .A(n5544), .B(n5598), .Z(n5597) );
  XOR U6070 ( .A(n5599), .B(n5600), .Z(n5470) );
  IV U6071 ( .A(n1083), .Z(n4461) );
  XNOR U6072 ( .A(n5468), .B(n5601), .Z(n1083) );
  XOR U6073 ( .A(n5602), .B(n5524), .Z(n5601) );
  XOR U6074 ( .A(n5543), .B(n5603), .Z(n5468) );
  XOR U6075 ( .A(n438), .B(n4452), .Z(n1068) );
  XOR U6076 ( .A(n5555), .B(n5596), .Z(n4452) );
  IV U6077 ( .A(n1072), .Z(n5596) );
  XNOR U6078 ( .A(n5604), .B(n5538), .Z(n1072) );
  XNOR U6079 ( .A(n390), .B(n5605), .Z(n5578) );
  XNOR U6080 ( .A(key[1187]), .B(n1033), .Z(n5605) );
  XOR U6081 ( .A(n5606), .B(n5607), .Z(n1033) );
  XNOR U6082 ( .A(n5608), .B(n5502), .Z(n5606) );
  XNOR U6083 ( .A(n5609), .B(n5610), .Z(n5502) );
  XNOR U6084 ( .A(n5611), .B(n5557), .Z(n5610) );
  ANDN U6085 ( .B(n5612), .A(n5613), .Z(n5557) );
  ANDN U6086 ( .B(n5614), .A(n5615), .Z(n5611) );
  IV U6087 ( .A(n1067), .Z(n390) );
  XNOR U6088 ( .A(n431), .B(n1031), .Z(n1067) );
  XNOR U6089 ( .A(n5616), .B(n5617), .Z(n1031) );
  XOR U6090 ( .A(n5603), .B(n5469), .Z(n5617) );
  XOR U6091 ( .A(n5618), .B(n5619), .Z(n5469) );
  XOR U6092 ( .A(n5620), .B(n5488), .Z(n5619) );
  NANDN U6093 ( .A(n5621), .B(n5622), .Z(n5488) );
  ANDN U6094 ( .B(n5623), .A(n5624), .Z(n5620) );
  XNOR U6095 ( .A(n5486), .B(n5625), .Z(n5603) );
  XNOR U6096 ( .A(n5626), .B(n5627), .Z(n5625) );
  NANDN U6097 ( .A(n5628), .B(n5629), .Z(n5627) );
  XNOR U6098 ( .A(n5602), .B(n5524), .Z(n5616) );
  XOR U6099 ( .A(n5618), .B(n5630), .Z(n5524) );
  XNOR U6100 ( .A(n5626), .B(n5631), .Z(n5630) );
  NANDN U6101 ( .A(n5521), .B(n5632), .Z(n5631) );
  OR U6102 ( .A(n5633), .B(n5634), .Z(n5626) );
  XNOR U6103 ( .A(n5486), .B(n5635), .Z(n5618) );
  XNOR U6104 ( .A(n5636), .B(n5637), .Z(n5635) );
  NAND U6105 ( .A(n5638), .B(n5639), .Z(n5637) );
  XOR U6106 ( .A(n5640), .B(n5636), .Z(n5486) );
  NANDN U6107 ( .A(n5641), .B(n5642), .Z(n5636) );
  ANDN U6108 ( .B(n5643), .A(n5644), .Z(n5640) );
  IV U6109 ( .A(n5523), .Z(n5602) );
  XOR U6110 ( .A(n5645), .B(n5646), .Z(n5523) );
  XNOR U6111 ( .A(n5647), .B(n5648), .Z(n5646) );
  NAND U6112 ( .A(n5649), .B(n5490), .Z(n5648) );
  XOR U6113 ( .A(n5525), .B(n5650), .Z(n431) );
  XNOR U6114 ( .A(n5600), .B(n5471), .Z(n5650) );
  XNOR U6115 ( .A(n5651), .B(n5652), .Z(n5471) );
  XNOR U6116 ( .A(n5653), .B(n5498), .Z(n5652) );
  ANDN U6117 ( .B(n5654), .A(n5655), .Z(n5498) );
  ANDN U6118 ( .B(n5656), .A(n5657), .Z(n5653) );
  XNOR U6119 ( .A(n5496), .B(n5658), .Z(n5600) );
  XNOR U6120 ( .A(n5659), .B(n5660), .Z(n5658) );
  NANDN U6121 ( .A(n5661), .B(n5662), .Z(n5660) );
  XNOR U6122 ( .A(n5544), .B(n5598), .Z(n5525) );
  XOR U6123 ( .A(n5651), .B(n5663), .Z(n5598) );
  XNOR U6124 ( .A(n5659), .B(n5664), .Z(n5663) );
  NANDN U6125 ( .A(n5531), .B(n5665), .Z(n5664) );
  OR U6126 ( .A(n5666), .B(n5667), .Z(n5659) );
  XNOR U6127 ( .A(n5496), .B(n5668), .Z(n5651) );
  XNOR U6128 ( .A(n5669), .B(n5670), .Z(n5668) );
  NAND U6129 ( .A(n5671), .B(n5672), .Z(n5670) );
  XOR U6130 ( .A(n5673), .B(n5669), .Z(n5496) );
  NANDN U6131 ( .A(n5674), .B(n5675), .Z(n5669) );
  ANDN U6132 ( .B(n5676), .A(n5677), .Z(n5673) );
  XNOR U6133 ( .A(n5678), .B(n5679), .Z(n5544) );
  XNOR U6134 ( .A(n5680), .B(n5681), .Z(n5679) );
  NAND U6135 ( .A(n5682), .B(n5500), .Z(n5681) );
  XNOR U6136 ( .A(n5683), .B(n5684), .Z(n893) );
  XNOR U6137 ( .A(n428), .B(n1055), .Z(n5684) );
  XNOR U6138 ( .A(n438), .B(n413), .Z(n1055) );
  IV U6139 ( .A(n1062), .Z(n413) );
  XOR U6140 ( .A(n5543), .B(n5484), .Z(n1062) );
  XOR U6141 ( .A(n5517), .B(n5685), .Z(n5484) );
  XOR U6142 ( .A(n5686), .B(n5647), .Z(n5685) );
  NANDN U6143 ( .A(n5687), .B(n5622), .Z(n5647) );
  XOR U6144 ( .A(n5623), .B(n5490), .Z(n5622) );
  ANDN U6145 ( .B(n5623), .A(n5688), .Z(n5686) );
  XNOR U6146 ( .A(n5645), .B(n5689), .Z(n5517) );
  XNOR U6147 ( .A(n5690), .B(n5691), .Z(n5689) );
  NAND U6148 ( .A(n5639), .B(n5692), .Z(n5691) );
  XOR U6149 ( .A(n5645), .B(n5693), .Z(n5543) );
  XOR U6150 ( .A(n5694), .B(n5519), .Z(n5693) );
  OR U6151 ( .A(n5695), .B(n5633), .Z(n5519) );
  XNOR U6152 ( .A(n5521), .B(n5628), .Z(n5633) );
  NOR U6153 ( .A(n5696), .B(n5628), .Z(n5694) );
  XOR U6154 ( .A(n5697), .B(n5690), .Z(n5645) );
  OR U6155 ( .A(n5641), .B(n5698), .Z(n5690) );
  XNOR U6156 ( .A(n5699), .B(n5639), .Z(n5641) );
  XNOR U6157 ( .A(n5628), .B(n5490), .Z(n5639) );
  XOR U6158 ( .A(n5700), .B(n5701), .Z(n5490) );
  NANDN U6159 ( .A(n5702), .B(n5703), .Z(n5701) );
  XNOR U6160 ( .A(n5704), .B(n5705), .Z(n5628) );
  OR U6161 ( .A(n5702), .B(n5706), .Z(n5705) );
  ANDN U6162 ( .B(n5699), .A(n5707), .Z(n5697) );
  IV U6163 ( .A(n5644), .Z(n5699) );
  XOR U6164 ( .A(n5521), .B(n5623), .Z(n5644) );
  XNOR U6165 ( .A(n5708), .B(n5700), .Z(n5623) );
  NANDN U6166 ( .A(n5709), .B(n5710), .Z(n5700) );
  ANDN U6167 ( .B(n5711), .A(n5712), .Z(n5708) );
  NANDN U6168 ( .A(n5709), .B(n5714), .Z(n5704) );
  XOR U6169 ( .A(n5715), .B(n5702), .Z(n5709) );
  XNOR U6170 ( .A(n5716), .B(n5717), .Z(n5702) );
  XOR U6171 ( .A(n5718), .B(n5711), .Z(n5717) );
  XNOR U6172 ( .A(n5719), .B(n5720), .Z(n5716) );
  XNOR U6173 ( .A(n5721), .B(n5722), .Z(n5720) );
  ANDN U6174 ( .B(n5711), .A(n5723), .Z(n5721) );
  IV U6175 ( .A(n5724), .Z(n5711) );
  ANDN U6176 ( .B(n5715), .A(n5723), .Z(n5713) );
  IV U6177 ( .A(n5719), .Z(n5723) );
  IV U6178 ( .A(n5712), .Z(n5715) );
  XNOR U6179 ( .A(n5718), .B(n5725), .Z(n5712) );
  XOR U6180 ( .A(n5726), .B(n5722), .Z(n5725) );
  NAND U6181 ( .A(n5714), .B(n5710), .Z(n5722) );
  XNOR U6182 ( .A(n5703), .B(n5724), .Z(n5710) );
  XOR U6183 ( .A(n5727), .B(n5728), .Z(n5724) );
  XOR U6184 ( .A(n5729), .B(n5730), .Z(n5728) );
  XNOR U6185 ( .A(n5629), .B(n5731), .Z(n5730) );
  XNOR U6186 ( .A(n5732), .B(n5733), .Z(n5727) );
  XNOR U6187 ( .A(n5734), .B(n5735), .Z(n5733) );
  ANDN U6188 ( .B(n5632), .A(n5522), .Z(n5734) );
  XNOR U6189 ( .A(n5719), .B(n5706), .Z(n5714) );
  XOR U6190 ( .A(n5736), .B(n5737), .Z(n5719) );
  XNOR U6191 ( .A(n5738), .B(n5731), .Z(n5737) );
  XOR U6192 ( .A(n5739), .B(n5740), .Z(n5731) );
  XNOR U6193 ( .A(n5741), .B(n5742), .Z(n5740) );
  NAND U6194 ( .A(n5692), .B(n5638), .Z(n5742) );
  XNOR U6195 ( .A(n5743), .B(n5744), .Z(n5736) );
  ANDN U6196 ( .B(n5745), .A(n5688), .Z(n5743) );
  ANDN U6197 ( .B(n5703), .A(n5706), .Z(n5726) );
  XOR U6198 ( .A(n5706), .B(n5703), .Z(n5718) );
  XNOR U6199 ( .A(n5746), .B(n5747), .Z(n5703) );
  XNOR U6200 ( .A(n5739), .B(n5748), .Z(n5747) );
  XNOR U6201 ( .A(n5738), .B(n5632), .Z(n5748) );
  XNOR U6202 ( .A(n5749), .B(n5750), .Z(n5746) );
  XNOR U6203 ( .A(n5751), .B(n5735), .Z(n5750) );
  OR U6204 ( .A(n5634), .B(n5695), .Z(n5735) );
  XNOR U6205 ( .A(n5749), .B(n5732), .Z(n5695) );
  XNOR U6206 ( .A(n5632), .B(n5629), .Z(n5634) );
  ANDN U6207 ( .B(n5629), .A(n5696), .Z(n5751) );
  XOR U6208 ( .A(n5752), .B(n5753), .Z(n5706) );
  XOR U6209 ( .A(n5739), .B(n5729), .Z(n5753) );
  XOR U6210 ( .A(n5649), .B(n5491), .Z(n5729) );
  XOR U6211 ( .A(n5754), .B(n5741), .Z(n5739) );
  NANDN U6212 ( .A(n5698), .B(n5642), .Z(n5741) );
  XOR U6213 ( .A(n5643), .B(n5638), .Z(n5642) );
  XNOR U6214 ( .A(n5745), .B(n5755), .Z(n5629) );
  XNOR U6215 ( .A(n5756), .B(n5757), .Z(n5755) );
  XOR U6216 ( .A(n5707), .B(n5692), .Z(n5698) );
  XNOR U6217 ( .A(n5696), .B(n5649), .Z(n5692) );
  IV U6218 ( .A(n5732), .Z(n5696) );
  XOR U6219 ( .A(n5758), .B(n5759), .Z(n5732) );
  XOR U6220 ( .A(n5760), .B(n5761), .Z(n5759) );
  XOR U6221 ( .A(n5749), .B(n5762), .Z(n5758) );
  ANDN U6222 ( .B(n5643), .A(n5707), .Z(n5754) );
  XNOR U6223 ( .A(n5749), .B(n5763), .Z(n5707) );
  XOR U6224 ( .A(n5745), .B(n5632), .Z(n5643) );
  XNOR U6225 ( .A(n5764), .B(n5765), .Z(n5632) );
  XOR U6226 ( .A(n5766), .B(n5761), .Z(n5765) );
  XNOR U6227 ( .A(n5767), .B(n5768), .Z(n5761) );
  XOR U6228 ( .A(n5242), .B(n5243), .Z(n5768) );
  XNOR U6229 ( .A(n3904), .B(n5222), .Z(n5243) );
  XNOR U6230 ( .A(n5769), .B(n5770), .Z(n3904) );
  XNOR U6231 ( .A(n5771), .B(n5772), .Z(n5770) );
  XNOR U6232 ( .A(n5773), .B(n5774), .Z(n5769) );
  XOR U6233 ( .A(n5775), .B(n5776), .Z(n5774) );
  ANDN U6234 ( .B(n5777), .A(n5778), .Z(n5776) );
  XNOR U6235 ( .A(key[1044]), .B(n3897), .Z(n5767) );
  XOR U6236 ( .A(n5779), .B(n5780), .Z(n3897) );
  XNOR U6237 ( .A(n3932), .B(n5212), .Z(n5780) );
  IV U6238 ( .A(n2671), .Z(n5212) );
  XOR U6239 ( .A(n5781), .B(n2644), .Z(n2671) );
  XNOR U6240 ( .A(n5782), .B(n3940), .Z(n3932) );
  XNOR U6241 ( .A(n5783), .B(n5226), .Z(n5779) );
  IV U6242 ( .A(n5624), .Z(n5745) );
  XOR U6243 ( .A(n5738), .B(n5784), .Z(n5752) );
  XNOR U6244 ( .A(n5785), .B(n5744), .Z(n5784) );
  OR U6245 ( .A(n5621), .B(n5687), .Z(n5744) );
  XNOR U6246 ( .A(n5763), .B(n5649), .Z(n5687) );
  XNOR U6247 ( .A(n5624), .B(n5491), .Z(n5621) );
  ANDN U6248 ( .B(n5649), .A(n5491), .Z(n5785) );
  XOR U6249 ( .A(n5764), .B(n5786), .Z(n5491) );
  XOR U6250 ( .A(n5756), .B(n5787), .Z(n5786) );
  XOR U6251 ( .A(n5766), .B(n5764), .Z(n5649) );
  XNOR U6252 ( .A(n5688), .B(n5624), .Z(n5738) );
  XOR U6253 ( .A(n5764), .B(n5788), .Z(n5624) );
  XNOR U6254 ( .A(n5766), .B(n5760), .Z(n5788) );
  XOR U6255 ( .A(n5789), .B(n5790), .Z(n5760) );
  XNOR U6256 ( .A(n5791), .B(n3912), .Z(n5790) );
  XOR U6257 ( .A(n3924), .B(n5232), .Z(n3912) );
  XNOR U6258 ( .A(n5792), .B(n5793), .Z(n5232) );
  XOR U6259 ( .A(n5794), .B(n5795), .Z(n5793) );
  XNOR U6260 ( .A(n5796), .B(n5797), .Z(n5792) );
  IV U6261 ( .A(n5220), .Z(n3924) );
  XNOR U6262 ( .A(n5798), .B(n5799), .Z(n5220) );
  XNOR U6263 ( .A(key[1047]), .B(n5238), .Z(n5789) );
  XNOR U6264 ( .A(n5802), .B(n5803), .Z(n5764) );
  XOR U6265 ( .A(n5226), .B(n5231), .Z(n5803) );
  XOR U6266 ( .A(n3907), .B(n3926), .Z(n5231) );
  XOR U6267 ( .A(n5804), .B(n5805), .Z(n3926) );
  IV U6268 ( .A(n5806), .Z(n3907) );
  XNOR U6269 ( .A(n5807), .B(n5808), .Z(n5226) );
  XNOR U6270 ( .A(n5809), .B(n5810), .Z(n5808) );
  XOR U6271 ( .A(n5811), .B(n5812), .Z(n5807) );
  XOR U6272 ( .A(n5813), .B(n5814), .Z(n5812) );
  ANDN U6273 ( .B(n5815), .A(n5816), .Z(n5814) );
  XNOR U6274 ( .A(key[1045]), .B(n3903), .Z(n5802) );
  XNOR U6275 ( .A(n3896), .B(n2659), .Z(n3903) );
  XOR U6276 ( .A(n5817), .B(n5818), .Z(n2659) );
  XOR U6277 ( .A(n5819), .B(n5781), .Z(n5818) );
  XNOR U6278 ( .A(n5796), .B(n5820), .Z(n5817) );
  XOR U6279 ( .A(n5821), .B(n5822), .Z(n5820) );
  ANDN U6280 ( .B(n5823), .A(n5824), .Z(n5822) );
  XNOR U6281 ( .A(n5825), .B(n5826), .Z(n5796) );
  XNOR U6282 ( .A(n5827), .B(n5828), .Z(n5826) );
  NANDN U6283 ( .A(n5829), .B(n5830), .Z(n5828) );
  XOR U6284 ( .A(n5831), .B(n5832), .Z(n3896) );
  XOR U6285 ( .A(n5800), .B(n5782), .Z(n5832) );
  XNOR U6286 ( .A(n5833), .B(n5834), .Z(n5800) );
  XNOR U6287 ( .A(n5835), .B(n5836), .Z(n5834) );
  NANDN U6288 ( .A(n5837), .B(n5838), .Z(n5836) );
  XNOR U6289 ( .A(n5839), .B(n5840), .Z(n5831) );
  XOR U6290 ( .A(n5841), .B(n5842), .Z(n5840) );
  ANDN U6291 ( .B(n5843), .A(n5844), .Z(n5842) );
  IV U6292 ( .A(n5763), .Z(n5688) );
  XNOR U6293 ( .A(n5757), .B(n5845), .Z(n5763) );
  XOR U6294 ( .A(n5762), .B(n5787), .Z(n5845) );
  IV U6295 ( .A(n5766), .Z(n5787) );
  XOR U6296 ( .A(n5846), .B(n5847), .Z(n5766) );
  XOR U6297 ( .A(n5230), .B(n5522), .Z(n5847) );
  IV U6298 ( .A(n5749), .Z(n5522) );
  XOR U6299 ( .A(n5848), .B(n5849), .Z(n5749) );
  XNOR U6300 ( .A(n3910), .B(n2680), .Z(n5849) );
  XNOR U6301 ( .A(n3944), .B(n3937), .Z(n2680) );
  XOR U6302 ( .A(n5850), .B(n5851), .Z(n3937) );
  XOR U6303 ( .A(n5852), .B(n5804), .Z(n5851) );
  XOR U6304 ( .A(n2689), .B(n3923), .Z(n3910) );
  IV U6305 ( .A(n2666), .Z(n3923) );
  XOR U6306 ( .A(n5853), .B(n5782), .Z(n2666) );
  XOR U6307 ( .A(n5833), .B(n5854), .Z(n5782) );
  XOR U6308 ( .A(n5855), .B(n5856), .Z(n5854) );
  ANDN U6309 ( .B(n5857), .A(n5858), .Z(n5855) );
  XNOR U6310 ( .A(n5859), .B(n5860), .Z(n5833) );
  XNOR U6311 ( .A(n5861), .B(n5862), .Z(n5860) );
  NANDN U6312 ( .A(n5863), .B(n5864), .Z(n5862) );
  XOR U6313 ( .A(key[1040]), .B(n5213), .Z(n5848) );
  XNOR U6314 ( .A(n5781), .B(n5865), .Z(n5213) );
  XOR U6315 ( .A(n5825), .B(n5866), .Z(n5781) );
  XOR U6316 ( .A(n5867), .B(n5868), .Z(n5866) );
  NOR U6317 ( .A(n5869), .B(n5870), .Z(n5867) );
  XNOR U6318 ( .A(n5871), .B(n5872), .Z(n5825) );
  XNOR U6319 ( .A(n5873), .B(n5874), .Z(n5872) );
  NANDN U6320 ( .A(n5875), .B(n5876), .Z(n5874) );
  XNOR U6321 ( .A(n5222), .B(n3911), .Z(n5230) );
  XNOR U6322 ( .A(n5877), .B(n5878), .Z(n3911) );
  XNOR U6323 ( .A(n5804), .B(n5850), .Z(n5878) );
  XNOR U6324 ( .A(n5773), .B(n5852), .Z(n5877) );
  XNOR U6325 ( .A(n5881), .B(n5882), .Z(n5773) );
  XNOR U6326 ( .A(n5883), .B(n5884), .Z(n5882) );
  NANDN U6327 ( .A(n5885), .B(n5886), .Z(n5884) );
  IV U6328 ( .A(n5238), .Z(n5222) );
  XNOR U6329 ( .A(n3922), .B(n5887), .Z(n5846) );
  XOR U6330 ( .A(key[1046]), .B(n5806), .Z(n5887) );
  XNOR U6331 ( .A(n5888), .B(n5889), .Z(n5806) );
  XNOR U6332 ( .A(n5791), .B(n2657), .Z(n3922) );
  XOR U6333 ( .A(n3905), .B(n2652), .Z(n2657) );
  IV U6334 ( .A(n5225), .Z(n2652) );
  XNOR U6335 ( .A(n5794), .B(n5890), .Z(n5225) );
  XOR U6336 ( .A(n5801), .B(n5891), .Z(n3905) );
  XOR U6337 ( .A(n2689), .B(n5221), .Z(n5791) );
  XOR U6338 ( .A(n5892), .B(n5893), .Z(n5221) );
  XNOR U6339 ( .A(n5888), .B(n5810), .Z(n5892) );
  XNOR U6340 ( .A(n5894), .B(n5895), .Z(n5810) );
  XNOR U6341 ( .A(n5896), .B(n5897), .Z(n5895) );
  NANDN U6342 ( .A(n5898), .B(n5899), .Z(n5897) );
  IV U6343 ( .A(n5783), .Z(n2689) );
  XOR U6344 ( .A(n5900), .B(n5901), .Z(n5762) );
  XNOR U6345 ( .A(n5756), .B(n5902), .Z(n5901) );
  XNOR U6346 ( .A(n3930), .B(n5211), .Z(n5902) );
  XOR U6347 ( .A(n3895), .B(n5238), .Z(n5211) );
  XOR U6348 ( .A(n5772), .B(n5880), .Z(n5238) );
  XOR U6349 ( .A(n5772), .B(n3919), .Z(n3895) );
  XOR U6350 ( .A(n5881), .B(n5903), .Z(n5772) );
  XOR U6351 ( .A(n5904), .B(n5905), .Z(n5903) );
  NOR U6352 ( .A(n5906), .B(n5907), .Z(n5904) );
  XNOR U6353 ( .A(n5908), .B(n5909), .Z(n5881) );
  XNOR U6354 ( .A(n5910), .B(n5911), .Z(n5909) );
  NANDN U6355 ( .A(n5912), .B(n5913), .Z(n5911) );
  XOR U6356 ( .A(n5783), .B(n5242), .Z(n3930) );
  XNOR U6357 ( .A(n5809), .B(n3938), .Z(n5242) );
  XNOR U6358 ( .A(n5894), .B(n5914), .Z(n5809) );
  XOR U6359 ( .A(n5915), .B(n5916), .Z(n5914) );
  ANDN U6360 ( .B(n5917), .A(n5918), .Z(n5915) );
  XNOR U6361 ( .A(n5919), .B(n5920), .Z(n5894) );
  XNOR U6362 ( .A(n5921), .B(n5922), .Z(n5920) );
  NANDN U6363 ( .A(n5923), .B(n5924), .Z(n5922) );
  XOR U6364 ( .A(n5926), .B(n5927), .Z(n5756) );
  XNOR U6365 ( .A(n2688), .B(n5201), .Z(n5927) );
  XNOR U6366 ( .A(n3919), .B(n3938), .Z(n5201) );
  XNOR U6367 ( .A(n5852), .B(n5880), .Z(n3919) );
  XNOR U6368 ( .A(n5908), .B(n5928), .Z(n5880) );
  XOR U6369 ( .A(n5929), .B(n5883), .Z(n5928) );
  OR U6370 ( .A(n5930), .B(n5931), .Z(n5883) );
  ANDN U6371 ( .B(n5932), .A(n5933), .Z(n5929) );
  XOR U6372 ( .A(n3943), .B(n2679), .Z(n2688) );
  IV U6373 ( .A(n5236), .Z(n2679) );
  XNOR U6374 ( .A(n5795), .B(n5934), .Z(n5236) );
  XNOR U6375 ( .A(n5797), .B(n5794), .Z(n5934) );
  XNOR U6376 ( .A(n5936), .B(n5937), .Z(n3943) );
  XNOR U6377 ( .A(n5801), .B(n5938), .Z(n5937) );
  XOR U6378 ( .A(n5853), .B(n5939), .Z(n5801) );
  XNOR U6379 ( .A(key[1041]), .B(n3944), .Z(n5926) );
  XNOR U6380 ( .A(n5940), .B(n5941), .Z(n3944) );
  XNOR U6381 ( .A(n5888), .B(n5942), .Z(n5941) );
  XOR U6382 ( .A(n5925), .B(n5943), .Z(n5888) );
  XNOR U6383 ( .A(n3933), .B(n5944), .Z(n5900) );
  XNOR U6384 ( .A(key[1043]), .B(n3916), .Z(n5944) );
  IV U6385 ( .A(n2642), .Z(n3933) );
  XOR U6386 ( .A(n3917), .B(n2684), .Z(n2642) );
  XOR U6387 ( .A(n5945), .B(n5946), .Z(n2684) );
  XOR U6388 ( .A(n5890), .B(n5795), .Z(n5946) );
  XNOR U6389 ( .A(n5947), .B(n5948), .Z(n5795) );
  XNOR U6390 ( .A(n5949), .B(n5950), .Z(n5948) );
  NANDN U6391 ( .A(n5951), .B(n5830), .Z(n5950) );
  XOR U6392 ( .A(n5947), .B(n5952), .Z(n5890) );
  XNOR U6393 ( .A(n5953), .B(n5821), .Z(n5952) );
  ANDN U6394 ( .B(n5954), .A(n5955), .Z(n5821) );
  NOR U6395 ( .A(n5956), .B(n5870), .Z(n5953) );
  XNOR U6396 ( .A(n5819), .B(n5957), .Z(n5947) );
  XNOR U6397 ( .A(n5958), .B(n5959), .Z(n5957) );
  NANDN U6398 ( .A(n5875), .B(n5960), .Z(n5959) );
  XOR U6399 ( .A(n5797), .B(n5935), .Z(n5945) );
  XOR U6400 ( .A(n5819), .B(n5961), .Z(n5935) );
  XNOR U6401 ( .A(n5949), .B(n5962), .Z(n5961) );
  NANDN U6402 ( .A(n5963), .B(n5964), .Z(n5962) );
  OR U6403 ( .A(n5965), .B(n5966), .Z(n5949) );
  XOR U6404 ( .A(n5967), .B(n5958), .Z(n5819) );
  NANDN U6405 ( .A(n5968), .B(n5969), .Z(n5958) );
  ANDN U6406 ( .B(n5970), .A(n5971), .Z(n5967) );
  XOR U6407 ( .A(n5972), .B(n5799), .Z(n3917) );
  XNOR U6408 ( .A(n5938), .B(n5936), .Z(n5799) );
  XNOR U6409 ( .A(n5973), .B(n5974), .Z(n5936) );
  XNOR U6410 ( .A(n5975), .B(n5976), .Z(n5974) );
  NANDN U6411 ( .A(n5977), .B(n5838), .Z(n5976) );
  XOR U6412 ( .A(n5939), .B(n5891), .Z(n5972) );
  XOR U6413 ( .A(n5973), .B(n5978), .Z(n5891) );
  XNOR U6414 ( .A(n5979), .B(n5841), .Z(n5978) );
  ANDN U6415 ( .B(n5980), .A(n5981), .Z(n5841) );
  ANDN U6416 ( .B(n5857), .A(n5982), .Z(n5979) );
  XNOR U6417 ( .A(n5839), .B(n5983), .Z(n5973) );
  XNOR U6418 ( .A(n5984), .B(n5985), .Z(n5983) );
  NANDN U6419 ( .A(n5863), .B(n5986), .Z(n5985) );
  XOR U6420 ( .A(n5839), .B(n5987), .Z(n5939) );
  XNOR U6421 ( .A(n5975), .B(n5988), .Z(n5987) );
  NANDN U6422 ( .A(n5989), .B(n5990), .Z(n5988) );
  OR U6423 ( .A(n5991), .B(n5992), .Z(n5975) );
  XOR U6424 ( .A(n5993), .B(n5984), .Z(n5839) );
  NANDN U6425 ( .A(n5994), .B(n5995), .Z(n5984) );
  ANDN U6426 ( .B(n5996), .A(n5997), .Z(n5993) );
  XOR U6427 ( .A(n5998), .B(n5999), .Z(n5757) );
  XNOR U6428 ( .A(n3938), .B(n2675), .Z(n5999) );
  XNOR U6429 ( .A(n3916), .B(n3931), .Z(n2675) );
  XNOR U6430 ( .A(n6000), .B(n6001), .Z(n3931) );
  XNOR U6431 ( .A(n5805), .B(n5850), .Z(n6001) );
  XNOR U6432 ( .A(n6002), .B(n6003), .Z(n5850) );
  XNOR U6433 ( .A(n6004), .B(n6005), .Z(n6003) );
  NANDN U6434 ( .A(n6006), .B(n5886), .Z(n6005) );
  XNOR U6435 ( .A(n6002), .B(n6007), .Z(n5805) );
  XNOR U6436 ( .A(n6008), .B(n5775), .Z(n6007) );
  ANDN U6437 ( .B(n6009), .A(n6010), .Z(n5775) );
  NOR U6438 ( .A(n6011), .B(n5907), .Z(n6008) );
  XNOR U6439 ( .A(n6012), .B(n6013), .Z(n6002) );
  XNOR U6440 ( .A(n6014), .B(n6015), .Z(n6013) );
  NANDN U6441 ( .A(n5912), .B(n6016), .Z(n6015) );
  XNOR U6442 ( .A(n5852), .B(n5879), .Z(n6000) );
  XNOR U6443 ( .A(n6012), .B(n6017), .Z(n5879) );
  XNOR U6444 ( .A(n6004), .B(n6018), .Z(n6017) );
  NANDN U6445 ( .A(n6019), .B(n5932), .Z(n6018) );
  OR U6446 ( .A(n5930), .B(n6020), .Z(n6004) );
  XNOR U6447 ( .A(n5886), .B(n5932), .Z(n5930) );
  IV U6448 ( .A(n5771), .Z(n6012) );
  XNOR U6449 ( .A(n6021), .B(n6014), .Z(n5771) );
  NANDN U6450 ( .A(n6022), .B(n6023), .Z(n6014) );
  ANDN U6451 ( .B(n6024), .A(n6025), .Z(n6021) );
  XOR U6452 ( .A(n5908), .B(n6026), .Z(n5852) );
  XNOR U6453 ( .A(n5905), .B(n6027), .Z(n6026) );
  NANDN U6454 ( .A(n6028), .B(n5777), .Z(n6027) );
  XNOR U6455 ( .A(n5907), .B(n5777), .Z(n6009) );
  XOR U6456 ( .A(n6030), .B(n5910), .Z(n5908) );
  OR U6457 ( .A(n6022), .B(n6031), .Z(n5910) );
  XOR U6458 ( .A(n6032), .B(n5912), .Z(n6022) );
  XNOR U6459 ( .A(n5932), .B(n5777), .Z(n5912) );
  XOR U6460 ( .A(n6033), .B(n6034), .Z(n5777) );
  NANDN U6461 ( .A(n6035), .B(n6036), .Z(n6034) );
  XOR U6462 ( .A(n6037), .B(n6038), .Z(n5932) );
  NANDN U6463 ( .A(n6035), .B(n6039), .Z(n6038) );
  ANDN U6464 ( .B(n6032), .A(n6040), .Z(n6030) );
  IV U6465 ( .A(n6025), .Z(n6032) );
  XOR U6466 ( .A(n5907), .B(n5886), .Z(n6025) );
  XNOR U6467 ( .A(n6041), .B(n6037), .Z(n5886) );
  NANDN U6468 ( .A(n6042), .B(n6043), .Z(n6037) );
  XOR U6469 ( .A(n6039), .B(n6044), .Z(n6043) );
  ANDN U6470 ( .B(n6044), .A(n6045), .Z(n6041) );
  XOR U6471 ( .A(n6046), .B(n6033), .Z(n5907) );
  NANDN U6472 ( .A(n6042), .B(n6047), .Z(n6033) );
  XOR U6473 ( .A(n6048), .B(n6036), .Z(n6047) );
  XNOR U6474 ( .A(n6049), .B(n6050), .Z(n6035) );
  XOR U6475 ( .A(n6051), .B(n6052), .Z(n6050) );
  XNOR U6476 ( .A(n6053), .B(n6054), .Z(n6049) );
  XNOR U6477 ( .A(n6055), .B(n6056), .Z(n6054) );
  ANDN U6478 ( .B(n6048), .A(n6052), .Z(n6055) );
  ANDN U6479 ( .B(n6048), .A(n6045), .Z(n6046) );
  XNOR U6480 ( .A(n6051), .B(n6057), .Z(n6045) );
  XOR U6481 ( .A(n6058), .B(n6056), .Z(n6057) );
  NAND U6482 ( .A(n6059), .B(n6060), .Z(n6056) );
  XNOR U6483 ( .A(n6053), .B(n6036), .Z(n6060) );
  IV U6484 ( .A(n6048), .Z(n6053) );
  XNOR U6485 ( .A(n6039), .B(n6052), .Z(n6059) );
  IV U6486 ( .A(n6044), .Z(n6052) );
  XOR U6487 ( .A(n6061), .B(n6062), .Z(n6044) );
  XNOR U6488 ( .A(n6063), .B(n6064), .Z(n6062) );
  XNOR U6489 ( .A(n6065), .B(n6066), .Z(n6061) );
  NOR U6490 ( .A(n6011), .B(n5906), .Z(n6065) );
  AND U6491 ( .A(n6036), .B(n6039), .Z(n6058) );
  XNOR U6492 ( .A(n6036), .B(n6039), .Z(n6051) );
  XNOR U6493 ( .A(n6067), .B(n6068), .Z(n6039) );
  XNOR U6494 ( .A(n6069), .B(n6064), .Z(n6068) );
  XOR U6495 ( .A(n6070), .B(n6071), .Z(n6067) );
  XNOR U6496 ( .A(n6072), .B(n6066), .Z(n6071) );
  OR U6497 ( .A(n6010), .B(n6029), .Z(n6066) );
  XNOR U6498 ( .A(n5906), .B(n6028), .Z(n6029) );
  XNOR U6499 ( .A(n6011), .B(n5778), .Z(n6010) );
  ANDN U6500 ( .B(n6073), .A(n6028), .Z(n6072) );
  XNOR U6501 ( .A(n6074), .B(n6075), .Z(n6036) );
  XNOR U6502 ( .A(n6064), .B(n6076), .Z(n6075) );
  XOR U6503 ( .A(n6006), .B(n6070), .Z(n6076) );
  XNOR U6504 ( .A(n5906), .B(n6077), .Z(n6064) );
  XOR U6505 ( .A(n5885), .B(n6078), .Z(n6074) );
  XNOR U6506 ( .A(n6079), .B(n6080), .Z(n6078) );
  ANDN U6507 ( .B(n6081), .A(n5933), .Z(n6079) );
  XNOR U6508 ( .A(n6082), .B(n6083), .Z(n6048) );
  XNOR U6509 ( .A(n6069), .B(n6084), .Z(n6083) );
  XNOR U6510 ( .A(n6019), .B(n6063), .Z(n6084) );
  XOR U6511 ( .A(n6070), .B(n6085), .Z(n6063) );
  XNOR U6512 ( .A(n6086), .B(n6087), .Z(n6085) );
  NAND U6513 ( .A(n5913), .B(n6016), .Z(n6087) );
  XNOR U6514 ( .A(n6088), .B(n6086), .Z(n6070) );
  NANDN U6515 ( .A(n6031), .B(n6023), .Z(n6086) );
  XOR U6516 ( .A(n6024), .B(n6016), .Z(n6023) );
  XNOR U6517 ( .A(n6081), .B(n5778), .Z(n6016) );
  XOR U6518 ( .A(n6040), .B(n5913), .Z(n6031) );
  XNOR U6519 ( .A(n5933), .B(n6089), .Z(n5913) );
  ANDN U6520 ( .B(n6024), .A(n6040), .Z(n6088) );
  XNOR U6521 ( .A(n5885), .B(n5906), .Z(n6040) );
  XOR U6522 ( .A(n6090), .B(n6091), .Z(n5906) );
  XNOR U6523 ( .A(n6092), .B(n6093), .Z(n6091) );
  XOR U6524 ( .A(n6089), .B(n6073), .Z(n6069) );
  IV U6525 ( .A(n5778), .Z(n6073) );
  XOR U6526 ( .A(n6094), .B(n6095), .Z(n5778) );
  XOR U6527 ( .A(n6096), .B(n6093), .Z(n6095) );
  IV U6528 ( .A(n6028), .Z(n6089) );
  XOR U6529 ( .A(n6093), .B(n6097), .Z(n6028) );
  XNOR U6530 ( .A(n6098), .B(n6099), .Z(n6082) );
  XNOR U6531 ( .A(n6100), .B(n6080), .Z(n6099) );
  OR U6532 ( .A(n6020), .B(n5931), .Z(n6080) );
  XNOR U6533 ( .A(n5885), .B(n5933), .Z(n5931) );
  IV U6534 ( .A(n6098), .Z(n5933) );
  XOR U6535 ( .A(n6006), .B(n6081), .Z(n6020) );
  IV U6536 ( .A(n6019), .Z(n6081) );
  XOR U6537 ( .A(n6077), .B(n6101), .Z(n6019) );
  XNOR U6538 ( .A(n6102), .B(n6090), .Z(n6101) );
  XOR U6539 ( .A(n6103), .B(n6104), .Z(n6090) );
  XNOR U6540 ( .A(n6105), .B(n6106), .Z(n6104) );
  XNOR U6541 ( .A(key[1010]), .B(n6107), .Z(n6103) );
  IV U6542 ( .A(n6011), .Z(n6077) );
  XOR U6543 ( .A(n6094), .B(n6108), .Z(n6011) );
  XOR U6544 ( .A(n6093), .B(n6109), .Z(n6108) );
  NOR U6545 ( .A(n6006), .B(n5885), .Z(n6100) );
  XOR U6546 ( .A(n6094), .B(n6110), .Z(n6006) );
  XOR U6547 ( .A(n6093), .B(n6111), .Z(n6110) );
  XOR U6548 ( .A(n6112), .B(n6113), .Z(n6093) );
  XNOR U6549 ( .A(n5885), .B(n6114), .Z(n6113) );
  XNOR U6550 ( .A(n6115), .B(n6116), .Z(n6112) );
  XNOR U6551 ( .A(key[1014]), .B(n6117), .Z(n6116) );
  IV U6552 ( .A(n6097), .Z(n6094) );
  XOR U6553 ( .A(n6118), .B(n6119), .Z(n6097) );
  XNOR U6554 ( .A(n6120), .B(n6121), .Z(n6119) );
  XNOR U6555 ( .A(key[1013]), .B(n6122), .Z(n6118) );
  XOR U6556 ( .A(n6123), .B(n6124), .Z(n6098) );
  XNOR U6557 ( .A(n6111), .B(n6109), .Z(n6124) );
  XNOR U6558 ( .A(n6125), .B(n6126), .Z(n6109) );
  XNOR U6559 ( .A(n6127), .B(n6128), .Z(n6126) );
  XNOR U6560 ( .A(key[1015]), .B(n6129), .Z(n6125) );
  XNOR U6561 ( .A(n6130), .B(n6131), .Z(n6111) );
  XNOR U6562 ( .A(n6132), .B(n6133), .Z(n6130) );
  XNOR U6563 ( .A(key[1012]), .B(n6134), .Z(n6133) );
  XNOR U6564 ( .A(n5885), .B(n6092), .Z(n6123) );
  XOR U6565 ( .A(n6135), .B(n6136), .Z(n6092) );
  XNOR U6566 ( .A(n6137), .B(n6138), .Z(n6136) );
  XNOR U6567 ( .A(n6139), .B(n6102), .Z(n6138) );
  IV U6568 ( .A(n6096), .Z(n6102) );
  XNOR U6569 ( .A(n6140), .B(n6141), .Z(n6096) );
  XOR U6570 ( .A(n6142), .B(n6143), .Z(n6141) );
  XOR U6571 ( .A(key[1009]), .B(n6144), .Z(n6140) );
  XOR U6572 ( .A(n6145), .B(n6146), .Z(n6135) );
  XNOR U6573 ( .A(key[1011]), .B(n6147), .Z(n6146) );
  XNOR U6574 ( .A(n6148), .B(n6149), .Z(n5885) );
  XNOR U6575 ( .A(n6150), .B(n6151), .Z(n6149) );
  XNOR U6576 ( .A(key[1008]), .B(n6152), .Z(n6148) );
  XOR U6577 ( .A(n6153), .B(n5893), .Z(n3916) );
  XOR U6578 ( .A(n5942), .B(n5940), .Z(n5893) );
  XOR U6579 ( .A(n6154), .B(n6155), .Z(n5940) );
  XNOR U6580 ( .A(n6156), .B(n6157), .Z(n6155) );
  NANDN U6581 ( .A(n6158), .B(n5899), .Z(n6157) );
  XOR U6582 ( .A(n5943), .B(n5889), .Z(n6153) );
  XOR U6583 ( .A(n6154), .B(n6159), .Z(n5889) );
  XNOR U6584 ( .A(n6160), .B(n5813), .Z(n6159) );
  ANDN U6585 ( .B(n6161), .A(n6162), .Z(n5813) );
  ANDN U6586 ( .B(n6163), .A(n5918), .Z(n6160) );
  IV U6587 ( .A(n6164), .Z(n5918) );
  XNOR U6588 ( .A(n5811), .B(n6165), .Z(n6154) );
  XNOR U6589 ( .A(n6166), .B(n6167), .Z(n6165) );
  NANDN U6590 ( .A(n5923), .B(n6168), .Z(n6167) );
  XNOR U6591 ( .A(n6156), .B(n6170), .Z(n6169) );
  NANDN U6592 ( .A(n6171), .B(n6172), .Z(n6170) );
  OR U6593 ( .A(n6173), .B(n6174), .Z(n6156) );
  XNOR U6594 ( .A(n6175), .B(n6166), .Z(n5811) );
  NANDN U6595 ( .A(n6176), .B(n6177), .Z(n6166) );
  ANDN U6596 ( .B(n6178), .A(n6179), .Z(n6175) );
  XNOR U6597 ( .A(n5925), .B(n5942), .Z(n3938) );
  XOR U6598 ( .A(n5919), .B(n6180), .Z(n5942) );
  XNOR U6599 ( .A(n5916), .B(n6181), .Z(n6180) );
  NANDN U6600 ( .A(n6182), .B(n5815), .Z(n6181) );
  XOR U6601 ( .A(n6164), .B(n5815), .Z(n6161) );
  XNOR U6602 ( .A(n5919), .B(n6184), .Z(n5925) );
  XOR U6603 ( .A(n6185), .B(n5896), .Z(n6184) );
  OR U6604 ( .A(n6186), .B(n6173), .Z(n5896) );
  XNOR U6605 ( .A(n5899), .B(n6172), .Z(n6173) );
  ANDN U6606 ( .B(n6172), .A(n6187), .Z(n6185) );
  XOR U6607 ( .A(n6188), .B(n5921), .Z(n5919) );
  OR U6608 ( .A(n6176), .B(n6189), .Z(n5921) );
  XNOR U6609 ( .A(n6179), .B(n5923), .Z(n6176) );
  XNOR U6610 ( .A(n6172), .B(n5815), .Z(n5923) );
  XOR U6611 ( .A(n6190), .B(n6191), .Z(n5815) );
  NANDN U6612 ( .A(n6192), .B(n6193), .Z(n6191) );
  XOR U6613 ( .A(n6194), .B(n6195), .Z(n6172) );
  NANDN U6614 ( .A(n6192), .B(n6196), .Z(n6195) );
  NOR U6615 ( .A(n6179), .B(n6197), .Z(n6188) );
  XNOR U6616 ( .A(n6164), .B(n5899), .Z(n6179) );
  XNOR U6617 ( .A(n6198), .B(n6194), .Z(n5899) );
  NANDN U6618 ( .A(n6199), .B(n6200), .Z(n6194) );
  XOR U6619 ( .A(n6196), .B(n6201), .Z(n6200) );
  ANDN U6620 ( .B(n6201), .A(n6202), .Z(n6198) );
  XNOR U6621 ( .A(n6203), .B(n6190), .Z(n6164) );
  NANDN U6622 ( .A(n6199), .B(n6204), .Z(n6190) );
  XOR U6623 ( .A(n6205), .B(n6193), .Z(n6204) );
  XNOR U6624 ( .A(n6206), .B(n6207), .Z(n6192) );
  XOR U6625 ( .A(n6208), .B(n6209), .Z(n6207) );
  XNOR U6626 ( .A(n6210), .B(n6211), .Z(n6206) );
  XNOR U6627 ( .A(n6212), .B(n6213), .Z(n6211) );
  ANDN U6628 ( .B(n6205), .A(n6209), .Z(n6212) );
  ANDN U6629 ( .B(n6205), .A(n6202), .Z(n6203) );
  XNOR U6630 ( .A(n6208), .B(n6214), .Z(n6202) );
  XOR U6631 ( .A(n6215), .B(n6213), .Z(n6214) );
  NAND U6632 ( .A(n6216), .B(n6217), .Z(n6213) );
  XNOR U6633 ( .A(n6210), .B(n6193), .Z(n6217) );
  IV U6634 ( .A(n6205), .Z(n6210) );
  XNOR U6635 ( .A(n6196), .B(n6209), .Z(n6216) );
  IV U6636 ( .A(n6201), .Z(n6209) );
  XOR U6637 ( .A(n6218), .B(n6219), .Z(n6201) );
  XNOR U6638 ( .A(n6220), .B(n6221), .Z(n6219) );
  XNOR U6639 ( .A(n6222), .B(n6223), .Z(n6218) );
  ANDN U6640 ( .B(n5917), .A(n6224), .Z(n6222) );
  AND U6641 ( .A(n6193), .B(n6196), .Z(n6215) );
  XNOR U6642 ( .A(n6193), .B(n6196), .Z(n6208) );
  XNOR U6643 ( .A(n6225), .B(n6226), .Z(n6196) );
  XNOR U6644 ( .A(n6227), .B(n6221), .Z(n6226) );
  XOR U6645 ( .A(n6228), .B(n6229), .Z(n6225) );
  XNOR U6646 ( .A(n6230), .B(n6223), .Z(n6229) );
  OR U6647 ( .A(n6162), .B(n6183), .Z(n6223) );
  XNOR U6648 ( .A(n5917), .B(n6231), .Z(n6183) );
  XNOR U6649 ( .A(n6224), .B(n5816), .Z(n6162) );
  ANDN U6650 ( .B(n6232), .A(n6182), .Z(n6230) );
  XNOR U6651 ( .A(n6233), .B(n6234), .Z(n6193) );
  XNOR U6652 ( .A(n6221), .B(n6235), .Z(n6234) );
  XOR U6653 ( .A(n6158), .B(n6228), .Z(n6235) );
  XNOR U6654 ( .A(n5917), .B(n6224), .Z(n6221) );
  XOR U6655 ( .A(n5898), .B(n6236), .Z(n6233) );
  XNOR U6656 ( .A(n6237), .B(n6238), .Z(n6236) );
  ANDN U6657 ( .B(n6239), .A(n6187), .Z(n6237) );
  XNOR U6658 ( .A(n6240), .B(n6241), .Z(n6205) );
  XNOR U6659 ( .A(n6227), .B(n6242), .Z(n6241) );
  XNOR U6660 ( .A(n6171), .B(n6220), .Z(n6242) );
  XOR U6661 ( .A(n6228), .B(n6243), .Z(n6220) );
  XNOR U6662 ( .A(n6244), .B(n6245), .Z(n6243) );
  NAND U6663 ( .A(n5924), .B(n6168), .Z(n6245) );
  XNOR U6664 ( .A(n6246), .B(n6244), .Z(n6228) );
  NANDN U6665 ( .A(n6189), .B(n6177), .Z(n6244) );
  XOR U6666 ( .A(n6178), .B(n6168), .Z(n6177) );
  XNOR U6667 ( .A(n6239), .B(n5816), .Z(n6168) );
  XOR U6668 ( .A(n6197), .B(n5924), .Z(n6189) );
  XNOR U6669 ( .A(n6187), .B(n6231), .Z(n5924) );
  ANDN U6670 ( .B(n6178), .A(n6197), .Z(n6246) );
  XOR U6671 ( .A(n5898), .B(n5917), .Z(n6197) );
  XNOR U6672 ( .A(n6247), .B(n6248), .Z(n5917) );
  XNOR U6673 ( .A(n6249), .B(n6250), .Z(n6248) );
  XOR U6674 ( .A(n6231), .B(n6232), .Z(n6227) );
  IV U6675 ( .A(n5816), .Z(n6232) );
  XOR U6676 ( .A(n6251), .B(n6252), .Z(n5816) );
  XOR U6677 ( .A(n6253), .B(n6250), .Z(n6252) );
  IV U6678 ( .A(n6182), .Z(n6231) );
  XOR U6679 ( .A(n6250), .B(n6254), .Z(n6182) );
  XNOR U6680 ( .A(n6255), .B(n6256), .Z(n6240) );
  XNOR U6681 ( .A(n6257), .B(n6238), .Z(n6256) );
  OR U6682 ( .A(n6174), .B(n6186), .Z(n6238) );
  XNOR U6683 ( .A(n5898), .B(n6187), .Z(n6186) );
  IV U6684 ( .A(n6255), .Z(n6187) );
  XOR U6685 ( .A(n6158), .B(n6239), .Z(n6174) );
  IV U6686 ( .A(n6171), .Z(n6239) );
  XOR U6687 ( .A(n6163), .B(n6258), .Z(n6171) );
  XNOR U6688 ( .A(n6259), .B(n6247), .Z(n6258) );
  XOR U6689 ( .A(n6260), .B(n6261), .Z(n6247) );
  XOR U6690 ( .A(n6262), .B(n6263), .Z(n6261) );
  XOR U6691 ( .A(n6264), .B(n6265), .Z(n6260) );
  XNOR U6692 ( .A(key[970]), .B(n6266), .Z(n6265) );
  IV U6693 ( .A(n6224), .Z(n6163) );
  XOR U6694 ( .A(n6251), .B(n6267), .Z(n6224) );
  XOR U6695 ( .A(n6250), .B(n6268), .Z(n6267) );
  NOR U6696 ( .A(n6158), .B(n5898), .Z(n6257) );
  XOR U6697 ( .A(n6251), .B(n6269), .Z(n6158) );
  XOR U6698 ( .A(n6250), .B(n6270), .Z(n6269) );
  XOR U6699 ( .A(n6271), .B(n6272), .Z(n6250) );
  XOR U6700 ( .A(n5898), .B(n6273), .Z(n6272) );
  XNOR U6701 ( .A(n6274), .B(n6275), .Z(n6271) );
  XOR U6702 ( .A(key[974]), .B(n6276), .Z(n6275) );
  IV U6703 ( .A(n6254), .Z(n6251) );
  XOR U6704 ( .A(n6277), .B(n6278), .Z(n6254) );
  XNOR U6705 ( .A(n6279), .B(n6280), .Z(n6278) );
  XNOR U6706 ( .A(n6281), .B(n6282), .Z(n6277) );
  XOR U6707 ( .A(key[973]), .B(n6283), .Z(n6282) );
  XOR U6708 ( .A(n6284), .B(n6285), .Z(n6255) );
  XNOR U6709 ( .A(n6270), .B(n6268), .Z(n6285) );
  XNOR U6710 ( .A(n6286), .B(n6287), .Z(n6268) );
  XOR U6711 ( .A(n6288), .B(n6289), .Z(n6287) );
  XOR U6712 ( .A(key[975]), .B(n6290), .Z(n6286) );
  XNOR U6713 ( .A(n6291), .B(n6292), .Z(n6270) );
  XNOR U6714 ( .A(n6293), .B(n6294), .Z(n6292) );
  XNOR U6715 ( .A(n6295), .B(n6296), .Z(n6291) );
  XNOR U6716 ( .A(key[972]), .B(n6297), .Z(n6296) );
  XNOR U6717 ( .A(n5898), .B(n6249), .Z(n6284) );
  XOR U6718 ( .A(n6298), .B(n6299), .Z(n6249) );
  XNOR U6719 ( .A(n6300), .B(n6301), .Z(n6299) );
  XNOR U6720 ( .A(n6302), .B(n6259), .Z(n6301) );
  IV U6721 ( .A(n6253), .Z(n6259) );
  XNOR U6722 ( .A(n6303), .B(n6304), .Z(n6253) );
  XNOR U6723 ( .A(n6305), .B(n6306), .Z(n6304) );
  XOR U6724 ( .A(n6307), .B(n6308), .Z(n6303) );
  XNOR U6725 ( .A(key[969]), .B(n6309), .Z(n6308) );
  XNOR U6726 ( .A(n6310), .B(n6311), .Z(n6298) );
  XNOR U6727 ( .A(key[971]), .B(n6312), .Z(n6311) );
  XNOR U6728 ( .A(n6313), .B(n6314), .Z(n5898) );
  XNOR U6729 ( .A(n6315), .B(n6316), .Z(n6314) );
  XOR U6730 ( .A(n6317), .B(n6318), .Z(n6313) );
  XNOR U6731 ( .A(key[968]), .B(n6319), .Z(n6318) );
  XOR U6732 ( .A(key[1042]), .B(n2681), .Z(n5998) );
  XOR U6733 ( .A(n3940), .B(n2644), .Z(n2681) );
  XNOR U6734 ( .A(n5797), .B(n5865), .Z(n2644) );
  XNOR U6735 ( .A(n5871), .B(n6320), .Z(n5865) );
  XOR U6736 ( .A(n6321), .B(n5827), .Z(n6320) );
  OR U6737 ( .A(n5965), .B(n6322), .Z(n5827) );
  XNOR U6738 ( .A(n5830), .B(n5964), .Z(n5965) );
  ANDN U6739 ( .B(n5964), .A(n6323), .Z(n6321) );
  XOR U6740 ( .A(n5871), .B(n6324), .Z(n5797) );
  XNOR U6741 ( .A(n5868), .B(n6325), .Z(n6324) );
  NANDN U6742 ( .A(n6326), .B(n5823), .Z(n6325) );
  XNOR U6743 ( .A(n5870), .B(n5823), .Z(n5954) );
  XOR U6744 ( .A(n6328), .B(n5873), .Z(n5871) );
  OR U6745 ( .A(n5968), .B(n6329), .Z(n5873) );
  XOR U6746 ( .A(n6330), .B(n5875), .Z(n5968) );
  XNOR U6747 ( .A(n5964), .B(n5823), .Z(n5875) );
  XOR U6748 ( .A(n6331), .B(n6332), .Z(n5823) );
  NANDN U6749 ( .A(n6333), .B(n6334), .Z(n6332) );
  XOR U6750 ( .A(n6335), .B(n6336), .Z(n5964) );
  NANDN U6751 ( .A(n6333), .B(n6337), .Z(n6336) );
  ANDN U6752 ( .B(n6330), .A(n6338), .Z(n6328) );
  IV U6753 ( .A(n5971), .Z(n6330) );
  XOR U6754 ( .A(n5870), .B(n5830), .Z(n5971) );
  XNOR U6755 ( .A(n6339), .B(n6335), .Z(n5830) );
  NANDN U6756 ( .A(n6340), .B(n6341), .Z(n6335) );
  XOR U6757 ( .A(n6337), .B(n6342), .Z(n6341) );
  ANDN U6758 ( .B(n6342), .A(n6343), .Z(n6339) );
  XOR U6759 ( .A(n6344), .B(n6331), .Z(n5870) );
  NANDN U6760 ( .A(n6340), .B(n6345), .Z(n6331) );
  XOR U6761 ( .A(n6346), .B(n6334), .Z(n6345) );
  XNOR U6762 ( .A(n6347), .B(n6348), .Z(n6333) );
  XOR U6763 ( .A(n6349), .B(n6350), .Z(n6348) );
  XNOR U6764 ( .A(n6351), .B(n6352), .Z(n6347) );
  XNOR U6765 ( .A(n6353), .B(n6354), .Z(n6352) );
  ANDN U6766 ( .B(n6346), .A(n6350), .Z(n6353) );
  ANDN U6767 ( .B(n6346), .A(n6343), .Z(n6344) );
  XNOR U6768 ( .A(n6349), .B(n6355), .Z(n6343) );
  XOR U6769 ( .A(n6356), .B(n6354), .Z(n6355) );
  NAND U6770 ( .A(n6357), .B(n6358), .Z(n6354) );
  XNOR U6771 ( .A(n6351), .B(n6334), .Z(n6358) );
  IV U6772 ( .A(n6346), .Z(n6351) );
  XNOR U6773 ( .A(n6337), .B(n6350), .Z(n6357) );
  IV U6774 ( .A(n6342), .Z(n6350) );
  XOR U6775 ( .A(n6359), .B(n6360), .Z(n6342) );
  XNOR U6776 ( .A(n6361), .B(n6362), .Z(n6360) );
  XNOR U6777 ( .A(n6363), .B(n6364), .Z(n6359) );
  NOR U6778 ( .A(n5956), .B(n5869), .Z(n6363) );
  AND U6779 ( .A(n6334), .B(n6337), .Z(n6356) );
  XNOR U6780 ( .A(n6334), .B(n6337), .Z(n6349) );
  XNOR U6781 ( .A(n6365), .B(n6366), .Z(n6337) );
  XNOR U6782 ( .A(n6367), .B(n6362), .Z(n6366) );
  XOR U6783 ( .A(n6368), .B(n6369), .Z(n6365) );
  XNOR U6784 ( .A(n6370), .B(n6364), .Z(n6369) );
  OR U6785 ( .A(n5955), .B(n6327), .Z(n6364) );
  XNOR U6786 ( .A(n5869), .B(n6326), .Z(n6327) );
  XNOR U6787 ( .A(n5956), .B(n5824), .Z(n5955) );
  ANDN U6788 ( .B(n6371), .A(n6326), .Z(n6370) );
  XNOR U6789 ( .A(n6372), .B(n6373), .Z(n6334) );
  XNOR U6790 ( .A(n6362), .B(n6374), .Z(n6373) );
  XOR U6791 ( .A(n5951), .B(n6368), .Z(n6374) );
  XNOR U6792 ( .A(n5869), .B(n6375), .Z(n6362) );
  XOR U6793 ( .A(n5829), .B(n6376), .Z(n6372) );
  XNOR U6794 ( .A(n6377), .B(n6378), .Z(n6376) );
  ANDN U6795 ( .B(n6379), .A(n6323), .Z(n6377) );
  XNOR U6796 ( .A(n6380), .B(n6381), .Z(n6346) );
  XNOR U6797 ( .A(n6367), .B(n6382), .Z(n6381) );
  XNOR U6798 ( .A(n5963), .B(n6361), .Z(n6382) );
  XOR U6799 ( .A(n6368), .B(n6383), .Z(n6361) );
  XNOR U6800 ( .A(n6384), .B(n6385), .Z(n6383) );
  NAND U6801 ( .A(n5876), .B(n5960), .Z(n6385) );
  XNOR U6802 ( .A(n6386), .B(n6384), .Z(n6368) );
  NANDN U6803 ( .A(n6329), .B(n5969), .Z(n6384) );
  XOR U6804 ( .A(n5970), .B(n5960), .Z(n5969) );
  XNOR U6805 ( .A(n6379), .B(n5824), .Z(n5960) );
  XOR U6806 ( .A(n6338), .B(n5876), .Z(n6329) );
  XNOR U6807 ( .A(n6323), .B(n6387), .Z(n5876) );
  ANDN U6808 ( .B(n5970), .A(n6338), .Z(n6386) );
  XNOR U6809 ( .A(n5829), .B(n5869), .Z(n6338) );
  XOR U6810 ( .A(n6388), .B(n6389), .Z(n5869) );
  XNOR U6811 ( .A(n6390), .B(n6391), .Z(n6389) );
  XOR U6812 ( .A(n6387), .B(n6371), .Z(n6367) );
  IV U6813 ( .A(n5824), .Z(n6371) );
  XOR U6814 ( .A(n6392), .B(n6393), .Z(n5824) );
  XOR U6815 ( .A(n6394), .B(n6391), .Z(n6393) );
  IV U6816 ( .A(n6326), .Z(n6387) );
  XOR U6817 ( .A(n6391), .B(n6395), .Z(n6326) );
  XNOR U6818 ( .A(n6396), .B(n6397), .Z(n6380) );
  XNOR U6819 ( .A(n6398), .B(n6378), .Z(n6397) );
  OR U6820 ( .A(n5966), .B(n6322), .Z(n6378) );
  XNOR U6821 ( .A(n5829), .B(n6323), .Z(n6322) );
  IV U6822 ( .A(n6396), .Z(n6323) );
  XOR U6823 ( .A(n5951), .B(n6379), .Z(n5966) );
  IV U6824 ( .A(n5963), .Z(n6379) );
  XOR U6825 ( .A(n6375), .B(n6399), .Z(n5963) );
  XOR U6826 ( .A(n6400), .B(n6401), .Z(n6388) );
  XNOR U6827 ( .A(n6402), .B(n6403), .Z(n6401) );
  XOR U6828 ( .A(n6404), .B(n6405), .Z(n6400) );
  XOR U6829 ( .A(key[922]), .B(n6406), .Z(n6405) );
  IV U6830 ( .A(n5956), .Z(n6375) );
  XOR U6831 ( .A(n6392), .B(n6407), .Z(n5956) );
  XOR U6832 ( .A(n6391), .B(n6408), .Z(n6407) );
  NOR U6833 ( .A(n5951), .B(n5829), .Z(n6398) );
  XOR U6834 ( .A(n6392), .B(n6409), .Z(n5951) );
  XOR U6835 ( .A(n6391), .B(n6410), .Z(n6409) );
  XOR U6836 ( .A(n6411), .B(n6412), .Z(n6391) );
  XOR U6837 ( .A(n5829), .B(n6413), .Z(n6412) );
  XNOR U6838 ( .A(n6414), .B(n6415), .Z(n6411) );
  XOR U6839 ( .A(key[926]), .B(n6416), .Z(n6415) );
  IV U6840 ( .A(n6395), .Z(n6392) );
  XOR U6841 ( .A(n6417), .B(n6418), .Z(n6395) );
  XNOR U6842 ( .A(n6419), .B(n6420), .Z(n6418) );
  XNOR U6843 ( .A(n6421), .B(n6422), .Z(n6417) );
  XOR U6844 ( .A(key[925]), .B(n6423), .Z(n6422) );
  XOR U6845 ( .A(n6424), .B(n6425), .Z(n6396) );
  XNOR U6846 ( .A(n6410), .B(n6408), .Z(n6425) );
  XNOR U6847 ( .A(n6426), .B(n6427), .Z(n6408) );
  XOR U6848 ( .A(n6428), .B(n6429), .Z(n6427) );
  XOR U6849 ( .A(key[927]), .B(n6430), .Z(n6426) );
  XNOR U6850 ( .A(n6431), .B(n6432), .Z(n6410) );
  XNOR U6851 ( .A(n6433), .B(n6434), .Z(n6432) );
  XNOR U6852 ( .A(n6435), .B(n6436), .Z(n6431) );
  XOR U6853 ( .A(key[924]), .B(n6437), .Z(n6436) );
  XNOR U6854 ( .A(n5829), .B(n6390), .Z(n6424) );
  XOR U6855 ( .A(n6438), .B(n6439), .Z(n6390) );
  XNOR U6856 ( .A(n6440), .B(n6441), .Z(n6439) );
  XOR U6857 ( .A(n6442), .B(n6394), .Z(n6441) );
  XNOR U6858 ( .A(n6443), .B(n6444), .Z(n6394) );
  XOR U6859 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U6860 ( .A(n6447), .B(n6448), .Z(n6443) );
  XNOR U6861 ( .A(key[921]), .B(n6449), .Z(n6448) );
  XNOR U6862 ( .A(n6450), .B(n6451), .Z(n6438) );
  XNOR U6863 ( .A(key[923]), .B(n6452), .Z(n6451) );
  XNOR U6864 ( .A(n6453), .B(n6454), .Z(n5829) );
  XNOR U6865 ( .A(n6455), .B(n6456), .Z(n6454) );
  XOR U6866 ( .A(n6457), .B(n6458), .Z(n6453) );
  XNOR U6867 ( .A(key[920]), .B(n6459), .Z(n6458) );
  XOR U6868 ( .A(n5853), .B(n5938), .Z(n3940) );
  XNOR U6869 ( .A(n5859), .B(n6460), .Z(n5938) );
  XNOR U6870 ( .A(n5856), .B(n6461), .Z(n6460) );
  NANDN U6871 ( .A(n6462), .B(n5843), .Z(n6461) );
  NANDN U6872 ( .A(n6463), .B(n5980), .Z(n5856) );
  XOR U6873 ( .A(n5857), .B(n5843), .Z(n5980) );
  XNOR U6874 ( .A(n5859), .B(n6464), .Z(n5853) );
  XOR U6875 ( .A(n6465), .B(n5835), .Z(n6464) );
  OR U6876 ( .A(n5991), .B(n6466), .Z(n5835) );
  XNOR U6877 ( .A(n5838), .B(n5990), .Z(n5991) );
  ANDN U6878 ( .B(n5990), .A(n6467), .Z(n6465) );
  XOR U6879 ( .A(n6468), .B(n5861), .Z(n5859) );
  OR U6880 ( .A(n5994), .B(n6469), .Z(n5861) );
  XOR U6881 ( .A(n6470), .B(n5863), .Z(n5994) );
  XNOR U6882 ( .A(n5990), .B(n5843), .Z(n5863) );
  XOR U6883 ( .A(n6471), .B(n6472), .Z(n5843) );
  NANDN U6884 ( .A(n6473), .B(n6474), .Z(n6472) );
  XOR U6885 ( .A(n6475), .B(n6476), .Z(n5990) );
  NANDN U6886 ( .A(n6473), .B(n6477), .Z(n6476) );
  ANDN U6887 ( .B(n6470), .A(n6478), .Z(n6468) );
  IV U6888 ( .A(n5997), .Z(n6470) );
  XNOR U6889 ( .A(n5857), .B(n5838), .Z(n5997) );
  XNOR U6890 ( .A(n6479), .B(n6475), .Z(n5838) );
  NANDN U6891 ( .A(n6480), .B(n6481), .Z(n6475) );
  XOR U6892 ( .A(n6477), .B(n6482), .Z(n6481) );
  ANDN U6893 ( .B(n6482), .A(n6483), .Z(n6479) );
  XNOR U6894 ( .A(n6484), .B(n6471), .Z(n5857) );
  NANDN U6895 ( .A(n6480), .B(n6485), .Z(n6471) );
  XOR U6896 ( .A(n6486), .B(n6474), .Z(n6485) );
  XNOR U6897 ( .A(n6487), .B(n6488), .Z(n6473) );
  XOR U6898 ( .A(n6489), .B(n6490), .Z(n6488) );
  XNOR U6899 ( .A(n6491), .B(n6492), .Z(n6487) );
  XNOR U6900 ( .A(n6493), .B(n6494), .Z(n6492) );
  ANDN U6901 ( .B(n6486), .A(n6490), .Z(n6493) );
  ANDN U6902 ( .B(n6486), .A(n6483), .Z(n6484) );
  XNOR U6903 ( .A(n6489), .B(n6495), .Z(n6483) );
  XOR U6904 ( .A(n6496), .B(n6494), .Z(n6495) );
  NAND U6905 ( .A(n6497), .B(n6498), .Z(n6494) );
  XNOR U6906 ( .A(n6491), .B(n6474), .Z(n6498) );
  IV U6907 ( .A(n6486), .Z(n6491) );
  XNOR U6908 ( .A(n6477), .B(n6490), .Z(n6497) );
  IV U6909 ( .A(n6482), .Z(n6490) );
  XOR U6910 ( .A(n6499), .B(n6500), .Z(n6482) );
  XNOR U6911 ( .A(n6501), .B(n6502), .Z(n6500) );
  XNOR U6912 ( .A(n6503), .B(n6504), .Z(n6499) );
  NOR U6913 ( .A(n5982), .B(n5858), .Z(n6503) );
  AND U6914 ( .A(n6474), .B(n6477), .Z(n6496) );
  XNOR U6915 ( .A(n6474), .B(n6477), .Z(n6489) );
  XNOR U6916 ( .A(n6505), .B(n6506), .Z(n6477) );
  XNOR U6917 ( .A(n6507), .B(n6502), .Z(n6506) );
  XOR U6918 ( .A(n6508), .B(n6509), .Z(n6505) );
  XNOR U6919 ( .A(n6510), .B(n6504), .Z(n6509) );
  OR U6920 ( .A(n5981), .B(n6463), .Z(n6504) );
  XNOR U6921 ( .A(n5858), .B(n6462), .Z(n6463) );
  XNOR U6922 ( .A(n5982), .B(n5844), .Z(n5981) );
  ANDN U6923 ( .B(n6511), .A(n6462), .Z(n6510) );
  XNOR U6924 ( .A(n6512), .B(n6513), .Z(n6474) );
  XNOR U6925 ( .A(n6502), .B(n6514), .Z(n6513) );
  XOR U6926 ( .A(n5977), .B(n6508), .Z(n6514) );
  XNOR U6927 ( .A(n5858), .B(n6515), .Z(n6502) );
  XOR U6928 ( .A(n5837), .B(n6516), .Z(n6512) );
  XNOR U6929 ( .A(n6517), .B(n6518), .Z(n6516) );
  ANDN U6930 ( .B(n6519), .A(n6467), .Z(n6517) );
  XNOR U6931 ( .A(n6520), .B(n6521), .Z(n6486) );
  XNOR U6932 ( .A(n6507), .B(n6522), .Z(n6521) );
  XNOR U6933 ( .A(n5989), .B(n6501), .Z(n6522) );
  XOR U6934 ( .A(n6508), .B(n6523), .Z(n6501) );
  XNOR U6935 ( .A(n6524), .B(n6525), .Z(n6523) );
  NAND U6936 ( .A(n5864), .B(n5986), .Z(n6525) );
  XNOR U6937 ( .A(n6526), .B(n6524), .Z(n6508) );
  NANDN U6938 ( .A(n6469), .B(n5995), .Z(n6524) );
  XOR U6939 ( .A(n5996), .B(n5986), .Z(n5995) );
  XNOR U6940 ( .A(n6519), .B(n5844), .Z(n5986) );
  XOR U6941 ( .A(n6478), .B(n5864), .Z(n6469) );
  XNOR U6942 ( .A(n6467), .B(n6527), .Z(n5864) );
  ANDN U6943 ( .B(n5996), .A(n6478), .Z(n6526) );
  XNOR U6944 ( .A(n5837), .B(n5858), .Z(n6478) );
  XOR U6945 ( .A(n6528), .B(n6529), .Z(n5858) );
  XNOR U6946 ( .A(n6530), .B(n6531), .Z(n6529) );
  XOR U6947 ( .A(n6527), .B(n6511), .Z(n6507) );
  IV U6948 ( .A(n5844), .Z(n6511) );
  XOR U6949 ( .A(n6532), .B(n6533), .Z(n5844) );
  XOR U6950 ( .A(n6534), .B(n6531), .Z(n6533) );
  IV U6951 ( .A(n6462), .Z(n6527) );
  XOR U6952 ( .A(n6531), .B(n6535), .Z(n6462) );
  XNOR U6953 ( .A(n6536), .B(n6537), .Z(n6520) );
  XNOR U6954 ( .A(n6538), .B(n6518), .Z(n6537) );
  OR U6955 ( .A(n5992), .B(n6466), .Z(n6518) );
  XNOR U6956 ( .A(n5837), .B(n6467), .Z(n6466) );
  IV U6957 ( .A(n6536), .Z(n6467) );
  XOR U6958 ( .A(n5977), .B(n6519), .Z(n5992) );
  IV U6959 ( .A(n5989), .Z(n6519) );
  XOR U6960 ( .A(n6515), .B(n6539), .Z(n5989) );
  XNOR U6961 ( .A(n6540), .B(n6528), .Z(n6539) );
  XOR U6962 ( .A(n6541), .B(n6542), .Z(n6528) );
  XNOR U6963 ( .A(n6543), .B(n6544), .Z(n6542) );
  XOR U6964 ( .A(key[930]), .B(n6545), .Z(n6541) );
  IV U6965 ( .A(n5982), .Z(n6515) );
  XOR U6966 ( .A(n6532), .B(n6546), .Z(n5982) );
  XOR U6967 ( .A(n6531), .B(n6547), .Z(n6546) );
  NOR U6968 ( .A(n5977), .B(n5837), .Z(n6538) );
  XOR U6969 ( .A(n6532), .B(n6548), .Z(n5977) );
  XOR U6970 ( .A(n6531), .B(n6549), .Z(n6548) );
  XOR U6971 ( .A(n6550), .B(n6551), .Z(n6531) );
  XNOR U6972 ( .A(n5837), .B(n6552), .Z(n6551) );
  XNOR U6973 ( .A(n6553), .B(n6554), .Z(n6550) );
  XNOR U6974 ( .A(key[934]), .B(n6555), .Z(n6554) );
  IV U6975 ( .A(n6535), .Z(n6532) );
  XOR U6976 ( .A(n6556), .B(n6557), .Z(n6535) );
  XNOR U6977 ( .A(n6558), .B(n6559), .Z(n6557) );
  XNOR U6978 ( .A(key[933]), .B(n6560), .Z(n6556) );
  XOR U6979 ( .A(n6561), .B(n6562), .Z(n6536) );
  XNOR U6980 ( .A(n6549), .B(n6547), .Z(n6562) );
  XNOR U6981 ( .A(n6563), .B(n6564), .Z(n6547) );
  XNOR U6982 ( .A(n6565), .B(n6566), .Z(n6564) );
  XNOR U6983 ( .A(key[935]), .B(n6567), .Z(n6563) );
  XNOR U6984 ( .A(n6568), .B(n6569), .Z(n6549) );
  XNOR U6985 ( .A(n6570), .B(n6571), .Z(n6568) );
  XNOR U6986 ( .A(key[932]), .B(n6572), .Z(n6571) );
  XNOR U6987 ( .A(n5837), .B(n6530), .Z(n6561) );
  XOR U6988 ( .A(n6573), .B(n6574), .Z(n6530) );
  XNOR U6989 ( .A(n6575), .B(n6576), .Z(n6574) );
  XNOR U6990 ( .A(n6577), .B(n6540), .Z(n6576) );
  IV U6991 ( .A(n6534), .Z(n6540) );
  XNOR U6992 ( .A(n6578), .B(n6579), .Z(n6534) );
  XOR U6993 ( .A(n6580), .B(n6581), .Z(n6579) );
  XOR U6994 ( .A(key[929]), .B(n6582), .Z(n6578) );
  XOR U6995 ( .A(n6583), .B(n6584), .Z(n6573) );
  XOR U6996 ( .A(key[931]), .B(n6585), .Z(n6584) );
  XNOR U6997 ( .A(n6586), .B(n6587), .Z(n5837) );
  XOR U6998 ( .A(n6588), .B(n6589), .Z(n6587) );
  XNOR U6999 ( .A(key[928]), .B(n6590), .Z(n6586) );
  IV U7000 ( .A(n5533), .Z(n438) );
  XOR U7001 ( .A(n5555), .B(n5604), .Z(n5533) );
  XNOR U7002 ( .A(n5549), .B(n6591), .Z(n5555) );
  XNOR U7003 ( .A(n6592), .B(n6593), .Z(n6591) );
  ANDN U7004 ( .B(n6594), .A(n5615), .Z(n6592) );
  IV U7005 ( .A(n6595), .Z(n5615) );
  XNOR U7006 ( .A(n6596), .B(n6597), .Z(n5549) );
  XNOR U7007 ( .A(n6598), .B(n6599), .Z(n6597) );
  NANDN U7008 ( .A(n6600), .B(n6601), .Z(n6599) );
  XNOR U7009 ( .A(n1080), .B(n1073), .Z(n428) );
  XNOR U7010 ( .A(n5475), .B(n5458), .Z(n1073) );
  XNOR U7011 ( .A(n5477), .B(n5478), .Z(n5458) );
  XOR U7012 ( .A(n5505), .B(n6602), .Z(n5478) );
  XNOR U7013 ( .A(n6603), .B(n6604), .Z(n6602) );
  NANDN U7014 ( .A(n6605), .B(n5570), .Z(n6604) );
  XNOR U7015 ( .A(n5564), .B(n6606), .Z(n5505) );
  XNOR U7016 ( .A(n6607), .B(n6608), .Z(n6606) );
  NANDN U7017 ( .A(n5591), .B(n6609), .Z(n6608) );
  XOR U7018 ( .A(n5587), .B(n6610), .Z(n5477) );
  XOR U7019 ( .A(n5584), .B(n6611), .Z(n6610) );
  NANDN U7020 ( .A(n6612), .B(n5574), .Z(n6611) );
  XOR U7021 ( .A(n5586), .B(n5574), .Z(n5576) );
  IV U7022 ( .A(n5504), .Z(n5475) );
  XOR U7023 ( .A(n5581), .B(n5459), .Z(n5504) );
  XOR U7024 ( .A(n5564), .B(n6614), .Z(n5459) );
  XNOR U7025 ( .A(n6603), .B(n6615), .Z(n6614) );
  NANDN U7026 ( .A(n6616), .B(n6617), .Z(n6615) );
  OR U7027 ( .A(n6618), .B(n6619), .Z(n6603) );
  XOR U7028 ( .A(n6620), .B(n6607), .Z(n5564) );
  NANDN U7029 ( .A(n6621), .B(n6622), .Z(n6607) );
  ANDN U7030 ( .B(n6623), .A(n6624), .Z(n6620) );
  XNOR U7031 ( .A(n5587), .B(n6625), .Z(n5581) );
  XOR U7032 ( .A(n6626), .B(n5567), .Z(n6625) );
  OR U7033 ( .A(n6627), .B(n6618), .Z(n5567) );
  XNOR U7034 ( .A(n5570), .B(n6617), .Z(n6618) );
  ANDN U7035 ( .B(n6628), .A(n6629), .Z(n6626) );
  XOR U7036 ( .A(n6630), .B(n5589), .Z(n5587) );
  OR U7037 ( .A(n6621), .B(n6631), .Z(n5589) );
  XNOR U7038 ( .A(n6624), .B(n5591), .Z(n6621) );
  XNOR U7039 ( .A(n6617), .B(n5574), .Z(n5591) );
  XOR U7040 ( .A(n6632), .B(n6633), .Z(n5574) );
  NANDN U7041 ( .A(n6634), .B(n6635), .Z(n6633) );
  IV U7042 ( .A(n6629), .Z(n6617) );
  XNOR U7043 ( .A(n6636), .B(n6637), .Z(n6629) );
  NANDN U7044 ( .A(n6634), .B(n6638), .Z(n6637) );
  NOR U7045 ( .A(n6624), .B(n6639), .Z(n6630) );
  XNOR U7046 ( .A(n5586), .B(n5570), .Z(n6624) );
  XNOR U7047 ( .A(n6640), .B(n6636), .Z(n5570) );
  NANDN U7048 ( .A(n6641), .B(n6642), .Z(n6636) );
  XOR U7049 ( .A(n6638), .B(n6643), .Z(n6642) );
  ANDN U7050 ( .B(n6643), .A(n6644), .Z(n6640) );
  XNOR U7051 ( .A(n6645), .B(n6632), .Z(n5586) );
  NANDN U7052 ( .A(n6641), .B(n6646), .Z(n6632) );
  XOR U7053 ( .A(n6647), .B(n6635), .Z(n6646) );
  XNOR U7054 ( .A(n6648), .B(n6649), .Z(n6634) );
  XOR U7055 ( .A(n6650), .B(n6651), .Z(n6649) );
  XNOR U7056 ( .A(n6652), .B(n6653), .Z(n6648) );
  XNOR U7057 ( .A(n6654), .B(n6655), .Z(n6653) );
  ANDN U7058 ( .B(n6647), .A(n6651), .Z(n6654) );
  ANDN U7059 ( .B(n6647), .A(n6644), .Z(n6645) );
  XNOR U7060 ( .A(n6650), .B(n6656), .Z(n6644) );
  XOR U7061 ( .A(n6657), .B(n6655), .Z(n6656) );
  NAND U7062 ( .A(n6658), .B(n6659), .Z(n6655) );
  XNOR U7063 ( .A(n6652), .B(n6635), .Z(n6659) );
  IV U7064 ( .A(n6647), .Z(n6652) );
  XNOR U7065 ( .A(n6638), .B(n6651), .Z(n6658) );
  IV U7066 ( .A(n6643), .Z(n6651) );
  XOR U7067 ( .A(n6660), .B(n6661), .Z(n6643) );
  XNOR U7068 ( .A(n6662), .B(n6663), .Z(n6661) );
  XNOR U7069 ( .A(n6664), .B(n6665), .Z(n6660) );
  ANDN U7070 ( .B(n5585), .A(n6666), .Z(n6664) );
  AND U7071 ( .A(n6635), .B(n6638), .Z(n6657) );
  XNOR U7072 ( .A(n6635), .B(n6638), .Z(n6650) );
  XNOR U7073 ( .A(n6667), .B(n6668), .Z(n6638) );
  XNOR U7074 ( .A(n6669), .B(n6663), .Z(n6668) );
  XOR U7075 ( .A(n6670), .B(n6671), .Z(n6667) );
  XNOR U7076 ( .A(n6672), .B(n6665), .Z(n6671) );
  OR U7077 ( .A(n5577), .B(n6613), .Z(n6665) );
  XNOR U7078 ( .A(n5585), .B(n6673), .Z(n6613) );
  XNOR U7079 ( .A(n6666), .B(n5575), .Z(n5577) );
  ANDN U7080 ( .B(n6674), .A(n6612), .Z(n6672) );
  XNOR U7081 ( .A(n6675), .B(n6676), .Z(n6635) );
  XNOR U7082 ( .A(n6663), .B(n6677), .Z(n6676) );
  XOR U7083 ( .A(n6605), .B(n6670), .Z(n6677) );
  XNOR U7084 ( .A(n5585), .B(n6666), .Z(n6663) );
  XNOR U7085 ( .A(n6678), .B(n6679), .Z(n6675) );
  XNOR U7086 ( .A(n6680), .B(n6681), .Z(n6679) );
  ANDN U7087 ( .B(n6628), .A(n6616), .Z(n6680) );
  XNOR U7088 ( .A(n6682), .B(n6683), .Z(n6647) );
  XNOR U7089 ( .A(n6669), .B(n6684), .Z(n6683) );
  XNOR U7090 ( .A(n6616), .B(n6662), .Z(n6684) );
  XOR U7091 ( .A(n6670), .B(n6685), .Z(n6662) );
  XNOR U7092 ( .A(n6686), .B(n6687), .Z(n6685) );
  NAND U7093 ( .A(n5592), .B(n6609), .Z(n6687) );
  XNOR U7094 ( .A(n6688), .B(n6686), .Z(n6670) );
  NANDN U7095 ( .A(n6631), .B(n6622), .Z(n6686) );
  XOR U7096 ( .A(n6623), .B(n6609), .Z(n6622) );
  XNOR U7097 ( .A(n6689), .B(n5575), .Z(n6609) );
  XOR U7098 ( .A(n6639), .B(n5592), .Z(n6631) );
  XOR U7099 ( .A(n6628), .B(n6673), .Z(n5592) );
  ANDN U7100 ( .B(n6623), .A(n6639), .Z(n6688) );
  XNOR U7101 ( .A(n6678), .B(n5585), .Z(n6639) );
  XNOR U7102 ( .A(n6690), .B(n6691), .Z(n5585) );
  XNOR U7103 ( .A(n6692), .B(n6693), .Z(n6691) );
  XOR U7104 ( .A(n6694), .B(n5509), .Z(n6623) );
  XOR U7105 ( .A(n6673), .B(n6674), .Z(n6669) );
  IV U7106 ( .A(n5575), .Z(n6674) );
  XOR U7107 ( .A(n6695), .B(n6696), .Z(n5575) );
  XNOR U7108 ( .A(n6697), .B(n6693), .Z(n6696) );
  IV U7109 ( .A(n6612), .Z(n6673) );
  XOR U7110 ( .A(n6693), .B(n6698), .Z(n6612) );
  XNOR U7111 ( .A(n6628), .B(n6699), .Z(n6682) );
  XNOR U7112 ( .A(n6700), .B(n6681), .Z(n6699) );
  OR U7113 ( .A(n6619), .B(n6627), .Z(n6681) );
  XNOR U7114 ( .A(n6678), .B(n6628), .Z(n6627) );
  XOR U7115 ( .A(n6605), .B(n6689), .Z(n6619) );
  IV U7116 ( .A(n6616), .Z(n6689) );
  XOR U7117 ( .A(n5509), .B(n6701), .Z(n6616) );
  XNOR U7118 ( .A(n6697), .B(n6690), .Z(n6701) );
  XOR U7119 ( .A(n6702), .B(n6703), .Z(n6690) );
  XNOR U7120 ( .A(n4067), .B(n3147), .Z(n6703) );
  XOR U7121 ( .A(n4104), .B(n4066), .Z(n3147) );
  XOR U7122 ( .A(n6704), .B(n6705), .Z(n4104) );
  XNOR U7123 ( .A(n6706), .B(n6707), .Z(n6705) );
  XNOR U7124 ( .A(n6708), .B(n6709), .Z(n6704) );
  IV U7125 ( .A(n3150), .Z(n4067) );
  XOR U7126 ( .A(n4111), .B(n3113), .Z(n3150) );
  XOR U7127 ( .A(key[1090]), .B(n4112), .Z(n6702) );
  IV U7128 ( .A(n6666), .Z(n5509) );
  XOR U7129 ( .A(n6695), .B(n6710), .Z(n6666) );
  XOR U7130 ( .A(n6693), .B(n6711), .Z(n6710) );
  ANDN U7131 ( .B(n6694), .A(n5569), .Z(n6700) );
  IV U7132 ( .A(n6605), .Z(n6694) );
  XOR U7133 ( .A(n6695), .B(n6712), .Z(n6605) );
  XOR U7134 ( .A(n6693), .B(n6713), .Z(n6712) );
  XOR U7135 ( .A(n6714), .B(n6715), .Z(n6693) );
  XOR U7136 ( .A(n5350), .B(n5569), .Z(n6715) );
  IV U7137 ( .A(n6678), .Z(n5569) );
  XOR U7138 ( .A(n5358), .B(n4093), .Z(n5350) );
  XNOR U7139 ( .A(n6716), .B(n6717), .Z(n4093) );
  XNOR U7140 ( .A(n6706), .B(n6718), .Z(n6717) );
  XNOR U7141 ( .A(n6719), .B(n6709), .Z(n6716) );
  XNOR U7142 ( .A(n4084), .B(n6720), .Z(n6714) );
  XNOR U7143 ( .A(key[1094]), .B(n4076), .Z(n6720) );
  XNOR U7144 ( .A(n3130), .B(n6721), .Z(n4076) );
  XOR U7145 ( .A(n4087), .B(n3123), .Z(n3130) );
  XNOR U7146 ( .A(n6722), .B(n6723), .Z(n3123) );
  XOR U7147 ( .A(n6724), .B(n6725), .Z(n6723) );
  XOR U7148 ( .A(n6726), .B(n6727), .Z(n4087) );
  IV U7149 ( .A(n6698), .Z(n6695) );
  XOR U7150 ( .A(n6728), .B(n6729), .Z(n6698) );
  XNOR U7151 ( .A(n4085), .B(n5351), .Z(n6729) );
  XNOR U7152 ( .A(n4079), .B(n4084), .Z(n5351) );
  XNOR U7153 ( .A(n6707), .B(n6732), .Z(n4079) );
  XOR U7154 ( .A(n6733), .B(n6708), .Z(n6732) );
  XNOR U7155 ( .A(n6734), .B(n6735), .Z(n6707) );
  XNOR U7156 ( .A(n6736), .B(n6737), .Z(n6735) );
  NANDN U7157 ( .A(n6738), .B(n6739), .Z(n6737) );
  XOR U7158 ( .A(n4101), .B(n3128), .Z(n4085) );
  XNOR U7159 ( .A(n6740), .B(n6741), .Z(n3128) );
  XNOR U7160 ( .A(n6742), .B(n6743), .Z(n6741) );
  XNOR U7161 ( .A(n6744), .B(n6745), .Z(n6740) );
  XOR U7162 ( .A(n6746), .B(n6747), .Z(n6745) );
  ANDN U7163 ( .B(n6748), .A(n6749), .Z(n6747) );
  XOR U7164 ( .A(n6750), .B(n6751), .Z(n4101) );
  XNOR U7165 ( .A(n6752), .B(n6753), .Z(n6751) );
  XNOR U7166 ( .A(n6754), .B(n6755), .Z(n6750) );
  XOR U7167 ( .A(n6756), .B(n6757), .Z(n6755) );
  ANDN U7168 ( .B(n6758), .A(n6759), .Z(n6757) );
  XNOR U7169 ( .A(key[1093]), .B(n5345), .Z(n6728) );
  XOR U7170 ( .A(n6760), .B(n6761), .Z(n6628) );
  XNOR U7171 ( .A(n6713), .B(n6711), .Z(n6761) );
  XNOR U7172 ( .A(n6762), .B(n6763), .Z(n6711) );
  XNOR U7173 ( .A(n6721), .B(n4094), .Z(n6763) );
  XNOR U7174 ( .A(n4078), .B(n5352), .Z(n4094) );
  XNOR U7175 ( .A(n6764), .B(n6765), .Z(n5352) );
  XOR U7176 ( .A(n6766), .B(n6743), .Z(n6765) );
  XNOR U7177 ( .A(n6767), .B(n6768), .Z(n6743) );
  XNOR U7178 ( .A(n6769), .B(n6770), .Z(n6768) );
  OR U7179 ( .A(n6771), .B(n6772), .Z(n6770) );
  XNOR U7180 ( .A(n6773), .B(n6774), .Z(n6764) );
  XNOR U7181 ( .A(n6775), .B(n6776), .Z(n4078) );
  XNOR U7182 ( .A(n6726), .B(n6753), .Z(n6776) );
  XNOR U7183 ( .A(n6777), .B(n6778), .Z(n6753) );
  XNOR U7184 ( .A(n6779), .B(n6780), .Z(n6778) );
  NANDN U7185 ( .A(n6781), .B(n6782), .Z(n6780) );
  XOR U7186 ( .A(n6783), .B(n6784), .Z(n6775) );
  XOR U7187 ( .A(n6785), .B(n5341), .Z(n6721) );
  XOR U7188 ( .A(n6786), .B(n6787), .Z(n5341) );
  XOR U7189 ( .A(n6731), .B(n6788), .Z(n6787) );
  XOR U7190 ( .A(n6789), .B(n6790), .Z(n6786) );
  XOR U7191 ( .A(key[1095]), .B(n5342), .Z(n6762) );
  IV U7192 ( .A(n5358), .Z(n5342) );
  XNOR U7193 ( .A(n6791), .B(n6792), .Z(n6713) );
  XOR U7194 ( .A(n4098), .B(n5331), .Z(n6792) );
  XOR U7195 ( .A(n5358), .B(n4083), .Z(n5331) );
  XNOR U7196 ( .A(n6793), .B(n6794), .Z(n4083) );
  XNOR U7197 ( .A(n6795), .B(n6718), .Z(n6794) );
  XNOR U7198 ( .A(n6796), .B(n6797), .Z(n6718) );
  XNOR U7199 ( .A(n6798), .B(n6799), .Z(n6797) );
  OR U7200 ( .A(n6800), .B(n6801), .Z(n6799) );
  XNOR U7201 ( .A(n6802), .B(n6803), .Z(n6793) );
  XNOR U7202 ( .A(n6804), .B(n6736), .Z(n6803) );
  NANDN U7203 ( .A(n6805), .B(n6806), .Z(n6736) );
  ANDN U7204 ( .B(n6807), .A(n6808), .Z(n6804) );
  XNOR U7205 ( .A(n4115), .B(n3140), .Z(n4098) );
  XNOR U7206 ( .A(n6744), .B(n3113), .Z(n3140) );
  XOR U7207 ( .A(n6724), .B(n6774), .Z(n3113) );
  XOR U7208 ( .A(n6754), .B(n4111), .Z(n4115) );
  XNOR U7209 ( .A(n6809), .B(n6783), .Z(n4111) );
  XNOR U7210 ( .A(n4099), .B(n6810), .Z(n6791) );
  XNOR U7211 ( .A(key[1092]), .B(n5329), .Z(n6810) );
  XOR U7212 ( .A(n6785), .B(n5345), .Z(n4099) );
  XOR U7213 ( .A(n6811), .B(n6812), .Z(n5345) );
  XNOR U7214 ( .A(n6813), .B(n6788), .Z(n6812) );
  XNOR U7215 ( .A(n6814), .B(n6815), .Z(n6788) );
  XNOR U7216 ( .A(n6816), .B(n6817), .Z(n6815) );
  OR U7217 ( .A(n6818), .B(n6819), .Z(n6817) );
  XNOR U7218 ( .A(n6820), .B(n6821), .Z(n6811) );
  XNOR U7219 ( .A(n6822), .B(n6823), .Z(n6821) );
  ANDN U7220 ( .B(n6824), .A(n6825), .Z(n6823) );
  XOR U7221 ( .A(n6678), .B(n6692), .Z(n6760) );
  XOR U7222 ( .A(n6826), .B(n6827), .Z(n6692) );
  XNOR U7223 ( .A(n6697), .B(n6828), .Z(n6827) );
  XOR U7224 ( .A(n4066), .B(n5365), .Z(n6828) );
  XNOR U7225 ( .A(n5358), .B(n4097), .Z(n5365) );
  XOR U7226 ( .A(n6802), .B(n4065), .Z(n4097) );
  XOR U7227 ( .A(n6733), .B(n6802), .Z(n5358) );
  XNOR U7228 ( .A(n6796), .B(n6829), .Z(n6802) );
  XNOR U7229 ( .A(n6830), .B(n6831), .Z(n6829) );
  ANDN U7230 ( .B(n6739), .A(n6832), .Z(n6830) );
  XNOR U7231 ( .A(n6833), .B(n6834), .Z(n6796) );
  XNOR U7232 ( .A(n6835), .B(n6836), .Z(n6834) );
  NANDN U7233 ( .A(n6837), .B(n6838), .Z(n6836) );
  XNOR U7234 ( .A(n6839), .B(n6840), .Z(n4066) );
  XOR U7235 ( .A(n6841), .B(n6730), .Z(n6840) );
  XOR U7236 ( .A(n6842), .B(n6843), .Z(n6730) );
  XOR U7237 ( .A(n6844), .B(n6822), .Z(n6843) );
  NANDN U7238 ( .A(n6845), .B(n6846), .Z(n6822) );
  ANDN U7239 ( .B(n6847), .A(n6848), .Z(n6844) );
  XNOR U7240 ( .A(n6849), .B(n6790), .Z(n6839) );
  XOR U7241 ( .A(n6850), .B(n6851), .Z(n6697) );
  XOR U7242 ( .A(n3159), .B(n3114), .Z(n6851) );
  XOR U7243 ( .A(n4112), .B(n4065), .Z(n3114) );
  XOR U7244 ( .A(n6733), .B(n6709), .Z(n4065) );
  IV U7245 ( .A(n6852), .Z(n6733) );
  XOR U7246 ( .A(n4118), .B(n3152), .Z(n3159) );
  IV U7247 ( .A(n5356), .Z(n3152) );
  XOR U7248 ( .A(n6766), .B(n6853), .Z(n5356) );
  XOR U7249 ( .A(n6773), .B(n6774), .Z(n6853) );
  XNOR U7250 ( .A(n6854), .B(n6725), .Z(n6773) );
  IV U7251 ( .A(n6855), .Z(n6766) );
  XNOR U7252 ( .A(n6726), .B(n6856), .Z(n4118) );
  XOR U7253 ( .A(n6783), .B(n6857), .Z(n6856) );
  XNOR U7254 ( .A(n6809), .B(n6858), .Z(n6726) );
  XNOR U7255 ( .A(key[1089]), .B(n4119), .Z(n6850) );
  XNOR U7256 ( .A(n4106), .B(n6859), .Z(n6826) );
  XNOR U7257 ( .A(key[1091]), .B(n4113), .Z(n6859) );
  XOR U7258 ( .A(n6785), .B(n5329), .Z(n4113) );
  XOR U7259 ( .A(n6813), .B(n4112), .Z(n5329) );
  XNOR U7260 ( .A(n6789), .B(n6860), .Z(n4112) );
  IV U7261 ( .A(n3115), .Z(n4106) );
  XOR U7262 ( .A(n4069), .B(n3153), .Z(n3115) );
  XOR U7263 ( .A(n6861), .B(n6862), .Z(n3153) );
  XNOR U7264 ( .A(n6855), .B(n6722), .Z(n6862) );
  XNOR U7265 ( .A(n6863), .B(n6864), .Z(n6722) );
  XNOR U7266 ( .A(n6865), .B(n6746), .Z(n6864) );
  NOR U7267 ( .A(n6866), .B(n6867), .Z(n6746) );
  NOR U7268 ( .A(n6868), .B(n6869), .Z(n6865) );
  XOR U7269 ( .A(n6871), .B(n6872), .Z(n6870) );
  NOR U7270 ( .A(n6873), .B(n6771), .Z(n6871) );
  XNOR U7271 ( .A(n6742), .B(n6874), .Z(n6863) );
  XNOR U7272 ( .A(n6875), .B(n6876), .Z(n6874) );
  NAND U7273 ( .A(n6877), .B(n6878), .Z(n6876) );
  XNOR U7274 ( .A(n6725), .B(n6774), .Z(n6861) );
  XOR U7275 ( .A(n6879), .B(n6880), .Z(n6774) );
  XNOR U7276 ( .A(n6881), .B(n6882), .Z(n6880) );
  NANDN U7277 ( .A(n6749), .B(n6883), .Z(n6882) );
  XNOR U7278 ( .A(n6742), .B(n6884), .Z(n6725) );
  XNOR U7279 ( .A(n6872), .B(n6885), .Z(n6884) );
  NANDN U7280 ( .A(n6886), .B(n6887), .Z(n6885) );
  OR U7281 ( .A(n6888), .B(n6889), .Z(n6872) );
  XOR U7282 ( .A(n6890), .B(n6875), .Z(n6742) );
  NANDN U7283 ( .A(n6891), .B(n6892), .Z(n6875) );
  AND U7284 ( .A(n6893), .B(n6894), .Z(n6890) );
  XOR U7285 ( .A(n6895), .B(n6896), .Z(n4069) );
  XNOR U7286 ( .A(n6858), .B(n6727), .Z(n6896) );
  XNOR U7287 ( .A(n6897), .B(n6898), .Z(n6727) );
  XNOR U7288 ( .A(n6899), .B(n6756), .Z(n6898) );
  ANDN U7289 ( .B(n6900), .A(n6901), .Z(n6756) );
  ANDN U7290 ( .B(n6902), .A(n6903), .Z(n6899) );
  XNOR U7291 ( .A(n6752), .B(n6904), .Z(n6858) );
  XNOR U7292 ( .A(n6905), .B(n6906), .Z(n6904) );
  NANDN U7293 ( .A(n6907), .B(n6908), .Z(n6906) );
  XNOR U7294 ( .A(n6783), .B(n6857), .Z(n6895) );
  IV U7295 ( .A(n6784), .Z(n6857) );
  XOR U7296 ( .A(n6897), .B(n6909), .Z(n6784) );
  XNOR U7297 ( .A(n6905), .B(n6910), .Z(n6909) );
  NANDN U7298 ( .A(n6911), .B(n6782), .Z(n6910) );
  OR U7299 ( .A(n6912), .B(n6913), .Z(n6905) );
  XNOR U7300 ( .A(n6752), .B(n6914), .Z(n6897) );
  XNOR U7301 ( .A(n6915), .B(n6916), .Z(n6914) );
  NANDN U7302 ( .A(n6917), .B(n6918), .Z(n6916) );
  XOR U7303 ( .A(n6919), .B(n6915), .Z(n6752) );
  NANDN U7304 ( .A(n6920), .B(n6921), .Z(n6915) );
  ANDN U7305 ( .B(n6922), .A(n6923), .Z(n6919) );
  XOR U7306 ( .A(n6924), .B(n6925), .Z(n6783) );
  XOR U7307 ( .A(n6926), .B(n6927), .Z(n6925) );
  NANDN U7308 ( .A(n6928), .B(n6758), .Z(n6927) );
  XOR U7309 ( .A(n6929), .B(n6930), .Z(n6678) );
  XNOR U7310 ( .A(n4092), .B(n3151), .Z(n6930) );
  XNOR U7311 ( .A(n4119), .B(n4109), .Z(n3151) );
  XOR U7312 ( .A(n6706), .B(n6931), .Z(n4109) );
  XOR U7313 ( .A(n6719), .B(n6709), .Z(n6931) );
  XOR U7314 ( .A(n6833), .B(n6932), .Z(n6709) );
  XOR U7315 ( .A(n6831), .B(n6933), .Z(n6932) );
  NAND U7316 ( .A(n6934), .B(n6807), .Z(n6933) );
  ANDN U7317 ( .B(n6806), .A(n6935), .Z(n6831) );
  XOR U7318 ( .A(n6739), .B(n6807), .Z(n6806) );
  XNOR U7319 ( .A(n6852), .B(n6708), .Z(n6719) );
  XNOR U7320 ( .A(n6795), .B(n6936), .Z(n6708) );
  XOR U7321 ( .A(n6937), .B(n6938), .Z(n6936) );
  AND U7322 ( .A(n6939), .B(n6940), .Z(n6937) );
  XNOR U7323 ( .A(n6833), .B(n6941), .Z(n6852) );
  XOR U7324 ( .A(n6942), .B(n6798), .Z(n6941) );
  OR U7325 ( .A(n6943), .B(n6944), .Z(n6798) );
  ANDN U7326 ( .B(n6940), .A(n6945), .Z(n6942) );
  XOR U7327 ( .A(n6946), .B(n6835), .Z(n6833) );
  OR U7328 ( .A(n6947), .B(n6948), .Z(n6835) );
  ANDN U7329 ( .B(n6949), .A(n6950), .Z(n6946) );
  XNOR U7330 ( .A(n6734), .B(n6951), .Z(n6706) );
  XNOR U7331 ( .A(n6938), .B(n6952), .Z(n6951) );
  OR U7332 ( .A(n6800), .B(n6953), .Z(n6952) );
  OR U7333 ( .A(n6944), .B(n6954), .Z(n6938) );
  XOR U7334 ( .A(n6800), .B(n6940), .Z(n6944) );
  XNOR U7335 ( .A(n6795), .B(n6955), .Z(n6734) );
  XNOR U7336 ( .A(n6956), .B(n6957), .Z(n6955) );
  NANDN U7337 ( .A(n6837), .B(n6958), .Z(n6957) );
  XOR U7338 ( .A(n6959), .B(n6956), .Z(n6795) );
  NANDN U7339 ( .A(n6947), .B(n6960), .Z(n6956) );
  XOR U7340 ( .A(n6949), .B(n6837), .Z(n6947) );
  XNOR U7341 ( .A(n6940), .B(n6807), .Z(n6837) );
  XOR U7342 ( .A(n6961), .B(n6962), .Z(n6807) );
  NANDN U7343 ( .A(n6963), .B(n6964), .Z(n6962) );
  XOR U7344 ( .A(n6965), .B(n6966), .Z(n6940) );
  OR U7345 ( .A(n6963), .B(n6967), .Z(n6966) );
  IV U7346 ( .A(n6968), .Z(n6949) );
  ANDN U7347 ( .B(n6969), .A(n6968), .Z(n6959) );
  XOR U7348 ( .A(n6800), .B(n6739), .Z(n6968) );
  XNOR U7349 ( .A(n6970), .B(n6961), .Z(n6739) );
  NANDN U7350 ( .A(n6971), .B(n6972), .Z(n6961) );
  ANDN U7351 ( .B(n6973), .A(n6974), .Z(n6970) );
  NANDN U7352 ( .A(n6971), .B(n6976), .Z(n6965) );
  XOR U7353 ( .A(n6977), .B(n6963), .Z(n6971) );
  XNOR U7354 ( .A(n6978), .B(n6979), .Z(n6963) );
  XOR U7355 ( .A(n6980), .B(n6973), .Z(n6979) );
  XNOR U7356 ( .A(n6981), .B(n6982), .Z(n6978) );
  XNOR U7357 ( .A(n6983), .B(n6984), .Z(n6982) );
  ANDN U7358 ( .B(n6973), .A(n6985), .Z(n6983) );
  IV U7359 ( .A(n6986), .Z(n6973) );
  ANDN U7360 ( .B(n6977), .A(n6985), .Z(n6975) );
  IV U7361 ( .A(n6981), .Z(n6985) );
  IV U7362 ( .A(n6974), .Z(n6977) );
  XNOR U7363 ( .A(n6980), .B(n6987), .Z(n6974) );
  XOR U7364 ( .A(n6988), .B(n6984), .Z(n6987) );
  NAND U7365 ( .A(n6976), .B(n6972), .Z(n6984) );
  XNOR U7366 ( .A(n6964), .B(n6986), .Z(n6972) );
  XOR U7367 ( .A(n6989), .B(n6990), .Z(n6986) );
  XOR U7368 ( .A(n6991), .B(n6992), .Z(n6990) );
  XNOR U7369 ( .A(n6939), .B(n6993), .Z(n6992) );
  XNOR U7370 ( .A(n6994), .B(n6995), .Z(n6989) );
  XNOR U7371 ( .A(n6996), .B(n6997), .Z(n6995) );
  ANDN U7372 ( .B(n6998), .A(n6801), .Z(n6996) );
  XNOR U7373 ( .A(n6981), .B(n6967), .Z(n6976) );
  XOR U7374 ( .A(n6999), .B(n7000), .Z(n6981) );
  XNOR U7375 ( .A(n7001), .B(n6993), .Z(n7000) );
  XOR U7376 ( .A(n7002), .B(n7003), .Z(n6993) );
  XNOR U7377 ( .A(n7004), .B(n7005), .Z(n7003) );
  NAND U7378 ( .A(n6838), .B(n6958), .Z(n7005) );
  XNOR U7379 ( .A(n7006), .B(n7007), .Z(n6999) );
  ANDN U7380 ( .B(n7008), .A(n6832), .Z(n7006) );
  ANDN U7381 ( .B(n6964), .A(n6967), .Z(n6988) );
  XOR U7382 ( .A(n6967), .B(n6964), .Z(n6980) );
  XNOR U7383 ( .A(n7009), .B(n7010), .Z(n6964) );
  XNOR U7384 ( .A(n7002), .B(n7011), .Z(n7010) );
  XOR U7385 ( .A(n7001), .B(n6953), .Z(n7011) );
  XOR U7386 ( .A(n6801), .B(n7012), .Z(n7009) );
  XNOR U7387 ( .A(n7013), .B(n6997), .Z(n7012) );
  OR U7388 ( .A(n6954), .B(n6943), .Z(n6997) );
  XNOR U7389 ( .A(n6801), .B(n6945), .Z(n6943) );
  XOR U7390 ( .A(n6953), .B(n6939), .Z(n6954) );
  ANDN U7391 ( .B(n6939), .A(n6945), .Z(n7013) );
  XOR U7392 ( .A(n7014), .B(n7015), .Z(n6967) );
  XOR U7393 ( .A(n7002), .B(n6991), .Z(n7015) );
  XOR U7394 ( .A(n6934), .B(n6808), .Z(n6991) );
  XOR U7395 ( .A(n7016), .B(n7004), .Z(n7002) );
  NANDN U7396 ( .A(n6948), .B(n6960), .Z(n7004) );
  XOR U7397 ( .A(n6969), .B(n6958), .Z(n6960) );
  XNOR U7398 ( .A(n7008), .B(n7017), .Z(n6939) );
  XOR U7399 ( .A(n7018), .B(n7019), .Z(n7017) );
  XOR U7400 ( .A(n6950), .B(n6838), .Z(n6948) );
  XNOR U7401 ( .A(n6945), .B(n6934), .Z(n6838) );
  IV U7402 ( .A(n6994), .Z(n6945) );
  XOR U7403 ( .A(n7020), .B(n7021), .Z(n6994) );
  XOR U7404 ( .A(n7022), .B(n7023), .Z(n7021) );
  XNOR U7405 ( .A(n6801), .B(n7024), .Z(n7020) );
  ANDN U7406 ( .B(n6969), .A(n6950), .Z(n7016) );
  XNOR U7407 ( .A(n6801), .B(n6832), .Z(n6950) );
  XOR U7408 ( .A(n7001), .B(n7025), .Z(n7014) );
  XNOR U7409 ( .A(n7026), .B(n7007), .Z(n7025) );
  OR U7410 ( .A(n6805), .B(n6935), .Z(n7007) );
  XNOR U7411 ( .A(n7027), .B(n6934), .Z(n6935) );
  XNOR U7412 ( .A(n6738), .B(n6808), .Z(n6805) );
  ANDN U7413 ( .B(n6934), .A(n6808), .Z(n7026) );
  XOR U7414 ( .A(n7028), .B(n7029), .Z(n6808) );
  XNOR U7415 ( .A(n7019), .B(n7030), .Z(n7029) );
  XOR U7416 ( .A(n7031), .B(n7028), .Z(n6934) );
  XNOR U7417 ( .A(n6832), .B(n6738), .Z(n7001) );
  IV U7418 ( .A(n7027), .Z(n6832) );
  XOR U7419 ( .A(n7030), .B(n7032), .Z(n7027) );
  XNOR U7420 ( .A(n7018), .B(n7024), .Z(n7032) );
  XOR U7421 ( .A(n7033), .B(n7034), .Z(n7024) );
  XNOR U7422 ( .A(n7035), .B(n7036), .Z(n7034) );
  XNOR U7423 ( .A(n7019), .B(n6106), .Z(n7036) );
  XNOR U7424 ( .A(n7037), .B(n7038), .Z(n7019) );
  XNOR U7425 ( .A(n6150), .B(n6105), .Z(n7038) );
  XNOR U7426 ( .A(key[993]), .B(n7039), .Z(n7037) );
  XNOR U7427 ( .A(n7040), .B(n7041), .Z(n7033) );
  XNOR U7428 ( .A(key[995]), .B(n7042), .Z(n7041) );
  XOR U7429 ( .A(n7043), .B(n7044), .Z(n7018) );
  XOR U7430 ( .A(n7045), .B(n6147), .Z(n7044) );
  XOR U7431 ( .A(key[994]), .B(n7046), .Z(n7043) );
  IV U7432 ( .A(n7031), .Z(n7030) );
  XOR U7433 ( .A(n7008), .B(n6998), .Z(n6969) );
  IV U7434 ( .A(n6953), .Z(n6998) );
  XOR U7435 ( .A(n7028), .B(n7047), .Z(n6953) );
  XOR U7436 ( .A(n7031), .B(n7023), .Z(n7047) );
  XNOR U7437 ( .A(n7048), .B(n7049), .Z(n7023) );
  XOR U7438 ( .A(n7050), .B(n7051), .Z(n7049) );
  XNOR U7439 ( .A(n7052), .B(n7053), .Z(n7048) );
  XNOR U7440 ( .A(key[996]), .B(n7054), .Z(n7053) );
  IV U7441 ( .A(n6738), .Z(n7008) );
  XOR U7442 ( .A(n7028), .B(n7055), .Z(n6738) );
  XNOR U7443 ( .A(n7031), .B(n7022), .Z(n7055) );
  XOR U7444 ( .A(n7056), .B(n7057), .Z(n7022) );
  XNOR U7445 ( .A(n7058), .B(n7059), .Z(n7057) );
  XNOR U7446 ( .A(key[999]), .B(n7060), .Z(n7056) );
  XOR U7447 ( .A(n7061), .B(n7062), .Z(n7031) );
  XOR U7448 ( .A(n7063), .B(n7064), .Z(n7062) );
  XNOR U7449 ( .A(n7065), .B(n7066), .Z(n7061) );
  XOR U7450 ( .A(key[998]), .B(n6801), .Z(n7066) );
  XNOR U7451 ( .A(n7067), .B(n7068), .Z(n6801) );
  XOR U7452 ( .A(n7069), .B(n6144), .Z(n7068) );
  XOR U7453 ( .A(key[992]), .B(n7070), .Z(n7067) );
  XNOR U7454 ( .A(n7071), .B(n7072), .Z(n7028) );
  XOR U7455 ( .A(n7073), .B(n7074), .Z(n7072) );
  XOR U7456 ( .A(key[997]), .B(n7075), .Z(n7071) );
  XOR U7457 ( .A(n6731), .B(n7076), .Z(n4119) );
  XOR U7458 ( .A(n6849), .B(n6790), .Z(n7076) );
  XOR U7459 ( .A(n6842), .B(n7077), .Z(n6790) );
  XNOR U7460 ( .A(n7078), .B(n7079), .Z(n7077) );
  NANDN U7461 ( .A(n6818), .B(n7080), .Z(n7079) );
  XNOR U7462 ( .A(n6820), .B(n7081), .Z(n6842) );
  XNOR U7463 ( .A(n7082), .B(n7083), .Z(n7081) );
  NAND U7464 ( .A(n7084), .B(n7085), .Z(n7083) );
  IV U7465 ( .A(n6789), .Z(n6849) );
  XOR U7466 ( .A(n7086), .B(n7087), .Z(n6789) );
  XNOR U7467 ( .A(n7088), .B(n7089), .Z(n7087) );
  NAND U7468 ( .A(n7090), .B(n6824), .Z(n7089) );
  XOR U7469 ( .A(n6841), .B(n6860), .Z(n6731) );
  XNOR U7470 ( .A(n6820), .B(n7091), .Z(n6841) );
  XNOR U7471 ( .A(n7078), .B(n7092), .Z(n7091) );
  NANDN U7472 ( .A(n7093), .B(n7094), .Z(n7092) );
  OR U7473 ( .A(n7095), .B(n7096), .Z(n7078) );
  XOR U7474 ( .A(n7097), .B(n7082), .Z(n6820) );
  NANDN U7475 ( .A(n7098), .B(n7099), .Z(n7082) );
  ANDN U7476 ( .B(n7100), .A(n7101), .Z(n7097) );
  XOR U7477 ( .A(n3137), .B(n6785), .Z(n4092) );
  IV U7478 ( .A(n3158), .Z(n6785) );
  XNOR U7479 ( .A(n6814), .B(n7102), .Z(n6813) );
  XOR U7480 ( .A(n7103), .B(n7088), .Z(n7102) );
  NANDN U7481 ( .A(n7104), .B(n6846), .Z(n7088) );
  XOR U7482 ( .A(n6847), .B(n6824), .Z(n6846) );
  ANDN U7483 ( .B(n6847), .A(n7105), .Z(n7103) );
  XNOR U7484 ( .A(n7086), .B(n7106), .Z(n6814) );
  XNOR U7485 ( .A(n7107), .B(n7108), .Z(n7106) );
  NAND U7486 ( .A(n7085), .B(n7109), .Z(n7108) );
  XNOR U7487 ( .A(n7086), .B(n7110), .Z(n6860) );
  XOR U7488 ( .A(n7111), .B(n6816), .Z(n7110) );
  OR U7489 ( .A(n7095), .B(n7112), .Z(n6816) );
  XNOR U7490 ( .A(n6818), .B(n7093), .Z(n7095) );
  NOR U7491 ( .A(n7113), .B(n7093), .Z(n7111) );
  XOR U7492 ( .A(n7114), .B(n7107), .Z(n7086) );
  OR U7493 ( .A(n7098), .B(n7115), .Z(n7107) );
  XOR U7494 ( .A(n7101), .B(n7085), .Z(n7098) );
  XNOR U7495 ( .A(n7093), .B(n6824), .Z(n7085) );
  XOR U7496 ( .A(n7116), .B(n7117), .Z(n6824) );
  NANDN U7497 ( .A(n7118), .B(n7119), .Z(n7117) );
  XNOR U7498 ( .A(n7120), .B(n7121), .Z(n7093) );
  OR U7499 ( .A(n7118), .B(n7122), .Z(n7121) );
  ANDN U7500 ( .B(n7123), .A(n7101), .Z(n7114) );
  XOR U7501 ( .A(n6818), .B(n6847), .Z(n7101) );
  XNOR U7502 ( .A(n7124), .B(n7116), .Z(n6847) );
  NANDN U7503 ( .A(n7125), .B(n7126), .Z(n7116) );
  ANDN U7504 ( .B(n7127), .A(n7128), .Z(n7124) );
  NANDN U7505 ( .A(n7125), .B(n7130), .Z(n7120) );
  XOR U7506 ( .A(n7131), .B(n7118), .Z(n7125) );
  XNOR U7507 ( .A(n7132), .B(n7133), .Z(n7118) );
  XOR U7508 ( .A(n7134), .B(n7127), .Z(n7133) );
  XNOR U7509 ( .A(n7135), .B(n7136), .Z(n7132) );
  XNOR U7510 ( .A(n7137), .B(n7138), .Z(n7136) );
  ANDN U7511 ( .B(n7127), .A(n7139), .Z(n7137) );
  IV U7512 ( .A(n7140), .Z(n7127) );
  ANDN U7513 ( .B(n7131), .A(n7139), .Z(n7129) );
  IV U7514 ( .A(n7135), .Z(n7139) );
  IV U7515 ( .A(n7128), .Z(n7131) );
  XNOR U7516 ( .A(n7134), .B(n7141), .Z(n7128) );
  XOR U7517 ( .A(n7142), .B(n7138), .Z(n7141) );
  NAND U7518 ( .A(n7130), .B(n7126), .Z(n7138) );
  XNOR U7519 ( .A(n7119), .B(n7140), .Z(n7126) );
  XOR U7520 ( .A(n7143), .B(n7144), .Z(n7140) );
  XOR U7521 ( .A(n7145), .B(n7146), .Z(n7144) );
  XNOR U7522 ( .A(n7094), .B(n7147), .Z(n7146) );
  XNOR U7523 ( .A(n7148), .B(n7149), .Z(n7143) );
  XNOR U7524 ( .A(n7150), .B(n7151), .Z(n7149) );
  ANDN U7525 ( .B(n7080), .A(n6819), .Z(n7150) );
  XNOR U7526 ( .A(n7135), .B(n7122), .Z(n7130) );
  XOR U7527 ( .A(n7152), .B(n7153), .Z(n7135) );
  XNOR U7528 ( .A(n7154), .B(n7147), .Z(n7153) );
  XOR U7529 ( .A(n7155), .B(n7156), .Z(n7147) );
  XNOR U7530 ( .A(n7157), .B(n7158), .Z(n7156) );
  NAND U7531 ( .A(n7109), .B(n7084), .Z(n7158) );
  XNOR U7532 ( .A(n7159), .B(n7160), .Z(n7152) );
  ANDN U7533 ( .B(n7161), .A(n7105), .Z(n7159) );
  ANDN U7534 ( .B(n7119), .A(n7122), .Z(n7142) );
  XOR U7535 ( .A(n7122), .B(n7119), .Z(n7134) );
  XNOR U7536 ( .A(n7162), .B(n7163), .Z(n7119) );
  XNOR U7537 ( .A(n7155), .B(n7164), .Z(n7163) );
  XNOR U7538 ( .A(n7154), .B(n7080), .Z(n7164) );
  XNOR U7539 ( .A(n7165), .B(n7166), .Z(n7162) );
  XNOR U7540 ( .A(n7167), .B(n7151), .Z(n7166) );
  OR U7541 ( .A(n7096), .B(n7112), .Z(n7151) );
  XNOR U7542 ( .A(n7165), .B(n7148), .Z(n7112) );
  XNOR U7543 ( .A(n7080), .B(n7094), .Z(n7096) );
  ANDN U7544 ( .B(n7094), .A(n7113), .Z(n7167) );
  XOR U7545 ( .A(n7168), .B(n7169), .Z(n7122) );
  XOR U7546 ( .A(n7155), .B(n7145), .Z(n7169) );
  XOR U7547 ( .A(n7090), .B(n6825), .Z(n7145) );
  XOR U7548 ( .A(n7170), .B(n7157), .Z(n7155) );
  NANDN U7549 ( .A(n7115), .B(n7099), .Z(n7157) );
  XOR U7550 ( .A(n7100), .B(n7084), .Z(n7099) );
  XNOR U7551 ( .A(n7161), .B(n7171), .Z(n7094) );
  XNOR U7552 ( .A(n7172), .B(n7173), .Z(n7171) );
  XNOR U7553 ( .A(n7123), .B(n7109), .Z(n7115) );
  XNOR U7554 ( .A(n7113), .B(n7090), .Z(n7109) );
  IV U7555 ( .A(n7148), .Z(n7113) );
  XOR U7556 ( .A(n7174), .B(n7175), .Z(n7148) );
  XOR U7557 ( .A(n7176), .B(n7177), .Z(n7175) );
  XOR U7558 ( .A(n7165), .B(n7178), .Z(n7174) );
  AND U7559 ( .A(n7100), .B(n7123), .Z(n7170) );
  XOR U7560 ( .A(n7161), .B(n7080), .Z(n7100) );
  XNOR U7561 ( .A(n7179), .B(n7180), .Z(n7080) );
  XOR U7562 ( .A(n7181), .B(n7177), .Z(n7180) );
  XNOR U7563 ( .A(n7182), .B(n7183), .Z(n7177) );
  XOR U7564 ( .A(n7184), .B(n7185), .Z(n7183) );
  XNOR U7565 ( .A(n7186), .B(n7187), .Z(n7182) );
  XNOR U7566 ( .A(key[988]), .B(n7188), .Z(n7187) );
  IV U7567 ( .A(n6848), .Z(n7161) );
  XOR U7568 ( .A(n7154), .B(n7189), .Z(n7168) );
  XNOR U7569 ( .A(n7190), .B(n7160), .Z(n7189) );
  OR U7570 ( .A(n6845), .B(n7104), .Z(n7160) );
  XNOR U7571 ( .A(n7191), .B(n7090), .Z(n7104) );
  XNOR U7572 ( .A(n6848), .B(n6825), .Z(n6845) );
  ANDN U7573 ( .B(n7090), .A(n6825), .Z(n7190) );
  XOR U7574 ( .A(n7179), .B(n7192), .Z(n6825) );
  XOR U7575 ( .A(n7172), .B(n7193), .Z(n7192) );
  XOR U7576 ( .A(n7181), .B(n7179), .Z(n7090) );
  XNOR U7577 ( .A(n7105), .B(n6848), .Z(n7154) );
  XOR U7578 ( .A(n7179), .B(n7194), .Z(n6848) );
  XNOR U7579 ( .A(n7181), .B(n7176), .Z(n7194) );
  XOR U7580 ( .A(n7195), .B(n7196), .Z(n7176) );
  XNOR U7581 ( .A(n7197), .B(n6316), .Z(n7196) );
  XOR U7582 ( .A(key[991]), .B(n7198), .Z(n7195) );
  XNOR U7583 ( .A(n7199), .B(n7200), .Z(n7179) );
  XOR U7584 ( .A(n7201), .B(n7202), .Z(n7200) );
  XOR U7585 ( .A(n7203), .B(n7204), .Z(n7199) );
  XOR U7586 ( .A(key[989]), .B(n6276), .Z(n7204) );
  XOR U7587 ( .A(n6819), .B(n7105), .Z(n7123) );
  IV U7588 ( .A(n7191), .Z(n7105) );
  XNOR U7589 ( .A(n7173), .B(n7205), .Z(n7191) );
  XOR U7590 ( .A(n7178), .B(n7193), .Z(n7205) );
  IV U7591 ( .A(n7181), .Z(n7193) );
  XOR U7592 ( .A(n7206), .B(n7207), .Z(n7181) );
  XNOR U7593 ( .A(n6283), .B(n7208), .Z(n7207) );
  XNOR U7594 ( .A(n7209), .B(n7210), .Z(n7206) );
  XNOR U7595 ( .A(key[990]), .B(n7165), .Z(n7210) );
  XOR U7596 ( .A(n7211), .B(n7212), .Z(n7178) );
  XNOR U7597 ( .A(n7213), .B(n7214), .Z(n7212) );
  XNOR U7598 ( .A(n7172), .B(n7215), .Z(n7214) );
  XOR U7599 ( .A(n7216), .B(n7217), .Z(n7172) );
  XOR U7600 ( .A(n6262), .B(n6315), .Z(n7217) );
  XNOR U7601 ( .A(n7218), .B(n7219), .Z(n7216) );
  XNOR U7602 ( .A(key[985]), .B(n7220), .Z(n7219) );
  XNOR U7603 ( .A(n7221), .B(n7222), .Z(n7211) );
  XNOR U7604 ( .A(key[987]), .B(n6266), .Z(n7222) );
  XOR U7605 ( .A(n7223), .B(n7224), .Z(n7173) );
  XOR U7606 ( .A(n7225), .B(n7226), .Z(n7224) );
  XOR U7607 ( .A(n6307), .B(n7227), .Z(n7223) );
  XOR U7608 ( .A(key[986]), .B(n7228), .Z(n7227) );
  IV U7609 ( .A(n7165), .Z(n6819) );
  XOR U7610 ( .A(n7229), .B(n7230), .Z(n7165) );
  XOR U7611 ( .A(n7231), .B(n7232), .Z(n7230) );
  XOR U7612 ( .A(n7233), .B(n7234), .Z(n7229) );
  XOR U7613 ( .A(key[984]), .B(n6290), .Z(n7234) );
  XOR U7614 ( .A(n6754), .B(n6809), .Z(n3137) );
  XNOR U7615 ( .A(n6924), .B(n7235), .Z(n6809) );
  XOR U7616 ( .A(n7236), .B(n6779), .Z(n7235) );
  OR U7617 ( .A(n7237), .B(n6912), .Z(n6779) );
  XNOR U7618 ( .A(n6782), .B(n6908), .Z(n6912) );
  ANDN U7619 ( .B(n6908), .A(n7238), .Z(n7236) );
  XNOR U7620 ( .A(n6777), .B(n7239), .Z(n6754) );
  XNOR U7621 ( .A(n7240), .B(n6926), .Z(n7239) );
  XOR U7622 ( .A(n7242), .B(n6758), .Z(n6900) );
  ANDN U7623 ( .B(n7243), .A(n6903), .Z(n7240) );
  IV U7624 ( .A(n7242), .Z(n6903) );
  XNOR U7625 ( .A(n6924), .B(n7244), .Z(n6777) );
  XNOR U7626 ( .A(n7245), .B(n7246), .Z(n7244) );
  NANDN U7627 ( .A(n6917), .B(n7247), .Z(n7246) );
  XOR U7628 ( .A(n7248), .B(n7245), .Z(n6924) );
  OR U7629 ( .A(n6920), .B(n7249), .Z(n7245) );
  XNOR U7630 ( .A(n6923), .B(n6917), .Z(n6920) );
  XNOR U7631 ( .A(n6908), .B(n6758), .Z(n6917) );
  XOR U7632 ( .A(n7250), .B(n7251), .Z(n6758) );
  NANDN U7633 ( .A(n7252), .B(n7253), .Z(n7251) );
  XOR U7634 ( .A(n7254), .B(n7255), .Z(n6908) );
  NANDN U7635 ( .A(n7252), .B(n7256), .Z(n7255) );
  NOR U7636 ( .A(n6923), .B(n7257), .Z(n7248) );
  XNOR U7637 ( .A(n7242), .B(n6782), .Z(n6923) );
  XNOR U7638 ( .A(n7258), .B(n7254), .Z(n6782) );
  NANDN U7639 ( .A(n7259), .B(n7260), .Z(n7254) );
  XOR U7640 ( .A(n7256), .B(n7261), .Z(n7260) );
  ANDN U7641 ( .B(n7261), .A(n7262), .Z(n7258) );
  XNOR U7642 ( .A(n7263), .B(n7250), .Z(n7242) );
  NANDN U7643 ( .A(n7259), .B(n7264), .Z(n7250) );
  XOR U7644 ( .A(n7265), .B(n7253), .Z(n7264) );
  XNOR U7645 ( .A(n7266), .B(n7267), .Z(n7252) );
  XOR U7646 ( .A(n7268), .B(n7269), .Z(n7267) );
  XNOR U7647 ( .A(n7270), .B(n7271), .Z(n7266) );
  XNOR U7648 ( .A(n7272), .B(n7273), .Z(n7271) );
  ANDN U7649 ( .B(n7265), .A(n7269), .Z(n7272) );
  ANDN U7650 ( .B(n7265), .A(n7262), .Z(n7263) );
  XNOR U7651 ( .A(n7268), .B(n7274), .Z(n7262) );
  XOR U7652 ( .A(n7275), .B(n7273), .Z(n7274) );
  NAND U7653 ( .A(n7276), .B(n7277), .Z(n7273) );
  XNOR U7654 ( .A(n7270), .B(n7253), .Z(n7277) );
  IV U7655 ( .A(n7265), .Z(n7270) );
  XNOR U7656 ( .A(n7256), .B(n7269), .Z(n7276) );
  IV U7657 ( .A(n7261), .Z(n7269) );
  XOR U7658 ( .A(n7278), .B(n7279), .Z(n7261) );
  XNOR U7659 ( .A(n7280), .B(n7281), .Z(n7279) );
  XNOR U7660 ( .A(n7282), .B(n7283), .Z(n7278) );
  ANDN U7661 ( .B(n7243), .A(n7284), .Z(n7282) );
  AND U7662 ( .A(n7253), .B(n7256), .Z(n7275) );
  XNOR U7663 ( .A(n7253), .B(n7256), .Z(n7268) );
  XNOR U7664 ( .A(n7285), .B(n7286), .Z(n7256) );
  XNOR U7665 ( .A(n7287), .B(n7281), .Z(n7286) );
  XOR U7666 ( .A(n7288), .B(n7289), .Z(n7285) );
  XNOR U7667 ( .A(n7290), .B(n7283), .Z(n7289) );
  OR U7668 ( .A(n6901), .B(n7241), .Z(n7283) );
  XNOR U7669 ( .A(n7243), .B(n7291), .Z(n7241) );
  XNOR U7670 ( .A(n7284), .B(n6759), .Z(n6901) );
  ANDN U7671 ( .B(n7292), .A(n6928), .Z(n7290) );
  XNOR U7672 ( .A(n7293), .B(n7294), .Z(n7253) );
  XNOR U7673 ( .A(n7281), .B(n7295), .Z(n7294) );
  XOR U7674 ( .A(n6911), .B(n7288), .Z(n7295) );
  XNOR U7675 ( .A(n7243), .B(n7284), .Z(n7281) );
  XOR U7676 ( .A(n6781), .B(n7296), .Z(n7293) );
  XNOR U7677 ( .A(n7297), .B(n7298), .Z(n7296) );
  ANDN U7678 ( .B(n7299), .A(n7238), .Z(n7297) );
  XNOR U7679 ( .A(n7300), .B(n7301), .Z(n7265) );
  XNOR U7680 ( .A(n7287), .B(n7302), .Z(n7301) );
  XNOR U7681 ( .A(n6907), .B(n7280), .Z(n7302) );
  XOR U7682 ( .A(n7288), .B(n7303), .Z(n7280) );
  XNOR U7683 ( .A(n7304), .B(n7305), .Z(n7303) );
  NAND U7684 ( .A(n7247), .B(n6918), .Z(n7305) );
  XNOR U7685 ( .A(n7306), .B(n7304), .Z(n7288) );
  NANDN U7686 ( .A(n7249), .B(n6921), .Z(n7304) );
  XOR U7687 ( .A(n6922), .B(n6918), .Z(n6921) );
  XNOR U7688 ( .A(n7299), .B(n6759), .Z(n6918) );
  XOR U7689 ( .A(n7257), .B(n7247), .Z(n7249) );
  XNOR U7690 ( .A(n7238), .B(n7291), .Z(n7247) );
  ANDN U7691 ( .B(n6922), .A(n7257), .Z(n7306) );
  XOR U7692 ( .A(n6781), .B(n7243), .Z(n7257) );
  XNOR U7693 ( .A(n7307), .B(n7308), .Z(n7243) );
  XNOR U7694 ( .A(n7309), .B(n7310), .Z(n7308) );
  XOR U7695 ( .A(n7291), .B(n7292), .Z(n7287) );
  IV U7696 ( .A(n6759), .Z(n7292) );
  XOR U7697 ( .A(n7311), .B(n7312), .Z(n6759) );
  XNOR U7698 ( .A(n7313), .B(n7310), .Z(n7312) );
  IV U7699 ( .A(n6928), .Z(n7291) );
  XOR U7700 ( .A(n7310), .B(n7314), .Z(n6928) );
  XNOR U7701 ( .A(n7315), .B(n7316), .Z(n7300) );
  XNOR U7702 ( .A(n7317), .B(n7298), .Z(n7316) );
  OR U7703 ( .A(n6913), .B(n7237), .Z(n7298) );
  XNOR U7704 ( .A(n6781), .B(n7238), .Z(n7237) );
  IV U7705 ( .A(n7315), .Z(n7238) );
  XOR U7706 ( .A(n6911), .B(n7299), .Z(n6913) );
  IV U7707 ( .A(n6907), .Z(n7299) );
  XOR U7708 ( .A(n6902), .B(n7318), .Z(n6907) );
  XNOR U7709 ( .A(n7313), .B(n7307), .Z(n7318) );
  XOR U7710 ( .A(n7319), .B(n7320), .Z(n7307) );
  XNOR U7711 ( .A(n6581), .B(n6583), .Z(n7320) );
  XOR U7712 ( .A(key[946]), .B(n7321), .Z(n7319) );
  IV U7713 ( .A(n7284), .Z(n6902) );
  XOR U7714 ( .A(n7311), .B(n7322), .Z(n7284) );
  XOR U7715 ( .A(n7310), .B(n7323), .Z(n7322) );
  NOR U7716 ( .A(n6911), .B(n6781), .Z(n7317) );
  XOR U7717 ( .A(n7311), .B(n7324), .Z(n6911) );
  XOR U7718 ( .A(n7310), .B(n7325), .Z(n7324) );
  XOR U7719 ( .A(n7326), .B(n7327), .Z(n7310) );
  XOR U7720 ( .A(n7328), .B(n7329), .Z(n7327) );
  XNOR U7721 ( .A(n7330), .B(n7331), .Z(n7326) );
  XOR U7722 ( .A(key[950]), .B(n6781), .Z(n7331) );
  IV U7723 ( .A(n7314), .Z(n7311) );
  XOR U7724 ( .A(n7332), .B(n7333), .Z(n7314) );
  XOR U7725 ( .A(n7334), .B(n7335), .Z(n7333) );
  XOR U7726 ( .A(key[949]), .B(n7336), .Z(n7332) );
  XOR U7727 ( .A(n7337), .B(n7338), .Z(n7315) );
  XNOR U7728 ( .A(n7325), .B(n7323), .Z(n7338) );
  XNOR U7729 ( .A(n7339), .B(n7340), .Z(n7323) );
  XNOR U7730 ( .A(n7341), .B(n7342), .Z(n7340) );
  XNOR U7731 ( .A(key[951]), .B(n7343), .Z(n7339) );
  XNOR U7732 ( .A(n7344), .B(n7345), .Z(n7325) );
  XOR U7733 ( .A(n7346), .B(n7347), .Z(n7345) );
  XNOR U7734 ( .A(n7348), .B(n7349), .Z(n7344) );
  XNOR U7735 ( .A(key[948]), .B(n7350), .Z(n7349) );
  XNOR U7736 ( .A(n6781), .B(n7309), .Z(n7337) );
  XOR U7737 ( .A(n7351), .B(n7352), .Z(n7309) );
  XNOR U7738 ( .A(n7353), .B(n7354), .Z(n7352) );
  XOR U7739 ( .A(n7313), .B(n7355), .Z(n7354) );
  XOR U7740 ( .A(n7356), .B(n7357), .Z(n7313) );
  XNOR U7741 ( .A(key[945]), .B(n7358), .Z(n7356) );
  XNOR U7742 ( .A(n7359), .B(n7360), .Z(n7351) );
  XNOR U7743 ( .A(key[947]), .B(n7361), .Z(n7360) );
  XNOR U7744 ( .A(n7362), .B(n7363), .Z(n6781) );
  XOR U7745 ( .A(n7364), .B(n6582), .Z(n7363) );
  XOR U7746 ( .A(key[944]), .B(n7365), .Z(n7362) );
  XNOR U7747 ( .A(key[1088]), .B(n5330), .Z(n6929) );
  XOR U7748 ( .A(n6724), .B(n6744), .Z(n5330) );
  XNOR U7749 ( .A(n6767), .B(n7366), .Z(n6744) );
  XNOR U7750 ( .A(n6881), .B(n7367), .Z(n7366) );
  OR U7751 ( .A(n6869), .B(n7368), .Z(n7367) );
  OR U7752 ( .A(n7369), .B(n6866), .Z(n6881) );
  XOR U7753 ( .A(n6869), .B(n7370), .Z(n6866) );
  XNOR U7754 ( .A(n6879), .B(n7371), .Z(n6767) );
  XNOR U7755 ( .A(n7372), .B(n7373), .Z(n7371) );
  NAND U7756 ( .A(n6878), .B(n7374), .Z(n7373) );
  IV U7757 ( .A(n6854), .Z(n6724) );
  XNOR U7758 ( .A(n6879), .B(n7375), .Z(n6854) );
  XOR U7759 ( .A(n7376), .B(n6769), .Z(n7375) );
  OR U7760 ( .A(n7377), .B(n6888), .Z(n6769) );
  XNOR U7761 ( .A(n6771), .B(n6886), .Z(n6888) );
  NOR U7762 ( .A(n7378), .B(n6886), .Z(n7376) );
  XOR U7763 ( .A(n7379), .B(n7372), .Z(n6879) );
  OR U7764 ( .A(n6891), .B(n7380), .Z(n7372) );
  XNOR U7765 ( .A(n6893), .B(n6878), .Z(n6891) );
  XOR U7766 ( .A(n6886), .B(n6749), .Z(n6878) );
  IV U7767 ( .A(n7370), .Z(n6749) );
  XOR U7768 ( .A(n7381), .B(n7382), .Z(n7370) );
  NANDN U7769 ( .A(n7383), .B(n7384), .Z(n7382) );
  XNOR U7770 ( .A(n7385), .B(n7386), .Z(n6886) );
  OR U7771 ( .A(n7383), .B(n7387), .Z(n7386) );
  ANDN U7772 ( .B(n6893), .A(n7388), .Z(n7379) );
  XOR U7773 ( .A(n6771), .B(n6869), .Z(n6893) );
  XNOR U7774 ( .A(n7381), .B(n7389), .Z(n6869) );
  NANDN U7775 ( .A(n7390), .B(n7391), .Z(n7389) );
  NANDN U7776 ( .A(n7392), .B(n7393), .Z(n7381) );
  OR U7777 ( .A(n7395), .B(n7392), .Z(n7385) );
  XOR U7778 ( .A(n7396), .B(n7383), .Z(n7392) );
  XNOR U7779 ( .A(n7397), .B(n7398), .Z(n7383) );
  XOR U7780 ( .A(n7399), .B(n7391), .Z(n7398) );
  XNOR U7781 ( .A(n7400), .B(n7401), .Z(n7397) );
  XNOR U7782 ( .A(n7402), .B(n7403), .Z(n7401) );
  ANDN U7783 ( .B(n7391), .A(n7404), .Z(n7402) );
  IV U7784 ( .A(n7405), .Z(n7391) );
  ANDN U7785 ( .B(n7396), .A(n7404), .Z(n7394) );
  IV U7786 ( .A(n7390), .Z(n7396) );
  XNOR U7787 ( .A(n7399), .B(n7406), .Z(n7390) );
  XNOR U7788 ( .A(n7403), .B(n7407), .Z(n7406) );
  NANDN U7789 ( .A(n7387), .B(n7384), .Z(n7407) );
  NANDN U7790 ( .A(n7395), .B(n7393), .Z(n7403) );
  XNOR U7791 ( .A(n7384), .B(n7405), .Z(n7393) );
  XOR U7792 ( .A(n7408), .B(n7409), .Z(n7405) );
  XOR U7793 ( .A(n7410), .B(n7411), .Z(n7409) );
  XNOR U7794 ( .A(n6887), .B(n7412), .Z(n7411) );
  XNOR U7795 ( .A(n7413), .B(n7414), .Z(n7408) );
  XNOR U7796 ( .A(n7415), .B(n7416), .Z(n7414) );
  ANDN U7797 ( .B(n7417), .A(n6772), .Z(n7415) );
  XNOR U7798 ( .A(n7404), .B(n7387), .Z(n7395) );
  IV U7799 ( .A(n7400), .Z(n7404) );
  XOR U7800 ( .A(n7418), .B(n7419), .Z(n7400) );
  XNOR U7801 ( .A(n7420), .B(n7412), .Z(n7419) );
  XOR U7802 ( .A(n7421), .B(n7422), .Z(n7412) );
  XNOR U7803 ( .A(n7423), .B(n7424), .Z(n7422) );
  NAND U7804 ( .A(n7374), .B(n6877), .Z(n7424) );
  XNOR U7805 ( .A(n7425), .B(n7426), .Z(n7418) );
  ANDN U7806 ( .B(n7427), .A(n7368), .Z(n7425) );
  XOR U7807 ( .A(n7387), .B(n7384), .Z(n7399) );
  XNOR U7808 ( .A(n7428), .B(n7429), .Z(n7384) );
  XNOR U7809 ( .A(n7421), .B(n7430), .Z(n7429) );
  XOR U7810 ( .A(n7420), .B(n6873), .Z(n7430) );
  XOR U7811 ( .A(n6772), .B(n7431), .Z(n7428) );
  XNOR U7812 ( .A(n7432), .B(n7416), .Z(n7431) );
  OR U7813 ( .A(n6889), .B(n7377), .Z(n7416) );
  XNOR U7814 ( .A(n6772), .B(n7378), .Z(n7377) );
  XOR U7815 ( .A(n6873), .B(n6887), .Z(n6889) );
  ANDN U7816 ( .B(n6887), .A(n7378), .Z(n7432) );
  XOR U7817 ( .A(n7433), .B(n7434), .Z(n7387) );
  XOR U7818 ( .A(n7421), .B(n7410), .Z(n7434) );
  XNOR U7819 ( .A(n6883), .B(n6748), .Z(n7410) );
  XOR U7820 ( .A(n7435), .B(n7423), .Z(n7421) );
  NANDN U7821 ( .A(n7380), .B(n6892), .Z(n7423) );
  XOR U7822 ( .A(n6894), .B(n6877), .Z(n6892) );
  XOR U7823 ( .A(n6748), .B(n6887), .Z(n6877) );
  XNOR U7824 ( .A(n7427), .B(n7436), .Z(n6887) );
  XOR U7825 ( .A(n7437), .B(n7438), .Z(n7436) );
  XOR U7826 ( .A(n7388), .B(n7374), .Z(n7380) );
  XNOR U7827 ( .A(n7378), .B(n6883), .Z(n7374) );
  IV U7828 ( .A(n7413), .Z(n7378) );
  XOR U7829 ( .A(n7439), .B(n7440), .Z(n7413) );
  XOR U7830 ( .A(n7441), .B(n7442), .Z(n7440) );
  XNOR U7831 ( .A(n6772), .B(n7443), .Z(n7439) );
  ANDN U7832 ( .B(n6894), .A(n7388), .Z(n7435) );
  XNOR U7833 ( .A(n6772), .B(n7368), .Z(n7388) );
  XOR U7834 ( .A(n7427), .B(n7417), .Z(n6894) );
  IV U7835 ( .A(n6873), .Z(n7417) );
  XOR U7836 ( .A(n7444), .B(n7445), .Z(n6873) );
  XOR U7837 ( .A(n7446), .B(n7442), .Z(n7445) );
  XNOR U7838 ( .A(n7447), .B(n7448), .Z(n7442) );
  XOR U7839 ( .A(n7449), .B(n7450), .Z(n7448) );
  XNOR U7840 ( .A(key[908]), .B(n7451), .Z(n7447) );
  XOR U7841 ( .A(n7420), .B(n7452), .Z(n7433) );
  XNOR U7842 ( .A(n7453), .B(n7426), .Z(n7452) );
  OR U7843 ( .A(n6867), .B(n7369), .Z(n7426) );
  XNOR U7844 ( .A(n7454), .B(n6883), .Z(n7369) );
  XNOR U7845 ( .A(n7427), .B(n6748), .Z(n6867) );
  IV U7846 ( .A(n6868), .Z(n7427) );
  AND U7847 ( .A(n6748), .B(n6883), .Z(n7453) );
  XOR U7848 ( .A(n7446), .B(n7444), .Z(n6883) );
  XNOR U7849 ( .A(n7444), .B(n7455), .Z(n6748) );
  XNOR U7850 ( .A(n7438), .B(n7456), .Z(n7455) );
  XNOR U7851 ( .A(n7368), .B(n6868), .Z(n7420) );
  XOR U7852 ( .A(n7444), .B(n7457), .Z(n6868) );
  XNOR U7853 ( .A(n7446), .B(n7441), .Z(n7457) );
  XOR U7854 ( .A(n7458), .B(n7459), .Z(n7441) );
  XNOR U7855 ( .A(n7460), .B(n6456), .Z(n7459) );
  XOR U7856 ( .A(key[911]), .B(n7461), .Z(n7458) );
  XNOR U7857 ( .A(n7462), .B(n7463), .Z(n7444) );
  XOR U7858 ( .A(n7464), .B(n7465), .Z(n7463) );
  XOR U7859 ( .A(n7466), .B(n7467), .Z(n7462) );
  XOR U7860 ( .A(key[909]), .B(n6416), .Z(n7467) );
  IV U7861 ( .A(n7454), .Z(n7368) );
  XOR U7862 ( .A(n7456), .B(n7468), .Z(n7454) );
  XNOR U7863 ( .A(n7437), .B(n7443), .Z(n7468) );
  XOR U7864 ( .A(n7469), .B(n7470), .Z(n7443) );
  XNOR U7865 ( .A(n7471), .B(n7472), .Z(n7470) );
  XNOR U7866 ( .A(n7438), .B(n6402), .Z(n7472) );
  XNOR U7867 ( .A(n7473), .B(n7474), .Z(n7438) );
  XNOR U7868 ( .A(n7475), .B(n6455), .Z(n7474) );
  XNOR U7869 ( .A(n7476), .B(n7477), .Z(n7473) );
  XOR U7870 ( .A(key[905]), .B(n6406), .Z(n7477) );
  XNOR U7871 ( .A(n7478), .B(n7479), .Z(n7469) );
  XNOR U7872 ( .A(key[907]), .B(n7480), .Z(n7479) );
  XOR U7873 ( .A(n7481), .B(n7482), .Z(n7437) );
  XOR U7874 ( .A(n7483), .B(n7484), .Z(n7482) );
  XOR U7875 ( .A(n7485), .B(n7486), .Z(n7481) );
  XOR U7876 ( .A(key[906]), .B(n6447), .Z(n7486) );
  IV U7877 ( .A(n7446), .Z(n7456) );
  XOR U7878 ( .A(n7487), .B(n7488), .Z(n7446) );
  XNOR U7879 ( .A(n6423), .B(n7489), .Z(n7488) );
  XNOR U7880 ( .A(n7490), .B(n7491), .Z(n7487) );
  XOR U7881 ( .A(key[910]), .B(n6772), .Z(n7491) );
  XNOR U7882 ( .A(n7492), .B(n7493), .Z(n6772) );
  XOR U7883 ( .A(n7494), .B(n7495), .Z(n7493) );
  XOR U7884 ( .A(n7496), .B(n7497), .Z(n7492) );
  XOR U7885 ( .A(key[904]), .B(n6430), .Z(n7497) );
  IV U7886 ( .A(n5595), .Z(n1080) );
  XOR U7887 ( .A(n5536), .B(n5607), .Z(n5595) );
  XNOR U7888 ( .A(n5538), .B(n5539), .Z(n5607) );
  XOR U7889 ( .A(n5609), .B(n7498), .Z(n5539) );
  XNOR U7890 ( .A(n7499), .B(n7500), .Z(n7498) );
  NANDN U7891 ( .A(n7501), .B(n5554), .Z(n7500) );
  XNOR U7892 ( .A(n5548), .B(n7502), .Z(n5609) );
  XNOR U7893 ( .A(n7503), .B(n7504), .Z(n7502) );
  NANDN U7894 ( .A(n6600), .B(n7505), .Z(n7504) );
  XOR U7895 ( .A(n6596), .B(n7506), .Z(n5538) );
  XOR U7896 ( .A(n6593), .B(n7507), .Z(n7506) );
  NANDN U7897 ( .A(n7508), .B(n5559), .Z(n7507) );
  XOR U7898 ( .A(n6595), .B(n5559), .Z(n5612) );
  IV U7899 ( .A(n5503), .Z(n5536) );
  XOR U7900 ( .A(n5604), .B(n5608), .Z(n5503) );
  XOR U7901 ( .A(n5548), .B(n7510), .Z(n5608) );
  XNOR U7902 ( .A(n7499), .B(n7511), .Z(n7510) );
  NANDN U7903 ( .A(n7512), .B(n7513), .Z(n7511) );
  OR U7904 ( .A(n7514), .B(n7515), .Z(n7499) );
  XOR U7905 ( .A(n7516), .B(n7503), .Z(n5548) );
  NANDN U7906 ( .A(n7517), .B(n7518), .Z(n7503) );
  ANDN U7907 ( .B(n7519), .A(n7520), .Z(n7516) );
  XNOR U7908 ( .A(n6596), .B(n7521), .Z(n5604) );
  XOR U7909 ( .A(n7522), .B(n5551), .Z(n7521) );
  OR U7910 ( .A(n7523), .B(n7514), .Z(n5551) );
  XNOR U7911 ( .A(n5554), .B(n7513), .Z(n7514) );
  ANDN U7912 ( .B(n7524), .A(n7525), .Z(n7522) );
  XOR U7913 ( .A(n7526), .B(n6598), .Z(n6596) );
  OR U7914 ( .A(n7517), .B(n7527), .Z(n6598) );
  XNOR U7915 ( .A(n7520), .B(n6600), .Z(n7517) );
  XNOR U7916 ( .A(n7513), .B(n5559), .Z(n6600) );
  XOR U7917 ( .A(n7528), .B(n7529), .Z(n5559) );
  NANDN U7918 ( .A(n7530), .B(n7531), .Z(n7529) );
  IV U7919 ( .A(n7525), .Z(n7513) );
  XNOR U7920 ( .A(n7532), .B(n7533), .Z(n7525) );
  NANDN U7921 ( .A(n7530), .B(n7534), .Z(n7533) );
  NOR U7922 ( .A(n7520), .B(n7535), .Z(n7526) );
  XNOR U7923 ( .A(n6595), .B(n5554), .Z(n7520) );
  XNOR U7924 ( .A(n7536), .B(n7532), .Z(n5554) );
  NANDN U7925 ( .A(n7537), .B(n7538), .Z(n7532) );
  XOR U7926 ( .A(n7534), .B(n7539), .Z(n7538) );
  ANDN U7927 ( .B(n7539), .A(n7540), .Z(n7536) );
  XNOR U7928 ( .A(n7541), .B(n7528), .Z(n6595) );
  NANDN U7929 ( .A(n7537), .B(n7542), .Z(n7528) );
  XOR U7930 ( .A(n7543), .B(n7531), .Z(n7542) );
  XNOR U7931 ( .A(n7544), .B(n7545), .Z(n7530) );
  XOR U7932 ( .A(n7546), .B(n7547), .Z(n7545) );
  XNOR U7933 ( .A(n7548), .B(n7549), .Z(n7544) );
  XNOR U7934 ( .A(n7550), .B(n7551), .Z(n7549) );
  ANDN U7935 ( .B(n7543), .A(n7547), .Z(n7550) );
  ANDN U7936 ( .B(n7543), .A(n7540), .Z(n7541) );
  XNOR U7937 ( .A(n7546), .B(n7552), .Z(n7540) );
  XOR U7938 ( .A(n7553), .B(n7551), .Z(n7552) );
  NAND U7939 ( .A(n7554), .B(n7555), .Z(n7551) );
  XNOR U7940 ( .A(n7548), .B(n7531), .Z(n7555) );
  IV U7941 ( .A(n7543), .Z(n7548) );
  XNOR U7942 ( .A(n7534), .B(n7547), .Z(n7554) );
  IV U7943 ( .A(n7539), .Z(n7547) );
  XOR U7944 ( .A(n7556), .B(n7557), .Z(n7539) );
  XNOR U7945 ( .A(n7558), .B(n7559), .Z(n7557) );
  XNOR U7946 ( .A(n7560), .B(n7561), .Z(n7556) );
  ANDN U7947 ( .B(n6594), .A(n7562), .Z(n7560) );
  AND U7948 ( .A(n7531), .B(n7534), .Z(n7553) );
  XNOR U7949 ( .A(n7531), .B(n7534), .Z(n7546) );
  XNOR U7950 ( .A(n7563), .B(n7564), .Z(n7534) );
  XNOR U7951 ( .A(n7565), .B(n7559), .Z(n7564) );
  XOR U7952 ( .A(n7566), .B(n7567), .Z(n7563) );
  XNOR U7953 ( .A(n7568), .B(n7561), .Z(n7567) );
  OR U7954 ( .A(n5613), .B(n7509), .Z(n7561) );
  XNOR U7955 ( .A(n6594), .B(n7569), .Z(n7509) );
  XNOR U7956 ( .A(n7562), .B(n5560), .Z(n5613) );
  ANDN U7957 ( .B(n7570), .A(n7508), .Z(n7568) );
  XNOR U7958 ( .A(n7571), .B(n7572), .Z(n7531) );
  XNOR U7959 ( .A(n7559), .B(n7573), .Z(n7572) );
  XOR U7960 ( .A(n7501), .B(n7566), .Z(n7573) );
  XNOR U7961 ( .A(n6594), .B(n7562), .Z(n7559) );
  XNOR U7962 ( .A(n7574), .B(n7575), .Z(n7571) );
  XNOR U7963 ( .A(n7576), .B(n7577), .Z(n7575) );
  ANDN U7964 ( .B(n7524), .A(n7512), .Z(n7576) );
  XNOR U7965 ( .A(n7578), .B(n7579), .Z(n7543) );
  XNOR U7966 ( .A(n7565), .B(n7580), .Z(n7579) );
  XNOR U7967 ( .A(n7512), .B(n7558), .Z(n7580) );
  XOR U7968 ( .A(n7566), .B(n7581), .Z(n7558) );
  XNOR U7969 ( .A(n7582), .B(n7583), .Z(n7581) );
  NAND U7970 ( .A(n6601), .B(n7505), .Z(n7583) );
  XNOR U7971 ( .A(n7584), .B(n7582), .Z(n7566) );
  NANDN U7972 ( .A(n7527), .B(n7518), .Z(n7582) );
  XOR U7973 ( .A(n7519), .B(n7505), .Z(n7518) );
  XNOR U7974 ( .A(n7585), .B(n5560), .Z(n7505) );
  XOR U7975 ( .A(n7535), .B(n6601), .Z(n7527) );
  XOR U7976 ( .A(n7524), .B(n7569), .Z(n6601) );
  ANDN U7977 ( .B(n7519), .A(n7535), .Z(n7584) );
  XNOR U7978 ( .A(n7574), .B(n6594), .Z(n7535) );
  XNOR U7979 ( .A(n7586), .B(n7587), .Z(n6594) );
  XNOR U7980 ( .A(n7588), .B(n7589), .Z(n7587) );
  XOR U7981 ( .A(n7590), .B(n5614), .Z(n7519) );
  XOR U7982 ( .A(n7569), .B(n7570), .Z(n7565) );
  IV U7983 ( .A(n5560), .Z(n7570) );
  XOR U7984 ( .A(n7591), .B(n7592), .Z(n5560) );
  XNOR U7985 ( .A(n7593), .B(n7589), .Z(n7592) );
  IV U7986 ( .A(n7508), .Z(n7569) );
  XOR U7987 ( .A(n7589), .B(n7594), .Z(n7508) );
  XNOR U7988 ( .A(n7524), .B(n7595), .Z(n7578) );
  XNOR U7989 ( .A(n7596), .B(n7577), .Z(n7595) );
  OR U7990 ( .A(n7515), .B(n7523), .Z(n7577) );
  XNOR U7991 ( .A(n7574), .B(n7524), .Z(n7523) );
  XOR U7992 ( .A(n7501), .B(n7585), .Z(n7515) );
  IV U7993 ( .A(n7512), .Z(n7585) );
  XOR U7994 ( .A(n5614), .B(n7597), .Z(n7512) );
  XNOR U7995 ( .A(n7593), .B(n7586), .Z(n7597) );
  XOR U7996 ( .A(n7598), .B(n7599), .Z(n7586) );
  XOR U7997 ( .A(n2822), .B(n2817), .Z(n7599) );
  XOR U7998 ( .A(n3803), .B(n7600), .Z(n7598) );
  XNOR U7999 ( .A(key[1082]), .B(n5084), .Z(n7600) );
  XOR U8000 ( .A(n7601), .B(n7602), .Z(n5084) );
  XNOR U8001 ( .A(n7603), .B(n7604), .Z(n7601) );
  XNOR U8002 ( .A(n2821), .B(n2778), .Z(n3803) );
  IV U8003 ( .A(n7562), .Z(n5614) );
  XOR U8004 ( .A(n7591), .B(n7605), .Z(n7562) );
  XOR U8005 ( .A(n7589), .B(n7606), .Z(n7605) );
  ANDN U8006 ( .B(n7590), .A(n5553), .Z(n7596) );
  IV U8007 ( .A(n7501), .Z(n7590) );
  XOR U8008 ( .A(n7591), .B(n7607), .Z(n7501) );
  XOR U8009 ( .A(n7589), .B(n7608), .Z(n7607) );
  XOR U8010 ( .A(n7609), .B(n7610), .Z(n7589) );
  XOR U8011 ( .A(n5087), .B(n5553), .Z(n7610) );
  IV U8012 ( .A(n7574), .Z(n5553) );
  XNOR U8013 ( .A(n3777), .B(n5078), .Z(n5087) );
  XNOR U8014 ( .A(n3810), .B(n3785), .Z(n5078) );
  XOR U8015 ( .A(n7611), .B(n7612), .Z(n3785) );
  XOR U8016 ( .A(n7613), .B(n7614), .Z(n7612) );
  XOR U8017 ( .A(n7615), .B(n7616), .Z(n7611) );
  IV U8018 ( .A(n7617), .Z(n3810) );
  XNOR U8019 ( .A(n2797), .B(n2790), .Z(n3777) );
  XNOR U8020 ( .A(n7618), .B(n7619), .Z(n2797) );
  XOR U8021 ( .A(n3771), .B(n7620), .Z(n7609) );
  XNOR U8022 ( .A(key[1086]), .B(n2799), .Z(n7620) );
  XOR U8023 ( .A(n7621), .B(n7622), .Z(n2799) );
  XNOR U8024 ( .A(n3789), .B(n2804), .Z(n3771) );
  IV U8025 ( .A(n7594), .Z(n7591) );
  XOR U8026 ( .A(n7623), .B(n7624), .Z(n7594) );
  XOR U8027 ( .A(n2790), .B(n5074), .Z(n7624) );
  XNOR U8028 ( .A(n3780), .B(n2795), .Z(n5074) );
  XOR U8029 ( .A(n7625), .B(n7626), .Z(n3780) );
  XNOR U8030 ( .A(n7627), .B(n7628), .Z(n7626) );
  XNOR U8031 ( .A(n7629), .B(n7630), .Z(n7625) );
  XOR U8032 ( .A(n7631), .B(n7632), .Z(n7630) );
  ANDN U8033 ( .B(n7633), .A(n7634), .Z(n7632) );
  XOR U8034 ( .A(n3778), .B(n7637), .Z(n7623) );
  XNOR U8035 ( .A(key[1085]), .B(n5075), .Z(n7637) );
  XNOR U8036 ( .A(n7604), .B(n7638), .Z(n5075) );
  XNOR U8037 ( .A(n7639), .B(n7640), .Z(n7604) );
  XNOR U8038 ( .A(n7641), .B(n7642), .Z(n7640) );
  ANDN U8039 ( .B(n7643), .A(n7644), .Z(n7641) );
  XNOR U8040 ( .A(n7645), .B(n7646), .Z(n3778) );
  XNOR U8041 ( .A(n7647), .B(n7648), .Z(n7646) );
  XNOR U8042 ( .A(n7649), .B(n7650), .Z(n7645) );
  XOR U8043 ( .A(n7651), .B(n7652), .Z(n7650) );
  ANDN U8044 ( .B(n7653), .A(n7654), .Z(n7652) );
  XOR U8045 ( .A(n7655), .B(n7656), .Z(n7524) );
  XNOR U8046 ( .A(n7608), .B(n7606), .Z(n7656) );
  XNOR U8047 ( .A(n7657), .B(n7658), .Z(n7606) );
  XOR U8048 ( .A(n5079), .B(n2832), .Z(n7658) );
  XOR U8049 ( .A(n7617), .B(n7659), .Z(n2832) );
  XOR U8050 ( .A(n3788), .B(n2804), .Z(n5079) );
  XNOR U8051 ( .A(n7660), .B(n7661), .Z(n2804) );
  XOR U8052 ( .A(n7636), .B(n7662), .Z(n7661) );
  XOR U8053 ( .A(n7663), .B(n7664), .Z(n7660) );
  XOR U8054 ( .A(n7665), .B(n7666), .Z(n3788) );
  XNOR U8055 ( .A(n7618), .B(n7628), .Z(n7666) );
  XNOR U8056 ( .A(n7667), .B(n7668), .Z(n7628) );
  XNOR U8057 ( .A(n7669), .B(n7670), .Z(n7668) );
  OR U8058 ( .A(n7671), .B(n7672), .Z(n7670) );
  XOR U8059 ( .A(key[1087]), .B(n3786), .Z(n7657) );
  XNOR U8060 ( .A(n7673), .B(n7674), .Z(n3786) );
  XOR U8061 ( .A(n7675), .B(n7648), .Z(n7674) );
  XNOR U8062 ( .A(n7676), .B(n7677), .Z(n7648) );
  XNOR U8063 ( .A(n7678), .B(n7679), .Z(n7677) );
  NANDN U8064 ( .A(n7680), .B(n7681), .Z(n7679) );
  XOR U8065 ( .A(n7682), .B(n7683), .Z(n7673) );
  XNOR U8066 ( .A(n7684), .B(n5065), .Z(n7608) );
  XOR U8067 ( .A(n7685), .B(n7686), .Z(n5065) );
  XOR U8068 ( .A(n3796), .B(n2813), .Z(n7686) );
  XOR U8069 ( .A(n7627), .B(n2821), .Z(n3796) );
  XNOR U8070 ( .A(n7687), .B(n7688), .Z(n2821) );
  XNOR U8071 ( .A(n7617), .B(n3779), .Z(n7685) );
  XNOR U8072 ( .A(n7689), .B(n7690), .Z(n3779) );
  XNOR U8073 ( .A(n7691), .B(n7614), .Z(n7690) );
  XNOR U8074 ( .A(n7692), .B(n7693), .Z(n7614) );
  XNOR U8075 ( .A(n7694), .B(n7695), .Z(n7693) );
  NANDN U8076 ( .A(n7696), .B(n7697), .Z(n7695) );
  XNOR U8077 ( .A(n7698), .B(n7699), .Z(n7689) );
  XOR U8078 ( .A(n7642), .B(n7700), .Z(n7699) );
  ANDN U8079 ( .B(n7701), .A(n7702), .Z(n7700) );
  ANDN U8080 ( .B(n7703), .A(n7704), .Z(n7642) );
  XNOR U8081 ( .A(n3792), .B(n7705), .Z(n7684) );
  XOR U8082 ( .A(key[1084]), .B(n3794), .Z(n7705) );
  XOR U8083 ( .A(n7649), .B(n2822), .Z(n3794) );
  XOR U8084 ( .A(n7706), .B(n7682), .Z(n2822) );
  XNOR U8085 ( .A(n7659), .B(n2795), .Z(n3792) );
  XNOR U8086 ( .A(n7707), .B(n7708), .Z(n2795) );
  XOR U8087 ( .A(n7709), .B(n7662), .Z(n7708) );
  XNOR U8088 ( .A(n7710), .B(n7711), .Z(n7662) );
  XNOR U8089 ( .A(n7712), .B(n7713), .Z(n7711) );
  OR U8090 ( .A(n7714), .B(n7715), .Z(n7713) );
  XNOR U8091 ( .A(n7716), .B(n7717), .Z(n7707) );
  XNOR U8092 ( .A(n7718), .B(n7719), .Z(n7717) );
  ANDN U8093 ( .B(n7720), .A(n7721), .Z(n7719) );
  XOR U8094 ( .A(n7574), .B(n7588), .Z(n7655) );
  XOR U8095 ( .A(n7722), .B(n7723), .Z(n7588) );
  XNOR U8096 ( .A(n7593), .B(n7724), .Z(n7723) );
  XNOR U8097 ( .A(n5098), .B(n5092), .Z(n7724) );
  XNOR U8098 ( .A(n7617), .B(n3793), .Z(n5092) );
  IV U8099 ( .A(n5067), .Z(n3793) );
  XOR U8100 ( .A(n7698), .B(n5096), .Z(n5067) );
  IV U8101 ( .A(n5083), .Z(n5096) );
  XOR U8102 ( .A(n7698), .B(n7725), .Z(n7617) );
  XNOR U8103 ( .A(n7692), .B(n7726), .Z(n7698) );
  XNOR U8104 ( .A(n7727), .B(n7728), .Z(n7726) );
  ANDN U8105 ( .B(n7729), .A(n7644), .Z(n7727) );
  IV U8106 ( .A(n7730), .Z(n7644) );
  XNOR U8107 ( .A(n7731), .B(n7732), .Z(n7692) );
  XNOR U8108 ( .A(n7733), .B(n7734), .Z(n7732) );
  NANDN U8109 ( .A(n7735), .B(n7736), .Z(n7734) );
  XNOR U8110 ( .A(n2780), .B(n2817), .Z(n5098) );
  XNOR U8111 ( .A(n7737), .B(n7738), .Z(n2817) );
  XOR U8112 ( .A(n7739), .B(n7635), .Z(n7738) );
  XOR U8113 ( .A(n7740), .B(n7741), .Z(n7635) );
  XOR U8114 ( .A(n7742), .B(n7718), .Z(n7741) );
  NANDN U8115 ( .A(n7743), .B(n7744), .Z(n7718) );
  ANDN U8116 ( .B(n7745), .A(n7746), .Z(n7742) );
  XNOR U8117 ( .A(n7747), .B(n7664), .Z(n7737) );
  XOR U8118 ( .A(n7665), .B(n7748), .Z(n2780) );
  XNOR U8119 ( .A(n7749), .B(n7619), .Z(n7748) );
  XNOR U8120 ( .A(n7750), .B(n7751), .Z(n7619) );
  XNOR U8121 ( .A(n7752), .B(n7631), .Z(n7751) );
  ANDN U8122 ( .B(n7753), .A(n7754), .Z(n7631) );
  ANDN U8123 ( .B(n7755), .A(n7756), .Z(n7752) );
  XNOR U8124 ( .A(n7687), .B(n7757), .Z(n7665) );
  XOR U8125 ( .A(n7758), .B(n7759), .Z(n7593) );
  XNOR U8126 ( .A(n2778), .B(n5083), .Z(n7759) );
  XNOR U8127 ( .A(n7725), .B(n7615), .Z(n5083) );
  XOR U8128 ( .A(n2831), .B(n7760), .Z(n7758) );
  XNOR U8129 ( .A(key[1081]), .B(n3808), .Z(n7760) );
  XNOR U8130 ( .A(n2825), .B(n2835), .Z(n3808) );
  XOR U8131 ( .A(n7618), .B(n7761), .Z(n2835) );
  XOR U8132 ( .A(n7687), .B(n7757), .Z(n7761) );
  XOR U8133 ( .A(n7750), .B(n7762), .Z(n7757) );
  XNOR U8134 ( .A(n7763), .B(n7764), .Z(n7762) );
  NANDN U8135 ( .A(n7671), .B(n7765), .Z(n7764) );
  XNOR U8136 ( .A(n7629), .B(n7766), .Z(n7750) );
  XNOR U8137 ( .A(n7767), .B(n7768), .Z(n7766) );
  NAND U8138 ( .A(n7769), .B(n7770), .Z(n7768) );
  XNOR U8139 ( .A(n7771), .B(n7772), .Z(n7687) );
  XNOR U8140 ( .A(n7773), .B(n7774), .Z(n7772) );
  NAND U8141 ( .A(n7775), .B(n7633), .Z(n7774) );
  XOR U8142 ( .A(n7776), .B(n7749), .Z(n7618) );
  XNOR U8143 ( .A(n7629), .B(n7777), .Z(n7749) );
  XNOR U8144 ( .A(n7763), .B(n7778), .Z(n7777) );
  NANDN U8145 ( .A(n7779), .B(n7780), .Z(n7778) );
  OR U8146 ( .A(n7781), .B(n7782), .Z(n7763) );
  XOR U8147 ( .A(n7783), .B(n7767), .Z(n7629) );
  NANDN U8148 ( .A(n7784), .B(n7785), .Z(n7767) );
  ANDN U8149 ( .B(n7786), .A(n7787), .Z(n7783) );
  IV U8150 ( .A(n7788), .Z(n2825) );
  XNOR U8151 ( .A(n7675), .B(n7789), .Z(n2831) );
  IV U8152 ( .A(n7622), .Z(n7675) );
  XOR U8153 ( .A(n7706), .B(n7790), .Z(n7622) );
  XNOR U8154 ( .A(n3799), .B(n7791), .Z(n7722) );
  XNOR U8155 ( .A(key[1083]), .B(n2782), .Z(n7791) );
  XOR U8156 ( .A(n7792), .B(n7789), .Z(n2782) );
  XNOR U8157 ( .A(n7682), .B(n7683), .Z(n7789) );
  XOR U8158 ( .A(n7793), .B(n7794), .Z(n7683) );
  XNOR U8159 ( .A(n7795), .B(n7796), .Z(n7794) );
  NANDN U8160 ( .A(n7797), .B(n7681), .Z(n7796) );
  XOR U8161 ( .A(n7798), .B(n7799), .Z(n7682) );
  XOR U8162 ( .A(n7800), .B(n7801), .Z(n7799) );
  NANDN U8163 ( .A(n7802), .B(n7653), .Z(n7801) );
  XOR U8164 ( .A(n7621), .B(n7790), .Z(n7792) );
  XOR U8165 ( .A(n7647), .B(n7803), .Z(n7790) );
  XNOR U8166 ( .A(n7795), .B(n7804), .Z(n7803) );
  NANDN U8167 ( .A(n7805), .B(n7806), .Z(n7804) );
  OR U8168 ( .A(n7807), .B(n7808), .Z(n7795) );
  XNOR U8169 ( .A(n7810), .B(n7651), .Z(n7809) );
  ANDN U8170 ( .B(n7811), .A(n7812), .Z(n7651) );
  ANDN U8171 ( .B(n7813), .A(n7814), .Z(n7810) );
  XNOR U8172 ( .A(n7647), .B(n7815), .Z(n7793) );
  XNOR U8173 ( .A(n7816), .B(n7817), .Z(n7815) );
  NANDN U8174 ( .A(n7818), .B(n7819), .Z(n7817) );
  XOR U8175 ( .A(n7820), .B(n7816), .Z(n7647) );
  NANDN U8176 ( .A(n7821), .B(n7822), .Z(n7816) );
  ANDN U8177 ( .B(n7823), .A(n7824), .Z(n7820) );
  XOR U8178 ( .A(n3789), .B(n2813), .Z(n3799) );
  XOR U8179 ( .A(n2778), .B(n7709), .Z(n2813) );
  XOR U8180 ( .A(n7663), .B(n7825), .Z(n2778) );
  XOR U8181 ( .A(n7826), .B(n7827), .Z(n7574) );
  XOR U8182 ( .A(n5101), .B(n3789), .Z(n7827) );
  IV U8183 ( .A(n7659), .Z(n3789) );
  XOR U8184 ( .A(n7825), .B(n7709), .Z(n7659) );
  XOR U8185 ( .A(n7710), .B(n7828), .Z(n7709) );
  XOR U8186 ( .A(n7829), .B(n7830), .Z(n7828) );
  ANDN U8187 ( .B(n7745), .A(n7831), .Z(n7829) );
  XNOR U8188 ( .A(n7832), .B(n7833), .Z(n7710) );
  XNOR U8189 ( .A(n7834), .B(n7835), .Z(n7833) );
  NAND U8190 ( .A(n7836), .B(n7837), .Z(n7835) );
  IV U8191 ( .A(n5095), .Z(n5101) );
  XOR U8192 ( .A(n7613), .B(n7602), .Z(n5095) );
  XNOR U8193 ( .A(n7615), .B(n7616), .Z(n7602) );
  XOR U8194 ( .A(n7639), .B(n7838), .Z(n7616) );
  XNOR U8195 ( .A(n7839), .B(n7840), .Z(n7838) );
  NANDN U8196 ( .A(n7841), .B(n7697), .Z(n7840) );
  XNOR U8197 ( .A(n7691), .B(n7842), .Z(n7639) );
  XNOR U8198 ( .A(n7843), .B(n7844), .Z(n7842) );
  NANDN U8199 ( .A(n7735), .B(n7845), .Z(n7844) );
  XOR U8200 ( .A(n7731), .B(n7846), .Z(n7615) );
  XOR U8201 ( .A(n7728), .B(n7847), .Z(n7846) );
  NANDN U8202 ( .A(n7848), .B(n7701), .Z(n7847) );
  XOR U8203 ( .A(n7730), .B(n7701), .Z(n7703) );
  IV U8204 ( .A(n7638), .Z(n7613) );
  XOR U8205 ( .A(n7725), .B(n7603), .Z(n7638) );
  XOR U8206 ( .A(n7691), .B(n7850), .Z(n7603) );
  XNOR U8207 ( .A(n7839), .B(n7851), .Z(n7850) );
  NANDN U8208 ( .A(n7852), .B(n7853), .Z(n7851) );
  OR U8209 ( .A(n7854), .B(n7855), .Z(n7839) );
  XOR U8210 ( .A(n7856), .B(n7843), .Z(n7691) );
  NANDN U8211 ( .A(n7857), .B(n7858), .Z(n7843) );
  ANDN U8212 ( .B(n7859), .A(n7860), .Z(n7856) );
  XNOR U8213 ( .A(n7731), .B(n7861), .Z(n7725) );
  XOR U8214 ( .A(n7862), .B(n7694), .Z(n7861) );
  OR U8215 ( .A(n7863), .B(n7854), .Z(n7694) );
  XNOR U8216 ( .A(n7697), .B(n7853), .Z(n7854) );
  ANDN U8217 ( .B(n7864), .A(n7865), .Z(n7862) );
  XOR U8218 ( .A(n7866), .B(n7733), .Z(n7731) );
  OR U8219 ( .A(n7857), .B(n7867), .Z(n7733) );
  XNOR U8220 ( .A(n7860), .B(n7735), .Z(n7857) );
  XNOR U8221 ( .A(n7853), .B(n7701), .Z(n7735) );
  XOR U8222 ( .A(n7868), .B(n7869), .Z(n7701) );
  NANDN U8223 ( .A(n7870), .B(n7871), .Z(n7869) );
  IV U8224 ( .A(n7865), .Z(n7853) );
  XNOR U8225 ( .A(n7872), .B(n7873), .Z(n7865) );
  NANDN U8226 ( .A(n7870), .B(n7874), .Z(n7873) );
  NOR U8227 ( .A(n7860), .B(n7875), .Z(n7866) );
  XNOR U8228 ( .A(n7730), .B(n7697), .Z(n7860) );
  XNOR U8229 ( .A(n7876), .B(n7872), .Z(n7697) );
  NANDN U8230 ( .A(n7877), .B(n7878), .Z(n7872) );
  XOR U8231 ( .A(n7874), .B(n7879), .Z(n7878) );
  ANDN U8232 ( .B(n7879), .A(n7880), .Z(n7876) );
  XNOR U8233 ( .A(n7881), .B(n7868), .Z(n7730) );
  NANDN U8234 ( .A(n7877), .B(n7882), .Z(n7868) );
  XOR U8235 ( .A(n7883), .B(n7871), .Z(n7882) );
  XNOR U8236 ( .A(n7884), .B(n7885), .Z(n7870) );
  XOR U8237 ( .A(n7886), .B(n7887), .Z(n7885) );
  XNOR U8238 ( .A(n7888), .B(n7889), .Z(n7884) );
  XNOR U8239 ( .A(n7890), .B(n7891), .Z(n7889) );
  ANDN U8240 ( .B(n7883), .A(n7887), .Z(n7890) );
  ANDN U8241 ( .B(n7883), .A(n7880), .Z(n7881) );
  XNOR U8242 ( .A(n7886), .B(n7892), .Z(n7880) );
  XOR U8243 ( .A(n7893), .B(n7891), .Z(n7892) );
  NAND U8244 ( .A(n7894), .B(n7895), .Z(n7891) );
  XNOR U8245 ( .A(n7888), .B(n7871), .Z(n7895) );
  IV U8246 ( .A(n7883), .Z(n7888) );
  XNOR U8247 ( .A(n7874), .B(n7887), .Z(n7894) );
  IV U8248 ( .A(n7879), .Z(n7887) );
  XOR U8249 ( .A(n7896), .B(n7897), .Z(n7879) );
  XNOR U8250 ( .A(n7898), .B(n7899), .Z(n7897) );
  XNOR U8251 ( .A(n7900), .B(n7901), .Z(n7896) );
  ANDN U8252 ( .B(n7729), .A(n7902), .Z(n7900) );
  AND U8253 ( .A(n7871), .B(n7874), .Z(n7893) );
  XNOR U8254 ( .A(n7871), .B(n7874), .Z(n7886) );
  XNOR U8255 ( .A(n7903), .B(n7904), .Z(n7874) );
  XNOR U8256 ( .A(n7905), .B(n7899), .Z(n7904) );
  XOR U8257 ( .A(n7906), .B(n7907), .Z(n7903) );
  XNOR U8258 ( .A(n7908), .B(n7901), .Z(n7907) );
  OR U8259 ( .A(n7704), .B(n7849), .Z(n7901) );
  XNOR U8260 ( .A(n7729), .B(n7909), .Z(n7849) );
  XNOR U8261 ( .A(n7902), .B(n7702), .Z(n7704) );
  ANDN U8262 ( .B(n7910), .A(n7848), .Z(n7908) );
  XNOR U8263 ( .A(n7911), .B(n7912), .Z(n7871) );
  XNOR U8264 ( .A(n7899), .B(n7913), .Z(n7912) );
  XOR U8265 ( .A(n7841), .B(n7906), .Z(n7913) );
  XNOR U8266 ( .A(n7729), .B(n7902), .Z(n7899) );
  XNOR U8267 ( .A(n7914), .B(n7915), .Z(n7911) );
  XNOR U8268 ( .A(n7916), .B(n7917), .Z(n7915) );
  ANDN U8269 ( .B(n7864), .A(n7852), .Z(n7916) );
  XNOR U8270 ( .A(n7918), .B(n7919), .Z(n7883) );
  XNOR U8271 ( .A(n7905), .B(n7920), .Z(n7919) );
  XNOR U8272 ( .A(n7852), .B(n7898), .Z(n7920) );
  XOR U8273 ( .A(n7906), .B(n7921), .Z(n7898) );
  XNOR U8274 ( .A(n7922), .B(n7923), .Z(n7921) );
  NAND U8275 ( .A(n7736), .B(n7845), .Z(n7923) );
  XNOR U8276 ( .A(n7924), .B(n7922), .Z(n7906) );
  NANDN U8277 ( .A(n7867), .B(n7858), .Z(n7922) );
  XOR U8278 ( .A(n7859), .B(n7845), .Z(n7858) );
  XNOR U8279 ( .A(n7925), .B(n7702), .Z(n7845) );
  XOR U8280 ( .A(n7875), .B(n7736), .Z(n7867) );
  XOR U8281 ( .A(n7864), .B(n7909), .Z(n7736) );
  ANDN U8282 ( .B(n7859), .A(n7875), .Z(n7924) );
  XNOR U8283 ( .A(n7914), .B(n7729), .Z(n7875) );
  XNOR U8284 ( .A(n7926), .B(n7927), .Z(n7729) );
  XNOR U8285 ( .A(n7928), .B(n7929), .Z(n7927) );
  XOR U8286 ( .A(n7930), .B(n7643), .Z(n7859) );
  XOR U8287 ( .A(n7909), .B(n7910), .Z(n7905) );
  IV U8288 ( .A(n7702), .Z(n7910) );
  XOR U8289 ( .A(n7931), .B(n7932), .Z(n7702) );
  XNOR U8290 ( .A(n7933), .B(n7929), .Z(n7932) );
  IV U8291 ( .A(n7848), .Z(n7909) );
  XOR U8292 ( .A(n7929), .B(n7934), .Z(n7848) );
  XNOR U8293 ( .A(n7864), .B(n7935), .Z(n7918) );
  XNOR U8294 ( .A(n7936), .B(n7917), .Z(n7935) );
  OR U8295 ( .A(n7855), .B(n7863), .Z(n7917) );
  XNOR U8296 ( .A(n7914), .B(n7864), .Z(n7863) );
  XOR U8297 ( .A(n7841), .B(n7925), .Z(n7855) );
  IV U8298 ( .A(n7852), .Z(n7925) );
  XOR U8299 ( .A(n7643), .B(n7937), .Z(n7852) );
  XNOR U8300 ( .A(n7933), .B(n7926), .Z(n7937) );
  XOR U8301 ( .A(n7938), .B(n7939), .Z(n7926) );
  XNOR U8302 ( .A(n7940), .B(n7941), .Z(n7939) );
  XOR U8303 ( .A(n6585), .B(n7942), .Z(n7938) );
  XOR U8304 ( .A(key[954]), .B(n6545), .Z(n7942) );
  XOR U8305 ( .A(n7321), .B(n7943), .Z(n6545) );
  IV U8306 ( .A(n7902), .Z(n7643) );
  XOR U8307 ( .A(n7931), .B(n7944), .Z(n7902) );
  XOR U8308 ( .A(n7929), .B(n7945), .Z(n7944) );
  ANDN U8309 ( .B(n7930), .A(n7696), .Z(n7936) );
  IV U8310 ( .A(n7841), .Z(n7930) );
  XOR U8311 ( .A(n7931), .B(n7946), .Z(n7841) );
  XOR U8312 ( .A(n7929), .B(n7947), .Z(n7946) );
  XOR U8313 ( .A(n7948), .B(n7949), .Z(n7929) );
  XNOR U8314 ( .A(n6552), .B(n7696), .Z(n7949) );
  IV U8315 ( .A(n7914), .Z(n7696) );
  XNOR U8316 ( .A(n7335), .B(n6565), .Z(n6552) );
  XOR U8317 ( .A(n7365), .B(n7950), .Z(n6565) );
  XNOR U8318 ( .A(n7330), .B(n7951), .Z(n7335) );
  XOR U8319 ( .A(n7329), .B(n7952), .Z(n7948) );
  XNOR U8320 ( .A(key[958]), .B(n7953), .Z(n7952) );
  XOR U8321 ( .A(n7954), .B(n7955), .Z(n7329) );
  IV U8322 ( .A(n7934), .Z(n7931) );
  XOR U8323 ( .A(n7956), .B(n7957), .Z(n7934) );
  XOR U8324 ( .A(n7951), .B(n6559), .Z(n7957) );
  XOR U8325 ( .A(n7336), .B(n7958), .Z(n6559) );
  XNOR U8326 ( .A(n7959), .B(n7960), .Z(n7956) );
  XOR U8327 ( .A(key[957]), .B(n7961), .Z(n7960) );
  XOR U8328 ( .A(n7962), .B(n7963), .Z(n7864) );
  XNOR U8329 ( .A(n7947), .B(n7945), .Z(n7963) );
  XNOR U8330 ( .A(n7964), .B(n7965), .Z(n7945) );
  XNOR U8331 ( .A(n6589), .B(n6566), .Z(n7965) );
  XOR U8332 ( .A(n7966), .B(n7955), .Z(n6566) );
  XOR U8333 ( .A(key[959]), .B(n7967), .Z(n7964) );
  XNOR U8334 ( .A(n7968), .B(n6569), .Z(n7947) );
  XOR U8335 ( .A(n7969), .B(n7970), .Z(n6569) );
  XOR U8336 ( .A(n7350), .B(n7971), .Z(n7970) );
  XNOR U8337 ( .A(n7365), .B(n6558), .Z(n7969) );
  XOR U8338 ( .A(n7347), .B(n7972), .Z(n7968) );
  XNOR U8339 ( .A(key[956]), .B(n7973), .Z(n7972) );
  XOR U8340 ( .A(n7954), .B(n7958), .Z(n7347) );
  XOR U8341 ( .A(n7914), .B(n7928), .Z(n7962) );
  XOR U8342 ( .A(n7974), .B(n7975), .Z(n7928) );
  XNOR U8343 ( .A(n7933), .B(n7976), .Z(n7975) );
  XOR U8344 ( .A(n6583), .B(n6575), .Z(n7976) );
  XOR U8345 ( .A(n7365), .B(n6572), .Z(n6575) );
  XNOR U8346 ( .A(n7359), .B(n7941), .Z(n6583) );
  XOR U8347 ( .A(n7977), .B(n7978), .Z(n7933) );
  XNOR U8348 ( .A(n7979), .B(n6544), .Z(n7978) );
  XNOR U8349 ( .A(n7980), .B(n7981), .Z(n7977) );
  XOR U8350 ( .A(key[953]), .B(n6582), .Z(n7981) );
  XOR U8351 ( .A(n7358), .B(n7982), .Z(n6582) );
  XNOR U8352 ( .A(n7353), .B(n7983), .Z(n7974) );
  XNOR U8353 ( .A(key[955]), .B(n7984), .Z(n7983) );
  XNOR U8354 ( .A(n7343), .B(n7971), .Z(n7353) );
  XOR U8355 ( .A(n7985), .B(n7986), .Z(n7914) );
  XOR U8356 ( .A(n7987), .B(n7343), .Z(n7986) );
  IV U8357 ( .A(n7954), .Z(n7343) );
  XNOR U8358 ( .A(n7982), .B(n7988), .Z(n7985) );
  XNOR U8359 ( .A(key[952]), .B(n7364), .Z(n7988) );
  XNOR U8360 ( .A(n3809), .B(n7989), .Z(n7826) );
  XNOR U8361 ( .A(key[1080]), .B(n7788), .Z(n7989) );
  XOR U8362 ( .A(n7636), .B(n7990), .Z(n7788) );
  XOR U8363 ( .A(n7747), .B(n7664), .Z(n7990) );
  XOR U8364 ( .A(n7740), .B(n7991), .Z(n7664) );
  XNOR U8365 ( .A(n7992), .B(n7993), .Z(n7991) );
  NANDN U8366 ( .A(n7714), .B(n7994), .Z(n7993) );
  XNOR U8367 ( .A(n7716), .B(n7995), .Z(n7740) );
  XNOR U8368 ( .A(n7996), .B(n7997), .Z(n7995) );
  NAND U8369 ( .A(n7998), .B(n7836), .Z(n7997) );
  IV U8370 ( .A(n7663), .Z(n7747) );
  XOR U8371 ( .A(n7832), .B(n7999), .Z(n7663) );
  XNOR U8372 ( .A(n7830), .B(n8000), .Z(n7999) );
  NAND U8373 ( .A(n8001), .B(n7720), .Z(n8000) );
  NANDN U8374 ( .A(n8002), .B(n7744), .Z(n7830) );
  XOR U8375 ( .A(n7745), .B(n7720), .Z(n7744) );
  XNOR U8376 ( .A(n7739), .B(n7825), .Z(n7636) );
  XOR U8377 ( .A(n7832), .B(n8003), .Z(n7825) );
  XOR U8378 ( .A(n8004), .B(n7712), .Z(n8003) );
  OR U8379 ( .A(n8005), .B(n8006), .Z(n7712) );
  NOR U8380 ( .A(n8007), .B(n8008), .Z(n8004) );
  XOR U8381 ( .A(n8009), .B(n7834), .Z(n7832) );
  OR U8382 ( .A(n8010), .B(n8011), .Z(n7834) );
  ANDN U8383 ( .B(n8012), .A(n8013), .Z(n8009) );
  XNOR U8384 ( .A(n7716), .B(n8014), .Z(n7739) );
  XNOR U8385 ( .A(n7992), .B(n8015), .Z(n8014) );
  NANDN U8386 ( .A(n8008), .B(n8016), .Z(n8015) );
  OR U8387 ( .A(n8005), .B(n8017), .Z(n7992) );
  XNOR U8388 ( .A(n7714), .B(n8008), .Z(n8005) );
  XOR U8389 ( .A(n8018), .B(n7996), .Z(n7716) );
  NANDN U8390 ( .A(n8010), .B(n8019), .Z(n7996) );
  XOR U8391 ( .A(n8013), .B(n7836), .Z(n8010) );
  XNOR U8392 ( .A(n8008), .B(n7720), .Z(n7836) );
  XOR U8393 ( .A(n8020), .B(n8021), .Z(n7720) );
  NANDN U8394 ( .A(n8022), .B(n8023), .Z(n8021) );
  XNOR U8395 ( .A(n8024), .B(n8025), .Z(n8008) );
  OR U8396 ( .A(n8022), .B(n8026), .Z(n8025) );
  ANDN U8397 ( .B(n8027), .A(n8013), .Z(n8018) );
  XOR U8398 ( .A(n7714), .B(n7745), .Z(n8013) );
  XNOR U8399 ( .A(n8028), .B(n8020), .Z(n7745) );
  NANDN U8400 ( .A(n8029), .B(n8030), .Z(n8020) );
  ANDN U8401 ( .B(n8031), .A(n8032), .Z(n8028) );
  NANDN U8402 ( .A(n8029), .B(n8034), .Z(n8024) );
  XOR U8403 ( .A(n8035), .B(n8022), .Z(n8029) );
  XNOR U8404 ( .A(n8036), .B(n8037), .Z(n8022) );
  XOR U8405 ( .A(n8038), .B(n8031), .Z(n8037) );
  XNOR U8406 ( .A(n8039), .B(n8040), .Z(n8036) );
  XNOR U8407 ( .A(n8041), .B(n8042), .Z(n8040) );
  ANDN U8408 ( .B(n8031), .A(n8043), .Z(n8041) );
  IV U8409 ( .A(n8044), .Z(n8031) );
  ANDN U8410 ( .B(n8035), .A(n8043), .Z(n8033) );
  IV U8411 ( .A(n8039), .Z(n8043) );
  IV U8412 ( .A(n8032), .Z(n8035) );
  XNOR U8413 ( .A(n8038), .B(n8045), .Z(n8032) );
  XOR U8414 ( .A(n8046), .B(n8042), .Z(n8045) );
  NAND U8415 ( .A(n8034), .B(n8030), .Z(n8042) );
  XNOR U8416 ( .A(n8023), .B(n8044), .Z(n8030) );
  XOR U8417 ( .A(n8047), .B(n8048), .Z(n8044) );
  XOR U8418 ( .A(n8049), .B(n8050), .Z(n8048) );
  XNOR U8419 ( .A(n8016), .B(n8051), .Z(n8050) );
  XNOR U8420 ( .A(n8052), .B(n8053), .Z(n8047) );
  XNOR U8421 ( .A(n8054), .B(n8055), .Z(n8053) );
  ANDN U8422 ( .B(n7994), .A(n7715), .Z(n8054) );
  XNOR U8423 ( .A(n8039), .B(n8026), .Z(n8034) );
  XOR U8424 ( .A(n8056), .B(n8057), .Z(n8039) );
  XNOR U8425 ( .A(n8058), .B(n8051), .Z(n8057) );
  XOR U8426 ( .A(n8059), .B(n8060), .Z(n8051) );
  XNOR U8427 ( .A(n8061), .B(n8062), .Z(n8060) );
  NAND U8428 ( .A(n7837), .B(n7998), .Z(n8062) );
  XNOR U8429 ( .A(n8063), .B(n8064), .Z(n8056) );
  ANDN U8430 ( .B(n8065), .A(n7831), .Z(n8063) );
  ANDN U8431 ( .B(n8023), .A(n8026), .Z(n8046) );
  XOR U8432 ( .A(n8026), .B(n8023), .Z(n8038) );
  XNOR U8433 ( .A(n8066), .B(n8067), .Z(n8023) );
  XNOR U8434 ( .A(n8059), .B(n8068), .Z(n8067) );
  XNOR U8435 ( .A(n8058), .B(n7994), .Z(n8068) );
  XNOR U8436 ( .A(n8069), .B(n8070), .Z(n8066) );
  XNOR U8437 ( .A(n8071), .B(n8055), .Z(n8070) );
  OR U8438 ( .A(n8017), .B(n8006), .Z(n8055) );
  XNOR U8439 ( .A(n8069), .B(n8052), .Z(n8006) );
  XNOR U8440 ( .A(n7994), .B(n8016), .Z(n8017) );
  ANDN U8441 ( .B(n8016), .A(n8007), .Z(n8071) );
  XOR U8442 ( .A(n8072), .B(n8073), .Z(n8026) );
  XOR U8443 ( .A(n8059), .B(n8049), .Z(n8073) );
  XOR U8444 ( .A(n8001), .B(n7721), .Z(n8049) );
  XOR U8445 ( .A(n8074), .B(n8061), .Z(n8059) );
  NANDN U8446 ( .A(n8011), .B(n8019), .Z(n8061) );
  XOR U8447 ( .A(n8027), .B(n7998), .Z(n8019) );
  XNOR U8448 ( .A(n8065), .B(n8075), .Z(n8016) );
  XNOR U8449 ( .A(n8076), .B(n8077), .Z(n8075) );
  XNOR U8450 ( .A(n8012), .B(n7837), .Z(n8011) );
  XNOR U8451 ( .A(n8007), .B(n8001), .Z(n7837) );
  IV U8452 ( .A(n8052), .Z(n8007) );
  XOR U8453 ( .A(n8078), .B(n8079), .Z(n8052) );
  XOR U8454 ( .A(n8080), .B(n8081), .Z(n8079) );
  XOR U8455 ( .A(n8069), .B(n8082), .Z(n8078) );
  AND U8456 ( .A(n8027), .B(n8012), .Z(n8074) );
  XOR U8457 ( .A(n7715), .B(n7831), .Z(n8012) );
  XOR U8458 ( .A(n8058), .B(n8083), .Z(n8072) );
  XNOR U8459 ( .A(n8084), .B(n8064), .Z(n8083) );
  OR U8460 ( .A(n7743), .B(n8002), .Z(n8064) );
  XNOR U8461 ( .A(n8085), .B(n8001), .Z(n8002) );
  XNOR U8462 ( .A(n7746), .B(n7721), .Z(n7743) );
  ANDN U8463 ( .B(n8001), .A(n7721), .Z(n8084) );
  XOR U8464 ( .A(n8086), .B(n8087), .Z(n7721) );
  XOR U8465 ( .A(n8076), .B(n8088), .Z(n8087) );
  XOR U8466 ( .A(n8089), .B(n8086), .Z(n8001) );
  XNOR U8467 ( .A(n7831), .B(n7746), .Z(n8058) );
  IV U8468 ( .A(n8085), .Z(n7831) );
  XNOR U8469 ( .A(n8077), .B(n8090), .Z(n8085) );
  XOR U8470 ( .A(n8082), .B(n8088), .Z(n8090) );
  IV U8471 ( .A(n8089), .Z(n8088) );
  XOR U8472 ( .A(n8091), .B(n8092), .Z(n8082) );
  XNOR U8473 ( .A(n8076), .B(n8093), .Z(n8092) );
  XNOR U8474 ( .A(n7471), .B(n6440), .Z(n8093) );
  XOR U8475 ( .A(n6459), .B(n7449), .Z(n6440) );
  XOR U8476 ( .A(n8094), .B(n8095), .Z(n7471) );
  XOR U8477 ( .A(n8096), .B(n8097), .Z(n8076) );
  XNOR U8478 ( .A(n7475), .B(n6403), .Z(n8097) );
  XNOR U8479 ( .A(key[913]), .B(n8098), .Z(n8096) );
  XNOR U8480 ( .A(n7478), .B(n8099), .Z(n8091) );
  XNOR U8481 ( .A(key[915]), .B(n7483), .Z(n8099) );
  XOR U8482 ( .A(n8100), .B(n8101), .Z(n8077) );
  XNOR U8483 ( .A(n7476), .B(n6442), .Z(n8101) );
  XOR U8484 ( .A(key[914]), .B(n7484), .Z(n8100) );
  XOR U8485 ( .A(n8065), .B(n7994), .Z(n8027) );
  XNOR U8486 ( .A(n8086), .B(n8102), .Z(n7994) );
  XOR U8487 ( .A(n8089), .B(n8081), .Z(n8102) );
  XNOR U8488 ( .A(n8103), .B(n8104), .Z(n8081) );
  XNOR U8489 ( .A(n7450), .B(n6434), .Z(n8104) );
  XNOR U8490 ( .A(n8105), .B(n7466), .Z(n6434) );
  XOR U8491 ( .A(n8106), .B(n8107), .Z(n7450) );
  XOR U8492 ( .A(n8108), .B(n8109), .Z(n8107) );
  XOR U8493 ( .A(n6437), .B(n8094), .Z(n8106) );
  XNOR U8494 ( .A(key[916]), .B(n8095), .Z(n8103) );
  IV U8495 ( .A(n7746), .Z(n8065) );
  XOR U8496 ( .A(n8086), .B(n8110), .Z(n7746) );
  XNOR U8497 ( .A(n8089), .B(n8080), .Z(n8110) );
  XOR U8498 ( .A(n8111), .B(n8112), .Z(n8080) );
  XOR U8499 ( .A(n8113), .B(n7460), .Z(n8112) );
  XOR U8500 ( .A(n6428), .B(n8114), .Z(n7460) );
  XOR U8501 ( .A(key[919]), .B(n8105), .Z(n8111) );
  XOR U8502 ( .A(n8115), .B(n8116), .Z(n8089) );
  XOR U8503 ( .A(n6413), .B(n7715), .Z(n8116) );
  IV U8504 ( .A(n8069), .Z(n7715) );
  XOR U8505 ( .A(n8117), .B(n8118), .Z(n8069) );
  XNOR U8506 ( .A(n6456), .B(n6446), .Z(n8118) );
  XNOR U8507 ( .A(n7494), .B(n8094), .Z(n6456) );
  XNOR U8508 ( .A(key[912]), .B(n8119), .Z(n8117) );
  XNOR U8509 ( .A(n8105), .B(n7461), .Z(n6413) );
  XNOR U8510 ( .A(n7464), .B(n8120), .Z(n8115) );
  XOR U8511 ( .A(key[918]), .B(n7489), .Z(n8120) );
  XOR U8512 ( .A(n8121), .B(n8113), .Z(n7489) );
  XNOR U8513 ( .A(n8094), .B(n8122), .Z(n8113) );
  XNOR U8514 ( .A(n8123), .B(n8124), .Z(n8086) );
  XOR U8515 ( .A(n7465), .B(n8125), .Z(n8124) );
  XNOR U8516 ( .A(n6419), .B(n8126), .Z(n7465) );
  XOR U8517 ( .A(key[917]), .B(n8109), .Z(n8123) );
  XOR U8518 ( .A(n2833), .B(n3787), .Z(n3809) );
  XOR U8519 ( .A(n7776), .B(n7627), .Z(n3787) );
  XNOR U8520 ( .A(n7667), .B(n8127), .Z(n7627) );
  XOR U8521 ( .A(n8128), .B(n7773), .Z(n8127) );
  XOR U8522 ( .A(n7755), .B(n7633), .Z(n7753) );
  ANDN U8523 ( .B(n7755), .A(n8130), .Z(n8128) );
  XNOR U8524 ( .A(n7771), .B(n8131), .Z(n7667) );
  XNOR U8525 ( .A(n8132), .B(n8133), .Z(n8131) );
  NAND U8526 ( .A(n7770), .B(n8134), .Z(n8133) );
  IV U8527 ( .A(n7688), .Z(n7776) );
  XNOR U8528 ( .A(n7771), .B(n8135), .Z(n7688) );
  XOR U8529 ( .A(n8136), .B(n7669), .Z(n8135) );
  OR U8530 ( .A(n8137), .B(n7781), .Z(n7669) );
  XNOR U8531 ( .A(n7671), .B(n7779), .Z(n7781) );
  NOR U8532 ( .A(n8138), .B(n7779), .Z(n8136) );
  XOR U8533 ( .A(n8139), .B(n8132), .Z(n7771) );
  OR U8534 ( .A(n7784), .B(n8140), .Z(n8132) );
  XNOR U8535 ( .A(n8141), .B(n7770), .Z(n7784) );
  XNOR U8536 ( .A(n7779), .B(n7633), .Z(n7770) );
  XOR U8537 ( .A(n8142), .B(n8143), .Z(n7633) );
  NANDN U8538 ( .A(n8144), .B(n8145), .Z(n8143) );
  XNOR U8539 ( .A(n8146), .B(n8147), .Z(n7779) );
  OR U8540 ( .A(n8144), .B(n8148), .Z(n8147) );
  ANDN U8541 ( .B(n8141), .A(n8149), .Z(n8139) );
  IV U8542 ( .A(n7787), .Z(n8141) );
  XOR U8543 ( .A(n7671), .B(n7755), .Z(n7787) );
  XNOR U8544 ( .A(n8150), .B(n8142), .Z(n7755) );
  NANDN U8545 ( .A(n8151), .B(n8152), .Z(n8142) );
  ANDN U8546 ( .B(n8153), .A(n8154), .Z(n8150) );
  NANDN U8547 ( .A(n8151), .B(n8156), .Z(n8146) );
  XOR U8548 ( .A(n8157), .B(n8144), .Z(n8151) );
  XNOR U8549 ( .A(n8158), .B(n8159), .Z(n8144) );
  XOR U8550 ( .A(n8160), .B(n8153), .Z(n8159) );
  XNOR U8551 ( .A(n8161), .B(n8162), .Z(n8158) );
  XNOR U8552 ( .A(n8163), .B(n8164), .Z(n8162) );
  ANDN U8553 ( .B(n8153), .A(n8165), .Z(n8163) );
  IV U8554 ( .A(n8166), .Z(n8153) );
  ANDN U8555 ( .B(n8157), .A(n8165), .Z(n8155) );
  IV U8556 ( .A(n8161), .Z(n8165) );
  IV U8557 ( .A(n8154), .Z(n8157) );
  XNOR U8558 ( .A(n8160), .B(n8167), .Z(n8154) );
  XOR U8559 ( .A(n8168), .B(n8164), .Z(n8167) );
  NAND U8560 ( .A(n8156), .B(n8152), .Z(n8164) );
  XNOR U8561 ( .A(n8145), .B(n8166), .Z(n8152) );
  XOR U8562 ( .A(n8169), .B(n8170), .Z(n8166) );
  XOR U8563 ( .A(n8171), .B(n8172), .Z(n8170) );
  XNOR U8564 ( .A(n7780), .B(n8173), .Z(n8172) );
  XNOR U8565 ( .A(n8174), .B(n8175), .Z(n8169) );
  XNOR U8566 ( .A(n8176), .B(n8177), .Z(n8175) );
  ANDN U8567 ( .B(n7765), .A(n7672), .Z(n8176) );
  XNOR U8568 ( .A(n8161), .B(n8148), .Z(n8156) );
  XOR U8569 ( .A(n8178), .B(n8179), .Z(n8161) );
  XNOR U8570 ( .A(n8180), .B(n8173), .Z(n8179) );
  XOR U8571 ( .A(n8181), .B(n8182), .Z(n8173) );
  XNOR U8572 ( .A(n8183), .B(n8184), .Z(n8182) );
  NAND U8573 ( .A(n8134), .B(n7769), .Z(n8184) );
  XNOR U8574 ( .A(n8185), .B(n8186), .Z(n8178) );
  ANDN U8575 ( .B(n8187), .A(n8130), .Z(n8185) );
  ANDN U8576 ( .B(n8145), .A(n8148), .Z(n8168) );
  XOR U8577 ( .A(n8148), .B(n8145), .Z(n8160) );
  XNOR U8578 ( .A(n8188), .B(n8189), .Z(n8145) );
  XNOR U8579 ( .A(n8181), .B(n8190), .Z(n8189) );
  XNOR U8580 ( .A(n8180), .B(n7765), .Z(n8190) );
  XNOR U8581 ( .A(n8191), .B(n8192), .Z(n8188) );
  XNOR U8582 ( .A(n8193), .B(n8177), .Z(n8192) );
  OR U8583 ( .A(n7782), .B(n8137), .Z(n8177) );
  XNOR U8584 ( .A(n8191), .B(n8174), .Z(n8137) );
  XNOR U8585 ( .A(n7765), .B(n7780), .Z(n7782) );
  ANDN U8586 ( .B(n7780), .A(n8138), .Z(n8193) );
  XOR U8587 ( .A(n8194), .B(n8195), .Z(n8148) );
  XOR U8588 ( .A(n8181), .B(n8171), .Z(n8195) );
  XOR U8589 ( .A(n7775), .B(n7634), .Z(n8171) );
  XOR U8590 ( .A(n8196), .B(n8183), .Z(n8181) );
  NANDN U8591 ( .A(n8140), .B(n7785), .Z(n8183) );
  XOR U8592 ( .A(n7786), .B(n7769), .Z(n7785) );
  XNOR U8593 ( .A(n8187), .B(n8197), .Z(n7780) );
  XNOR U8594 ( .A(n8198), .B(n8199), .Z(n8197) );
  XOR U8595 ( .A(n8149), .B(n8134), .Z(n8140) );
  XNOR U8596 ( .A(n8138), .B(n7775), .Z(n8134) );
  IV U8597 ( .A(n8174), .Z(n8138) );
  XOR U8598 ( .A(n8200), .B(n8201), .Z(n8174) );
  XOR U8599 ( .A(n8202), .B(n8203), .Z(n8201) );
  XOR U8600 ( .A(n8191), .B(n8204), .Z(n8200) );
  ANDN U8601 ( .B(n7786), .A(n8149), .Z(n8196) );
  XNOR U8602 ( .A(n8191), .B(n8205), .Z(n8149) );
  XOR U8603 ( .A(n8187), .B(n7765), .Z(n7786) );
  XNOR U8604 ( .A(n8206), .B(n8207), .Z(n7765) );
  XOR U8605 ( .A(n8208), .B(n8203), .Z(n8207) );
  XNOR U8606 ( .A(n8209), .B(n6131), .Z(n8203) );
  XOR U8607 ( .A(n8210), .B(n8211), .Z(n6131) );
  XOR U8608 ( .A(n7054), .B(n8212), .Z(n8211) );
  XOR U8609 ( .A(n8213), .B(n6120), .Z(n8210) );
  XOR U8610 ( .A(n7051), .B(n8214), .Z(n8209) );
  XNOR U8611 ( .A(key[1004]), .B(n8215), .Z(n8214) );
  XOR U8612 ( .A(n8216), .B(n8217), .Z(n7051) );
  IV U8613 ( .A(n7756), .Z(n8187) );
  XOR U8614 ( .A(n8180), .B(n8218), .Z(n8194) );
  XNOR U8615 ( .A(n8219), .B(n8186), .Z(n8218) );
  OR U8616 ( .A(n7754), .B(n8129), .Z(n8186) );
  XNOR U8617 ( .A(n8205), .B(n7775), .Z(n8129) );
  XNOR U8618 ( .A(n7756), .B(n7634), .Z(n7754) );
  ANDN U8619 ( .B(n7775), .A(n7634), .Z(n8219) );
  XOR U8620 ( .A(n8206), .B(n8220), .Z(n7634) );
  XOR U8621 ( .A(n8198), .B(n8221), .Z(n8220) );
  XOR U8622 ( .A(n8208), .B(n8206), .Z(n7775) );
  XNOR U8623 ( .A(n8130), .B(n7756), .Z(n8180) );
  XOR U8624 ( .A(n8206), .B(n8222), .Z(n7756) );
  XNOR U8625 ( .A(n8208), .B(n8202), .Z(n8222) );
  XOR U8626 ( .A(n8223), .B(n8224), .Z(n8202) );
  XNOR U8627 ( .A(n6151), .B(n6128), .Z(n8224) );
  XOR U8628 ( .A(n8225), .B(n8226), .Z(n6128) );
  XOR U8629 ( .A(key[1007]), .B(n8227), .Z(n8223) );
  XNOR U8630 ( .A(n8228), .B(n8229), .Z(n8206) );
  XOR U8631 ( .A(n8230), .B(n6121), .Z(n8229) );
  XOR U8632 ( .A(n7075), .B(n8217), .Z(n6121) );
  XNOR U8633 ( .A(n8231), .B(n8232), .Z(n8228) );
  XOR U8634 ( .A(key[1005]), .B(n8233), .Z(n8232) );
  IV U8635 ( .A(n8205), .Z(n8130) );
  XNOR U8636 ( .A(n8199), .B(n8234), .Z(n8205) );
  XOR U8637 ( .A(n8204), .B(n8221), .Z(n8234) );
  IV U8638 ( .A(n8208), .Z(n8221) );
  XOR U8639 ( .A(n8235), .B(n8236), .Z(n8208) );
  XNOR U8640 ( .A(n6114), .B(n7672), .Z(n8236) );
  IV U8641 ( .A(n8191), .Z(n7672) );
  XOR U8642 ( .A(n8237), .B(n8238), .Z(n8191) );
  XNOR U8643 ( .A(n6143), .B(n8216), .Z(n8238) );
  XNOR U8644 ( .A(n8239), .B(n8240), .Z(n8237) );
  XNOR U8645 ( .A(key[1000]), .B(n7069), .Z(n8240) );
  XNOR U8646 ( .A(n7074), .B(n6127), .Z(n6114) );
  XNOR U8647 ( .A(n8213), .B(n8241), .Z(n6127) );
  XNOR U8648 ( .A(n7065), .B(n8230), .Z(n7074) );
  XOR U8649 ( .A(n7064), .B(n8242), .Z(n8235) );
  XNOR U8650 ( .A(key[1006]), .B(n8243), .Z(n8242) );
  XOR U8651 ( .A(n8216), .B(n8226), .Z(n7064) );
  XOR U8652 ( .A(n8244), .B(n8245), .Z(n8204) );
  XNOR U8653 ( .A(n8198), .B(n8246), .Z(n8245) );
  XNOR U8654 ( .A(n7035), .B(n6137), .Z(n8246) );
  XNOR U8655 ( .A(n8213), .B(n6134), .Z(n6137) );
  XNOR U8656 ( .A(n7060), .B(n8212), .Z(n7035) );
  IV U8657 ( .A(n8216), .Z(n7060) );
  XOR U8658 ( .A(n8247), .B(n8248), .Z(n8198) );
  XNOR U8659 ( .A(n8249), .B(n8250), .Z(n8248) );
  XOR U8660 ( .A(n8251), .B(n8252), .Z(n8247) );
  XOR U8661 ( .A(key[1001]), .B(n6144), .Z(n8252) );
  XOR U8662 ( .A(n7039), .B(n8239), .Z(n6144) );
  XNOR U8663 ( .A(n8253), .B(n8254), .Z(n8244) );
  XNOR U8664 ( .A(key[1003]), .B(n6147), .Z(n8254) );
  XOR U8665 ( .A(n7042), .B(n8255), .Z(n6147) );
  XOR U8666 ( .A(n8256), .B(n8257), .Z(n8199) );
  XNOR U8667 ( .A(n6105), .B(n6145), .Z(n8257) );
  XNOR U8668 ( .A(n7045), .B(n8250), .Z(n6105) );
  XOR U8669 ( .A(n8255), .B(n8258), .Z(n8256) );
  XOR U8670 ( .A(key[1002]), .B(n8259), .Z(n8258) );
  XOR U8671 ( .A(n7649), .B(n7706), .Z(n2833) );
  XNOR U8672 ( .A(n7798), .B(n8260), .Z(n7706) );
  XOR U8673 ( .A(n8261), .B(n7678), .Z(n8260) );
  OR U8674 ( .A(n8262), .B(n7807), .Z(n7678) );
  XNOR U8675 ( .A(n7681), .B(n7806), .Z(n7807) );
  ANDN U8676 ( .B(n8263), .A(n8264), .Z(n8261) );
  XNOR U8677 ( .A(n7676), .B(n8265), .Z(n7649) );
  XNOR U8678 ( .A(n8266), .B(n7800), .Z(n8265) );
  XOR U8679 ( .A(n8268), .B(n7653), .Z(n7811) );
  ANDN U8680 ( .B(n8269), .A(n7814), .Z(n8266) );
  IV U8681 ( .A(n8268), .Z(n7814) );
  XNOR U8682 ( .A(n7798), .B(n8270), .Z(n7676) );
  XNOR U8683 ( .A(n8271), .B(n8272), .Z(n8270) );
  NANDN U8684 ( .A(n7818), .B(n8273), .Z(n8272) );
  XOR U8685 ( .A(n8274), .B(n8271), .Z(n7798) );
  OR U8686 ( .A(n7821), .B(n8275), .Z(n8271) );
  XNOR U8687 ( .A(n7824), .B(n7818), .Z(n7821) );
  XNOR U8688 ( .A(n7806), .B(n7653), .Z(n7818) );
  XOR U8689 ( .A(n8276), .B(n8277), .Z(n7653) );
  NANDN U8690 ( .A(n8278), .B(n8279), .Z(n8277) );
  IV U8691 ( .A(n8264), .Z(n7806) );
  XNOR U8692 ( .A(n8280), .B(n8281), .Z(n8264) );
  NANDN U8693 ( .A(n8278), .B(n8282), .Z(n8281) );
  NOR U8694 ( .A(n7824), .B(n8283), .Z(n8274) );
  XNOR U8695 ( .A(n8268), .B(n7681), .Z(n7824) );
  XNOR U8696 ( .A(n8284), .B(n8280), .Z(n7681) );
  NANDN U8697 ( .A(n8285), .B(n8286), .Z(n8280) );
  XOR U8698 ( .A(n8282), .B(n8287), .Z(n8286) );
  ANDN U8699 ( .B(n8287), .A(n8288), .Z(n8284) );
  XNOR U8700 ( .A(n8289), .B(n8276), .Z(n8268) );
  NANDN U8701 ( .A(n8285), .B(n8290), .Z(n8276) );
  XOR U8702 ( .A(n8291), .B(n8279), .Z(n8290) );
  XNOR U8703 ( .A(n8292), .B(n8293), .Z(n8278) );
  XOR U8704 ( .A(n8294), .B(n8295), .Z(n8293) );
  XNOR U8705 ( .A(n8296), .B(n8297), .Z(n8292) );
  XNOR U8706 ( .A(n8298), .B(n8299), .Z(n8297) );
  ANDN U8707 ( .B(n8291), .A(n8295), .Z(n8298) );
  ANDN U8708 ( .B(n8291), .A(n8288), .Z(n8289) );
  XNOR U8709 ( .A(n8294), .B(n8300), .Z(n8288) );
  XOR U8710 ( .A(n8301), .B(n8299), .Z(n8300) );
  NAND U8711 ( .A(n8302), .B(n8303), .Z(n8299) );
  XNOR U8712 ( .A(n8296), .B(n8279), .Z(n8303) );
  IV U8713 ( .A(n8291), .Z(n8296) );
  XNOR U8714 ( .A(n8282), .B(n8295), .Z(n8302) );
  IV U8715 ( .A(n8287), .Z(n8295) );
  XOR U8716 ( .A(n8304), .B(n8305), .Z(n8287) );
  XNOR U8717 ( .A(n8306), .B(n8307), .Z(n8305) );
  XNOR U8718 ( .A(n8308), .B(n8309), .Z(n8304) );
  ANDN U8719 ( .B(n8269), .A(n8310), .Z(n8308) );
  AND U8720 ( .A(n8279), .B(n8282), .Z(n8301) );
  XNOR U8721 ( .A(n8279), .B(n8282), .Z(n8294) );
  XNOR U8722 ( .A(n8311), .B(n8312), .Z(n8282) );
  XNOR U8723 ( .A(n8313), .B(n8307), .Z(n8312) );
  XOR U8724 ( .A(n8314), .B(n8315), .Z(n8311) );
  XNOR U8725 ( .A(n8316), .B(n8309), .Z(n8315) );
  OR U8726 ( .A(n7812), .B(n8267), .Z(n8309) );
  XNOR U8727 ( .A(n8269), .B(n8317), .Z(n8267) );
  XNOR U8728 ( .A(n8310), .B(n7654), .Z(n7812) );
  ANDN U8729 ( .B(n8318), .A(n7802), .Z(n8316) );
  XNOR U8730 ( .A(n8319), .B(n8320), .Z(n8279) );
  XNOR U8731 ( .A(n8307), .B(n8321), .Z(n8320) );
  XOR U8732 ( .A(n7797), .B(n8314), .Z(n8321) );
  XNOR U8733 ( .A(n8269), .B(n8310), .Z(n8307) );
  XNOR U8734 ( .A(n8322), .B(n8323), .Z(n8319) );
  XNOR U8735 ( .A(n8324), .B(n8325), .Z(n8323) );
  ANDN U8736 ( .B(n8263), .A(n7805), .Z(n8324) );
  XNOR U8737 ( .A(n8326), .B(n8327), .Z(n8291) );
  XNOR U8738 ( .A(n8313), .B(n8328), .Z(n8327) );
  XNOR U8739 ( .A(n7805), .B(n8306), .Z(n8328) );
  XOR U8740 ( .A(n8314), .B(n8329), .Z(n8306) );
  XNOR U8741 ( .A(n8330), .B(n8331), .Z(n8329) );
  NAND U8742 ( .A(n8273), .B(n7819), .Z(n8331) );
  XNOR U8743 ( .A(n8332), .B(n8330), .Z(n8314) );
  NANDN U8744 ( .A(n8275), .B(n7822), .Z(n8330) );
  XOR U8745 ( .A(n7823), .B(n7819), .Z(n7822) );
  XNOR U8746 ( .A(n8333), .B(n7654), .Z(n7819) );
  XOR U8747 ( .A(n8283), .B(n8273), .Z(n8275) );
  XOR U8748 ( .A(n8263), .B(n8317), .Z(n8273) );
  ANDN U8749 ( .B(n7823), .A(n8283), .Z(n8332) );
  XNOR U8750 ( .A(n8322), .B(n8269), .Z(n8283) );
  XNOR U8751 ( .A(n8334), .B(n8335), .Z(n8269) );
  XNOR U8752 ( .A(n8336), .B(n8337), .Z(n8335) );
  XOR U8753 ( .A(n8338), .B(n7813), .Z(n7823) );
  XOR U8754 ( .A(n8317), .B(n8318), .Z(n8313) );
  IV U8755 ( .A(n7654), .Z(n8318) );
  XOR U8756 ( .A(n8339), .B(n8340), .Z(n7654) );
  XNOR U8757 ( .A(n8341), .B(n8337), .Z(n8340) );
  IV U8758 ( .A(n7802), .Z(n8317) );
  XOR U8759 ( .A(n8337), .B(n8342), .Z(n7802) );
  XNOR U8760 ( .A(n8263), .B(n8343), .Z(n8326) );
  XNOR U8761 ( .A(n8344), .B(n8325), .Z(n8343) );
  OR U8762 ( .A(n7808), .B(n8262), .Z(n8325) );
  XNOR U8763 ( .A(n8322), .B(n8263), .Z(n8262) );
  XOR U8764 ( .A(n7797), .B(n8333), .Z(n7808) );
  IV U8765 ( .A(n7805), .Z(n8333) );
  XOR U8766 ( .A(n7813), .B(n8345), .Z(n7805) );
  XNOR U8767 ( .A(n8341), .B(n8334), .Z(n8345) );
  XOR U8768 ( .A(n8346), .B(n8347), .Z(n8334) );
  XNOR U8769 ( .A(n7226), .B(n8348), .Z(n8347) );
  XNOR U8770 ( .A(key[962]), .B(n7220), .Z(n8346) );
  IV U8771 ( .A(n8310), .Z(n7813) );
  XOR U8772 ( .A(n8339), .B(n8349), .Z(n8310) );
  XOR U8773 ( .A(n8337), .B(n8350), .Z(n8349) );
  ANDN U8774 ( .B(n8338), .A(n7680), .Z(n8344) );
  IV U8775 ( .A(n7797), .Z(n8338) );
  XOR U8776 ( .A(n8339), .B(n8351), .Z(n7797) );
  XOR U8777 ( .A(n8337), .B(n8352), .Z(n8351) );
  XOR U8778 ( .A(n8353), .B(n8354), .Z(n8337) );
  XOR U8779 ( .A(n6273), .B(n7680), .Z(n8354) );
  IV U8780 ( .A(n8322), .Z(n7680) );
  XNOR U8781 ( .A(n8355), .B(n7198), .Z(n6273) );
  XNOR U8782 ( .A(n7201), .B(n8356), .Z(n8353) );
  XOR U8783 ( .A(key[966]), .B(n7208), .Z(n8356) );
  XOR U8784 ( .A(n8357), .B(n8358), .Z(n7208) );
  IV U8785 ( .A(n8342), .Z(n8339) );
  XOR U8786 ( .A(n8359), .B(n8360), .Z(n8342) );
  XOR U8787 ( .A(n7202), .B(n8361), .Z(n8360) );
  XNOR U8788 ( .A(n6279), .B(n8362), .Z(n7202) );
  XOR U8789 ( .A(key[965]), .B(n8363), .Z(n8359) );
  XOR U8790 ( .A(n8364), .B(n8365), .Z(n8263) );
  XNOR U8791 ( .A(n8352), .B(n8350), .Z(n8365) );
  XNOR U8792 ( .A(n8366), .B(n8367), .Z(n8350) );
  XOR U8793 ( .A(n8358), .B(n7197), .Z(n8367) );
  XOR U8794 ( .A(n6288), .B(n8368), .Z(n7197) );
  XOR U8795 ( .A(n8369), .B(n8370), .Z(n8358) );
  XOR U8796 ( .A(key[967]), .B(n8355), .Z(n8366) );
  XNOR U8797 ( .A(n8371), .B(n8372), .Z(n8352) );
  XOR U8798 ( .A(n7185), .B(n6294), .Z(n8372) );
  XNOR U8799 ( .A(n8355), .B(n7203), .Z(n6294) );
  XOR U8800 ( .A(n6297), .B(n8373), .Z(n7185) );
  XNOR U8801 ( .A(n7184), .B(n8374), .Z(n8371) );
  XNOR U8802 ( .A(key[964]), .B(n8375), .Z(n8374) );
  XOR U8803 ( .A(n8369), .B(n8363), .Z(n7184) );
  XOR U8804 ( .A(n8322), .B(n8336), .Z(n8364) );
  XOR U8805 ( .A(n8376), .B(n8377), .Z(n8336) );
  XNOR U8806 ( .A(n8341), .B(n8378), .Z(n8377) );
  XNOR U8807 ( .A(n7225), .B(n6300), .Z(n8378) );
  XNOR U8808 ( .A(n6319), .B(n7186), .Z(n6300) );
  IV U8809 ( .A(n8355), .Z(n6319) );
  XOR U8810 ( .A(n8379), .B(n8380), .Z(n8341) );
  XOR U8811 ( .A(n7218), .B(n6263), .Z(n8380) );
  XNOR U8812 ( .A(key[961]), .B(n8381), .Z(n8379) );
  XNOR U8813 ( .A(n7213), .B(n8382), .Z(n8376) );
  XNOR U8814 ( .A(key[963]), .B(n7221), .Z(n8382) );
  XNOR U8815 ( .A(n8369), .B(n8375), .Z(n7213) );
  XOR U8816 ( .A(n8383), .B(n8384), .Z(n8322) );
  XNOR U8817 ( .A(n6316), .B(n6306), .Z(n8384) );
  XOR U8818 ( .A(n7231), .B(n8369), .Z(n6316) );
  XNOR U8819 ( .A(key[960]), .B(n8385), .Z(n8383) );
  XNOR U8820 ( .A(key[1184]), .B(n4437), .Z(n5683) );
  XOR U8821 ( .A(n5599), .B(n5494), .Z(n4437) );
  XNOR U8822 ( .A(n5527), .B(n8386), .Z(n5494) );
  XOR U8823 ( .A(n8387), .B(n5680), .Z(n8386) );
  XOR U8824 ( .A(n5656), .B(n5500), .Z(n5654) );
  ANDN U8825 ( .B(n5656), .A(n8389), .Z(n8387) );
  XNOR U8826 ( .A(n5678), .B(n8390), .Z(n5527) );
  XNOR U8827 ( .A(n8391), .B(n8392), .Z(n8390) );
  NAND U8828 ( .A(n5672), .B(n8393), .Z(n8392) );
  IV U8829 ( .A(n5545), .Z(n5599) );
  XNOR U8830 ( .A(n5678), .B(n8394), .Z(n5545) );
  XOR U8831 ( .A(n8395), .B(n5529), .Z(n8394) );
  OR U8832 ( .A(n8396), .B(n5666), .Z(n5529) );
  XNOR U8833 ( .A(n5531), .B(n5661), .Z(n5666) );
  NOR U8834 ( .A(n8397), .B(n5661), .Z(n8395) );
  XOR U8835 ( .A(n8398), .B(n8391), .Z(n5678) );
  OR U8836 ( .A(n5674), .B(n8399), .Z(n8391) );
  XNOR U8837 ( .A(n8400), .B(n5672), .Z(n5674) );
  XNOR U8838 ( .A(n5661), .B(n5500), .Z(n5672) );
  XOR U8839 ( .A(n8401), .B(n8402), .Z(n5500) );
  NANDN U8840 ( .A(n8403), .B(n8404), .Z(n8402) );
  XNOR U8841 ( .A(n8405), .B(n8406), .Z(n5661) );
  OR U8842 ( .A(n8403), .B(n8407), .Z(n8406) );
  ANDN U8843 ( .B(n8400), .A(n8408), .Z(n8398) );
  IV U8844 ( .A(n5677), .Z(n8400) );
  XOR U8845 ( .A(n5531), .B(n5656), .Z(n5677) );
  XNOR U8846 ( .A(n8409), .B(n8401), .Z(n5656) );
  NANDN U8847 ( .A(n8410), .B(n8411), .Z(n8401) );
  ANDN U8848 ( .B(n8412), .A(n8413), .Z(n8409) );
  NANDN U8849 ( .A(n8410), .B(n8415), .Z(n8405) );
  XOR U8850 ( .A(n8416), .B(n8403), .Z(n8410) );
  XNOR U8851 ( .A(n8417), .B(n8418), .Z(n8403) );
  XOR U8852 ( .A(n8419), .B(n8412), .Z(n8418) );
  XNOR U8853 ( .A(n8420), .B(n8421), .Z(n8417) );
  XNOR U8854 ( .A(n8422), .B(n8423), .Z(n8421) );
  ANDN U8855 ( .B(n8412), .A(n8424), .Z(n8422) );
  IV U8856 ( .A(n8425), .Z(n8412) );
  ANDN U8857 ( .B(n8416), .A(n8424), .Z(n8414) );
  IV U8858 ( .A(n8420), .Z(n8424) );
  IV U8859 ( .A(n8413), .Z(n8416) );
  XNOR U8860 ( .A(n8419), .B(n8426), .Z(n8413) );
  XOR U8861 ( .A(n8427), .B(n8423), .Z(n8426) );
  NAND U8862 ( .A(n8415), .B(n8411), .Z(n8423) );
  XNOR U8863 ( .A(n8404), .B(n8425), .Z(n8411) );
  XOR U8864 ( .A(n8428), .B(n8429), .Z(n8425) );
  XOR U8865 ( .A(n8430), .B(n8431), .Z(n8429) );
  XNOR U8866 ( .A(n5662), .B(n8432), .Z(n8431) );
  XNOR U8867 ( .A(n8433), .B(n8434), .Z(n8428) );
  XNOR U8868 ( .A(n8435), .B(n8436), .Z(n8434) );
  ANDN U8869 ( .B(n5665), .A(n5532), .Z(n8435) );
  XNOR U8870 ( .A(n8420), .B(n8407), .Z(n8415) );
  XOR U8871 ( .A(n8437), .B(n8438), .Z(n8420) );
  XNOR U8872 ( .A(n8439), .B(n8432), .Z(n8438) );
  XOR U8873 ( .A(n8440), .B(n8441), .Z(n8432) );
  XNOR U8874 ( .A(n8442), .B(n8443), .Z(n8441) );
  NAND U8875 ( .A(n8393), .B(n5671), .Z(n8443) );
  XNOR U8876 ( .A(n8444), .B(n8445), .Z(n8437) );
  ANDN U8877 ( .B(n8446), .A(n8389), .Z(n8444) );
  ANDN U8878 ( .B(n8404), .A(n8407), .Z(n8427) );
  XOR U8879 ( .A(n8407), .B(n8404), .Z(n8419) );
  XNOR U8880 ( .A(n8447), .B(n8448), .Z(n8404) );
  XNOR U8881 ( .A(n8440), .B(n8449), .Z(n8448) );
  XNOR U8882 ( .A(n8439), .B(n5665), .Z(n8449) );
  XNOR U8883 ( .A(n8450), .B(n8451), .Z(n8447) );
  XNOR U8884 ( .A(n8452), .B(n8436), .Z(n8451) );
  OR U8885 ( .A(n5667), .B(n8396), .Z(n8436) );
  XNOR U8886 ( .A(n8450), .B(n8433), .Z(n8396) );
  XNOR U8887 ( .A(n5665), .B(n5662), .Z(n5667) );
  ANDN U8888 ( .B(n5662), .A(n8397), .Z(n8452) );
  XOR U8889 ( .A(n8453), .B(n8454), .Z(n8407) );
  XOR U8890 ( .A(n8440), .B(n8430), .Z(n8454) );
  XOR U8891 ( .A(n5682), .B(n5501), .Z(n8430) );
  XOR U8892 ( .A(n8455), .B(n8442), .Z(n8440) );
  NANDN U8893 ( .A(n8399), .B(n5675), .Z(n8442) );
  XOR U8894 ( .A(n5676), .B(n5671), .Z(n5675) );
  XNOR U8895 ( .A(n8446), .B(n8456), .Z(n5662) );
  XNOR U8896 ( .A(n8457), .B(n8458), .Z(n8456) );
  XOR U8897 ( .A(n8408), .B(n8393), .Z(n8399) );
  XNOR U8898 ( .A(n8397), .B(n5682), .Z(n8393) );
  IV U8899 ( .A(n8433), .Z(n8397) );
  XOR U8900 ( .A(n8459), .B(n8460), .Z(n8433) );
  XOR U8901 ( .A(n8461), .B(n8462), .Z(n8460) );
  XOR U8902 ( .A(n8450), .B(n8463), .Z(n8459) );
  ANDN U8903 ( .B(n5676), .A(n8408), .Z(n8455) );
  XNOR U8904 ( .A(n8450), .B(n8464), .Z(n8408) );
  XOR U8905 ( .A(n8446), .B(n5665), .Z(n5676) );
  XNOR U8906 ( .A(n8465), .B(n8466), .Z(n5665) );
  XOR U8907 ( .A(n8467), .B(n8462), .Z(n8466) );
  XNOR U8908 ( .A(n8468), .B(n8469), .Z(n8462) );
  XOR U8909 ( .A(n4923), .B(n4922), .Z(n8469) );
  XNOR U8910 ( .A(n4235), .B(n2974), .Z(n4922) );
  XOR U8911 ( .A(n8470), .B(n3012), .Z(n4235) );
  XOR U8912 ( .A(n4275), .B(n4254), .Z(n4923) );
  IV U8913 ( .A(n4938), .Z(n4254) );
  XOR U8914 ( .A(n8471), .B(n8472), .Z(n4938) );
  XNOR U8915 ( .A(n8473), .B(n8474), .Z(n8472) );
  XNOR U8916 ( .A(n8475), .B(n8476), .Z(n8471) );
  XOR U8917 ( .A(n8477), .B(n8478), .Z(n8476) );
  ANDN U8918 ( .B(n8479), .A(n8480), .Z(n8478) );
  XOR U8919 ( .A(n4233), .B(n8481), .Z(n8468) );
  XNOR U8920 ( .A(key[1132]), .B(n4231), .Z(n8481) );
  XNOR U8921 ( .A(n4249), .B(n2979), .Z(n4231) );
  XNOR U8922 ( .A(n8482), .B(n3010), .Z(n4233) );
  IV U8923 ( .A(n5657), .Z(n8446) );
  XOR U8924 ( .A(n8439), .B(n8483), .Z(n8453) );
  XNOR U8925 ( .A(n8484), .B(n8445), .Z(n8483) );
  OR U8926 ( .A(n5655), .B(n8388), .Z(n8445) );
  XNOR U8927 ( .A(n8464), .B(n5682), .Z(n8388) );
  XNOR U8928 ( .A(n5657), .B(n5501), .Z(n5655) );
  ANDN U8929 ( .B(n5682), .A(n5501), .Z(n8484) );
  XOR U8930 ( .A(n8465), .B(n8485), .Z(n5501) );
  XOR U8931 ( .A(n8457), .B(n8486), .Z(n8485) );
  XOR U8932 ( .A(n8467), .B(n8465), .Z(n5682) );
  XNOR U8933 ( .A(n8389), .B(n5657), .Z(n8439) );
  XOR U8934 ( .A(n8465), .B(n8487), .Z(n5657) );
  XNOR U8935 ( .A(n8467), .B(n8461), .Z(n8487) );
  XOR U8936 ( .A(n8488), .B(n8489), .Z(n8461) );
  XOR U8937 ( .A(n4948), .B(n4934), .Z(n8489) );
  XNOR U8938 ( .A(n2986), .B(n4270), .Z(n4934) );
  XNOR U8939 ( .A(n8490), .B(n8491), .Z(n4270) );
  XNOR U8940 ( .A(n8492), .B(n8493), .Z(n8491) );
  XNOR U8941 ( .A(n8494), .B(n8495), .Z(n8490) );
  XOR U8942 ( .A(n4275), .B(n4249), .Z(n4948) );
  XOR U8943 ( .A(key[1135]), .B(n4248), .Z(n8488) );
  XNOR U8944 ( .A(n8496), .B(n8497), .Z(n4248) );
  XNOR U8945 ( .A(n8498), .B(n8499), .Z(n8497) );
  XNOR U8946 ( .A(n8500), .B(n8501), .Z(n8496) );
  XNOR U8947 ( .A(n8502), .B(n8503), .Z(n8465) );
  XOR U8948 ( .A(n8504), .B(n4939), .Z(n8503) );
  XOR U8949 ( .A(n4237), .B(n2979), .Z(n4939) );
  XNOR U8950 ( .A(n8505), .B(n8506), .Z(n2979) );
  XNOR U8951 ( .A(n8507), .B(n8508), .Z(n8506) );
  XNOR U8952 ( .A(n8509), .B(n8510), .Z(n8505) );
  XOR U8953 ( .A(n8511), .B(n8512), .Z(n8510) );
  ANDN U8954 ( .B(n8513), .A(n8514), .Z(n8512) );
  XNOR U8955 ( .A(n8515), .B(n8516), .Z(n4237) );
  XNOR U8956 ( .A(n8470), .B(n8493), .Z(n8516) );
  XNOR U8957 ( .A(n8517), .B(n8518), .Z(n8493) );
  XNOR U8958 ( .A(n8519), .B(n8520), .Z(n8518) );
  NANDN U8959 ( .A(n8521), .B(n8522), .Z(n8520) );
  XNOR U8960 ( .A(n8523), .B(n8524), .Z(n8515) );
  XOR U8961 ( .A(n8525), .B(n8526), .Z(n8524) );
  ANDN U8962 ( .B(n8527), .A(n8528), .Z(n8526) );
  XOR U8963 ( .A(n4253), .B(n8529), .Z(n8502) );
  XNOR U8964 ( .A(key[1133]), .B(n4940), .Z(n8529) );
  XOR U8965 ( .A(n8530), .B(n8531), .Z(n4940) );
  XNOR U8966 ( .A(n8532), .B(n8533), .Z(n4253) );
  XNOR U8967 ( .A(n8534), .B(n8499), .Z(n8533) );
  XNOR U8968 ( .A(n8535), .B(n8536), .Z(n8499) );
  XNOR U8969 ( .A(n8537), .B(n8538), .Z(n8536) );
  NANDN U8970 ( .A(n8539), .B(n8540), .Z(n8538) );
  XNOR U8971 ( .A(n8482), .B(n8541), .Z(n8532) );
  XOR U8972 ( .A(n8542), .B(n8543), .Z(n8541) );
  ANDN U8973 ( .B(n8544), .A(n8545), .Z(n8543) );
  IV U8974 ( .A(n8464), .Z(n8389) );
  XNOR U8975 ( .A(n8458), .B(n8546), .Z(n8464) );
  XOR U8976 ( .A(n8463), .B(n8486), .Z(n8546) );
  IV U8977 ( .A(n8467), .Z(n8486) );
  XOR U8978 ( .A(n8547), .B(n8548), .Z(n8467) );
  XNOR U8979 ( .A(n4944), .B(n5532), .Z(n8548) );
  IV U8980 ( .A(n8450), .Z(n5532) );
  XOR U8981 ( .A(n8549), .B(n8550), .Z(n8450) );
  XOR U8982 ( .A(n4249), .B(n4949), .Z(n8550) );
  XNOR U8983 ( .A(n8530), .B(n8551), .Z(n4949) );
  XNOR U8984 ( .A(n8552), .B(n8553), .Z(n8551) );
  XNOR U8985 ( .A(n4276), .B(n8554), .Z(n8549) );
  XNOR U8986 ( .A(key[1128]), .B(n8555), .Z(n8554) );
  XNOR U8987 ( .A(n4950), .B(n3022), .Z(n4276) );
  IV U8988 ( .A(n4935), .Z(n3022) );
  XOR U8989 ( .A(n8556), .B(n8482), .Z(n4935) );
  XNOR U8990 ( .A(n8535), .B(n8557), .Z(n8482) );
  XNOR U8991 ( .A(n8558), .B(n8559), .Z(n8557) );
  ANDN U8992 ( .B(n8560), .A(n8561), .Z(n8558) );
  XNOR U8993 ( .A(n8562), .B(n8563), .Z(n8535) );
  XNOR U8994 ( .A(n8564), .B(n8565), .Z(n8563) );
  NANDN U8995 ( .A(n8566), .B(n8567), .Z(n8565) );
  IV U8996 ( .A(n4236), .Z(n4950) );
  XNOR U8997 ( .A(n8517), .B(n8568), .Z(n8470) );
  XOR U8998 ( .A(n8569), .B(n8570), .Z(n8568) );
  ANDN U8999 ( .B(n8571), .A(n8572), .Z(n8569) );
  XNOR U9000 ( .A(n8573), .B(n8574), .Z(n8517) );
  XNOR U9001 ( .A(n8575), .B(n8576), .Z(n8574) );
  NAND U9002 ( .A(n8577), .B(n8578), .Z(n8576) );
  XOR U9003 ( .A(n4252), .B(n4933), .Z(n4944) );
  XOR U9004 ( .A(n4275), .B(n4247), .Z(n4933) );
  XNOR U9005 ( .A(n8580), .B(n8581), .Z(n4247) );
  XNOR U9006 ( .A(n8530), .B(n8474), .Z(n8581) );
  XNOR U9007 ( .A(n8582), .B(n8583), .Z(n8474) );
  XNOR U9008 ( .A(n8584), .B(n8585), .Z(n8583) );
  NANDN U9009 ( .A(n8586), .B(n8587), .Z(n8585) );
  XOR U9010 ( .A(n8588), .B(n8589), .Z(n8530) );
  XOR U9011 ( .A(n8552), .B(n8553), .Z(n8580) );
  XOR U9012 ( .A(n2981), .B(n8504), .Z(n4252) );
  IV U9013 ( .A(n3000), .Z(n8504) );
  XOR U9014 ( .A(n8590), .B(n8591), .Z(n3000) );
  XOR U9015 ( .A(n8494), .B(n8592), .Z(n2981) );
  XNOR U9016 ( .A(n2983), .B(n8593), .Z(n8547) );
  XNOR U9017 ( .A(key[1134]), .B(n4271), .Z(n8593) );
  XOR U9018 ( .A(n4249), .B(n2986), .Z(n4271) );
  XOR U9019 ( .A(n8594), .B(n8595), .Z(n2986) );
  XNOR U9020 ( .A(n8590), .B(n8508), .Z(n8595) );
  XNOR U9021 ( .A(n8596), .B(n8597), .Z(n8508) );
  XNOR U9022 ( .A(n8598), .B(n8599), .Z(n8597) );
  NANDN U9023 ( .A(n8600), .B(n8601), .Z(n8599) );
  IV U9024 ( .A(n8602), .Z(n8590) );
  XNOR U9025 ( .A(n8603), .B(n8604), .Z(n8594) );
  XOR U9026 ( .A(n8501), .B(n8605), .Z(n2983) );
  XOR U9027 ( .A(n8606), .B(n8607), .Z(n8463) );
  XNOR U9028 ( .A(n8457), .B(n8608), .Z(n8607) );
  XNOR U9029 ( .A(n2993), .B(n4954), .Z(n8608) );
  XNOR U9030 ( .A(n4275), .B(n4232), .Z(n4954) );
  XNOR U9031 ( .A(n8475), .B(n4957), .Z(n4232) );
  XOR U9032 ( .A(n8588), .B(n8475), .Z(n4275) );
  XNOR U9033 ( .A(n8582), .B(n8609), .Z(n8475) );
  XNOR U9034 ( .A(n8610), .B(n8611), .Z(n8609) );
  ANDN U9035 ( .B(n8612), .A(n8613), .Z(n8610) );
  XNOR U9036 ( .A(n8614), .B(n8615), .Z(n8582) );
  XNOR U9037 ( .A(n8616), .B(n8617), .Z(n8615) );
  NANDN U9038 ( .A(n8618), .B(n8619), .Z(n8617) );
  IV U9039 ( .A(n8620), .Z(n8588) );
  XNOR U9040 ( .A(n8621), .B(n8622), .Z(n2993) );
  XOR U9041 ( .A(n8498), .B(n8605), .Z(n8622) );
  XOR U9042 ( .A(n8623), .B(n8624), .Z(n8605) );
  XNOR U9043 ( .A(n8625), .B(n8542), .Z(n8624) );
  ANDN U9044 ( .B(n8626), .A(n8627), .Z(n8542) );
  ANDN U9045 ( .B(n8628), .A(n8561), .Z(n8625) );
  IV U9046 ( .A(n8629), .Z(n8561) );
  XOR U9047 ( .A(n8630), .B(n8631), .Z(n8621) );
  XOR U9048 ( .A(n8632), .B(n8633), .Z(n8457) );
  XNOR U9049 ( .A(n2992), .B(n3020), .Z(n8633) );
  XOR U9050 ( .A(n8498), .B(n8634), .Z(n3020) );
  XNOR U9051 ( .A(n8630), .B(n8501), .Z(n8634) );
  XOR U9052 ( .A(n8556), .B(n8631), .Z(n8501) );
  XNOR U9053 ( .A(n8534), .B(n8635), .Z(n8631) );
  XNOR U9054 ( .A(n8636), .B(n8637), .Z(n8635) );
  NANDN U9055 ( .A(n8638), .B(n8639), .Z(n8637) );
  IV U9056 ( .A(n8640), .Z(n8556) );
  XNOR U9057 ( .A(n8623), .B(n8641), .Z(n8498) );
  XNOR U9058 ( .A(n8636), .B(n8642), .Z(n8641) );
  NANDN U9059 ( .A(n8643), .B(n8540), .Z(n8642) );
  OR U9060 ( .A(n8644), .B(n8645), .Z(n8636) );
  XNOR U9061 ( .A(n8534), .B(n8646), .Z(n8623) );
  XNOR U9062 ( .A(n8647), .B(n8648), .Z(n8646) );
  NANDN U9063 ( .A(n8566), .B(n8649), .Z(n8648) );
  XOR U9064 ( .A(n8650), .B(n8647), .Z(n8534) );
  NANDN U9065 ( .A(n8651), .B(n8652), .Z(n8647) );
  ANDN U9066 ( .B(n8653), .A(n8654), .Z(n8650) );
  XOR U9067 ( .A(n4957), .B(n8655), .Z(n8632) );
  XNOR U9068 ( .A(key[1129]), .B(n4277), .Z(n8655) );
  XNOR U9069 ( .A(n3014), .B(n3024), .Z(n4277) );
  XNOR U9070 ( .A(n8656), .B(n8657), .Z(n3024) );
  XOR U9071 ( .A(n8579), .B(n8658), .Z(n8494) );
  IV U9072 ( .A(n8555), .Z(n3014) );
  XOR U9073 ( .A(n8602), .B(n8659), .Z(n8555) );
  XOR U9074 ( .A(n8603), .B(n8604), .Z(n8659) );
  IV U9075 ( .A(n8660), .Z(n8603) );
  XOR U9076 ( .A(n8661), .B(n8662), .Z(n8602) );
  XNOR U9077 ( .A(n8620), .B(n8552), .Z(n4957) );
  XNOR U9078 ( .A(n8614), .B(n8663), .Z(n8620) );
  XOR U9079 ( .A(n8664), .B(n8584), .Z(n8663) );
  OR U9080 ( .A(n8665), .B(n8666), .Z(n8584) );
  ANDN U9081 ( .B(n8667), .A(n8668), .Z(n8664) );
  XNOR U9082 ( .A(n4259), .B(n8669), .Z(n8606) );
  XOR U9083 ( .A(key[1131]), .B(n4960), .Z(n8669) );
  XOR U9084 ( .A(n2996), .B(n3017), .Z(n4960) );
  XOR U9085 ( .A(n8670), .B(n8671), .Z(n2996) );
  XNOR U9086 ( .A(n8656), .B(n8592), .Z(n8671) );
  XNOR U9087 ( .A(n8672), .B(n8673), .Z(n8592) );
  XNOR U9088 ( .A(n8674), .B(n8525), .Z(n8673) );
  ANDN U9089 ( .B(n8675), .A(n8676), .Z(n8525) );
  NOR U9090 ( .A(n8677), .B(n8572), .Z(n8674) );
  IV U9091 ( .A(n8492), .Z(n8656) );
  XOR U9092 ( .A(n8672), .B(n8678), .Z(n8492) );
  XNOR U9093 ( .A(n8679), .B(n8680), .Z(n8678) );
  NANDN U9094 ( .A(n8681), .B(n8522), .Z(n8680) );
  XOR U9095 ( .A(n8523), .B(n8682), .Z(n8672) );
  XNOR U9096 ( .A(n8683), .B(n8684), .Z(n8682) );
  NAND U9097 ( .A(n8685), .B(n8577), .Z(n8684) );
  XOR U9098 ( .A(n8658), .B(n8495), .Z(n8670) );
  XNOR U9099 ( .A(n8523), .B(n8686), .Z(n8658) );
  XNOR U9100 ( .A(n8679), .B(n8687), .Z(n8686) );
  NANDN U9101 ( .A(n8688), .B(n8689), .Z(n8687) );
  OR U9102 ( .A(n8690), .B(n8691), .Z(n8679) );
  XOR U9103 ( .A(n8692), .B(n8683), .Z(n8523) );
  NANDN U9104 ( .A(n8693), .B(n8694), .Z(n8683) );
  ANDN U9105 ( .B(n8695), .A(n8696), .Z(n8692) );
  XOR U9106 ( .A(n4249), .B(n2974), .Z(n4259) );
  XOR U9107 ( .A(n8507), .B(n2992), .Z(n2974) );
  XOR U9108 ( .A(n8661), .B(n8507), .Z(n4249) );
  XNOR U9109 ( .A(n8596), .B(n8697), .Z(n8507) );
  XNOR U9110 ( .A(n8698), .B(n8699), .Z(n8697) );
  ANDN U9111 ( .B(n8700), .A(n8701), .Z(n8698) );
  XNOR U9112 ( .A(n8702), .B(n8703), .Z(n8596) );
  XNOR U9113 ( .A(n8704), .B(n8705), .Z(n8703) );
  NANDN U9114 ( .A(n8706), .B(n8707), .Z(n8705) );
  XOR U9115 ( .A(n8708), .B(n8709), .Z(n8458) );
  XOR U9116 ( .A(n4963), .B(n4958), .Z(n8709) );
  XOR U9117 ( .A(n8710), .B(n8711), .Z(n4958) );
  XOR U9118 ( .A(n8589), .B(n8531), .Z(n8711) );
  XOR U9119 ( .A(n8712), .B(n8713), .Z(n8531) );
  XNOR U9120 ( .A(n8714), .B(n8477), .Z(n8713) );
  ANDN U9121 ( .B(n8715), .A(n8716), .Z(n8477) );
  ANDN U9122 ( .B(n8717), .A(n8613), .Z(n8714) );
  IV U9123 ( .A(n8718), .Z(n8613) );
  XNOR U9124 ( .A(n8473), .B(n8719), .Z(n8589) );
  XNOR U9125 ( .A(n8720), .B(n8721), .Z(n8719) );
  NANDN U9126 ( .A(n8722), .B(n8667), .Z(n8721) );
  XOR U9127 ( .A(n8712), .B(n8723), .Z(n8553) );
  XNOR U9128 ( .A(n8720), .B(n8724), .Z(n8723) );
  NANDN U9129 ( .A(n8725), .B(n8587), .Z(n8724) );
  OR U9130 ( .A(n8666), .B(n8726), .Z(n8720) );
  XNOR U9131 ( .A(n8587), .B(n8667), .Z(n8666) );
  XNOR U9132 ( .A(n8473), .B(n8727), .Z(n8712) );
  XNOR U9133 ( .A(n8728), .B(n8729), .Z(n8727) );
  NANDN U9134 ( .A(n8618), .B(n8730), .Z(n8729) );
  XOR U9135 ( .A(n8731), .B(n8728), .Z(n8473) );
  NANDN U9136 ( .A(n8732), .B(n8733), .Z(n8728) );
  ANDN U9137 ( .B(n8734), .A(n8735), .Z(n8731) );
  XOR U9138 ( .A(n8614), .B(n8736), .Z(n8552) );
  XOR U9139 ( .A(n8611), .B(n8737), .Z(n8736) );
  NANDN U9140 ( .A(n8738), .B(n8479), .Z(n8737) );
  XOR U9141 ( .A(n8718), .B(n8479), .Z(n8715) );
  XOR U9142 ( .A(n8740), .B(n8616), .Z(n8614) );
  OR U9143 ( .A(n8732), .B(n8741), .Z(n8616) );
  XNOR U9144 ( .A(n8735), .B(n8618), .Z(n8732) );
  XNOR U9145 ( .A(n8667), .B(n8479), .Z(n8618) );
  XOR U9146 ( .A(n8742), .B(n8743), .Z(n8479) );
  NANDN U9147 ( .A(n8744), .B(n8745), .Z(n8743) );
  XOR U9148 ( .A(n8746), .B(n8747), .Z(n8667) );
  NANDN U9149 ( .A(n8744), .B(n8748), .Z(n8747) );
  NOR U9150 ( .A(n8735), .B(n8749), .Z(n8740) );
  XNOR U9151 ( .A(n8718), .B(n8587), .Z(n8735) );
  XNOR U9152 ( .A(n8750), .B(n8746), .Z(n8587) );
  NANDN U9153 ( .A(n8751), .B(n8752), .Z(n8746) );
  XOR U9154 ( .A(n8748), .B(n8753), .Z(n8752) );
  ANDN U9155 ( .B(n8753), .A(n8754), .Z(n8750) );
  XNOR U9156 ( .A(n8755), .B(n8742), .Z(n8718) );
  NANDN U9157 ( .A(n8751), .B(n8756), .Z(n8742) );
  XOR U9158 ( .A(n8757), .B(n8745), .Z(n8756) );
  XNOR U9159 ( .A(n8758), .B(n8759), .Z(n8744) );
  XOR U9160 ( .A(n8760), .B(n8761), .Z(n8759) );
  XNOR U9161 ( .A(n8762), .B(n8763), .Z(n8758) );
  XNOR U9162 ( .A(n8764), .B(n8765), .Z(n8763) );
  ANDN U9163 ( .B(n8757), .A(n8761), .Z(n8764) );
  ANDN U9164 ( .B(n8757), .A(n8754), .Z(n8755) );
  XNOR U9165 ( .A(n8760), .B(n8766), .Z(n8754) );
  XOR U9166 ( .A(n8767), .B(n8765), .Z(n8766) );
  NAND U9167 ( .A(n8768), .B(n8769), .Z(n8765) );
  XNOR U9168 ( .A(n8762), .B(n8745), .Z(n8769) );
  IV U9169 ( .A(n8757), .Z(n8762) );
  XNOR U9170 ( .A(n8748), .B(n8761), .Z(n8768) );
  IV U9171 ( .A(n8753), .Z(n8761) );
  XOR U9172 ( .A(n8770), .B(n8771), .Z(n8753) );
  XNOR U9173 ( .A(n8772), .B(n8773), .Z(n8771) );
  XNOR U9174 ( .A(n8774), .B(n8775), .Z(n8770) );
  ANDN U9175 ( .B(n8612), .A(n8776), .Z(n8774) );
  AND U9176 ( .A(n8745), .B(n8748), .Z(n8767) );
  XNOR U9177 ( .A(n8745), .B(n8748), .Z(n8760) );
  XNOR U9178 ( .A(n8777), .B(n8778), .Z(n8748) );
  XNOR U9179 ( .A(n8779), .B(n8773), .Z(n8778) );
  XOR U9180 ( .A(n8780), .B(n8781), .Z(n8777) );
  XNOR U9181 ( .A(n8782), .B(n8775), .Z(n8781) );
  OR U9182 ( .A(n8716), .B(n8739), .Z(n8775) );
  XNOR U9183 ( .A(n8612), .B(n8783), .Z(n8739) );
  XNOR U9184 ( .A(n8776), .B(n8480), .Z(n8716) );
  ANDN U9185 ( .B(n8784), .A(n8738), .Z(n8782) );
  XNOR U9186 ( .A(n8785), .B(n8786), .Z(n8745) );
  XNOR U9187 ( .A(n8773), .B(n8787), .Z(n8786) );
  XOR U9188 ( .A(n8725), .B(n8780), .Z(n8787) );
  XNOR U9189 ( .A(n8612), .B(n8776), .Z(n8773) );
  XOR U9190 ( .A(n8586), .B(n8788), .Z(n8785) );
  XNOR U9191 ( .A(n8789), .B(n8790), .Z(n8788) );
  ANDN U9192 ( .B(n8791), .A(n8668), .Z(n8789) );
  XNOR U9193 ( .A(n8792), .B(n8793), .Z(n8757) );
  XNOR U9194 ( .A(n8779), .B(n8794), .Z(n8793) );
  XNOR U9195 ( .A(n8722), .B(n8772), .Z(n8794) );
  XOR U9196 ( .A(n8780), .B(n8795), .Z(n8772) );
  XNOR U9197 ( .A(n8796), .B(n8797), .Z(n8795) );
  NAND U9198 ( .A(n8619), .B(n8730), .Z(n8797) );
  XNOR U9199 ( .A(n8798), .B(n8796), .Z(n8780) );
  NANDN U9200 ( .A(n8741), .B(n8733), .Z(n8796) );
  XOR U9201 ( .A(n8734), .B(n8730), .Z(n8733) );
  XNOR U9202 ( .A(n8791), .B(n8480), .Z(n8730) );
  XOR U9203 ( .A(n8749), .B(n8619), .Z(n8741) );
  XNOR U9204 ( .A(n8668), .B(n8783), .Z(n8619) );
  ANDN U9205 ( .B(n8734), .A(n8749), .Z(n8798) );
  XOR U9206 ( .A(n8586), .B(n8612), .Z(n8749) );
  XNOR U9207 ( .A(n8799), .B(n8800), .Z(n8612) );
  XNOR U9208 ( .A(n8801), .B(n8802), .Z(n8800) );
  XOR U9209 ( .A(n8783), .B(n8784), .Z(n8779) );
  IV U9210 ( .A(n8480), .Z(n8784) );
  XOR U9211 ( .A(n8803), .B(n8804), .Z(n8480) );
  XNOR U9212 ( .A(n8805), .B(n8802), .Z(n8804) );
  IV U9213 ( .A(n8738), .Z(n8783) );
  XOR U9214 ( .A(n8802), .B(n8806), .Z(n8738) );
  XNOR U9215 ( .A(n8807), .B(n8808), .Z(n8792) );
  XNOR U9216 ( .A(n8809), .B(n8790), .Z(n8808) );
  OR U9217 ( .A(n8726), .B(n8665), .Z(n8790) );
  XNOR U9218 ( .A(n8586), .B(n8668), .Z(n8665) );
  IV U9219 ( .A(n8807), .Z(n8668) );
  XOR U9220 ( .A(n8725), .B(n8791), .Z(n8726) );
  IV U9221 ( .A(n8722), .Z(n8791) );
  XOR U9222 ( .A(n8717), .B(n8810), .Z(n8722) );
  XNOR U9223 ( .A(n8805), .B(n8799), .Z(n8810) );
  XOR U9224 ( .A(n8811), .B(n8812), .Z(n8799) );
  XOR U9225 ( .A(n7984), .B(n6581), .Z(n8812) );
  XOR U9226 ( .A(n8813), .B(n7940), .Z(n6581) );
  XNOR U9227 ( .A(n7979), .B(n8814), .Z(n8811) );
  XNOR U9228 ( .A(key[938]), .B(n7359), .Z(n8814) );
  XOR U9229 ( .A(n8815), .B(n8816), .Z(n7359) );
  XOR U9230 ( .A(n8817), .B(n8818), .Z(n8816) );
  IV U9231 ( .A(n8776), .Z(n8717) );
  XOR U9232 ( .A(n8803), .B(n8819), .Z(n8776) );
  XOR U9233 ( .A(n8802), .B(n8820), .Z(n8819) );
  NOR U9234 ( .A(n8725), .B(n8586), .Z(n8809) );
  XOR U9235 ( .A(n8803), .B(n8821), .Z(n8725) );
  XOR U9236 ( .A(n8802), .B(n8822), .Z(n8821) );
  XOR U9237 ( .A(n8823), .B(n8824), .Z(n8802) );
  XOR U9238 ( .A(n8586), .B(n6553), .Z(n8824) );
  XOR U9239 ( .A(n8825), .B(n8826), .Z(n6553) );
  XNOR U9240 ( .A(n7951), .B(n8827), .Z(n8823) );
  XNOR U9241 ( .A(key[942]), .B(n7328), .Z(n8827) );
  XOR U9242 ( .A(n6560), .B(n7341), .Z(n7328) );
  XNOR U9243 ( .A(n8815), .B(n8828), .Z(n7966) );
  XOR U9244 ( .A(n8829), .B(n8830), .Z(n8828) );
  XOR U9245 ( .A(n8831), .B(n8832), .Z(n8815) );
  XOR U9246 ( .A(n7953), .B(n7961), .Z(n6560) );
  IV U9247 ( .A(n6555), .Z(n7961) );
  XOR U9248 ( .A(n8833), .B(n8834), .Z(n6555) );
  XOR U9249 ( .A(n8835), .B(n8836), .Z(n7951) );
  IV U9250 ( .A(n8806), .Z(n8803) );
  XOR U9251 ( .A(n8837), .B(n8838), .Z(n8806) );
  XNOR U9252 ( .A(n7958), .B(n7334), .Z(n8838) );
  XNOR U9253 ( .A(n7959), .B(n6558), .Z(n7334) );
  XNOR U9254 ( .A(n8839), .B(n8840), .Z(n6558) );
  XNOR U9255 ( .A(n8841), .B(n8842), .Z(n8840) );
  XNOR U9256 ( .A(n8843), .B(n8844), .Z(n8839) );
  XOR U9257 ( .A(n8845), .B(n8846), .Z(n8844) );
  ANDN U9258 ( .B(n8847), .A(n8848), .Z(n8846) );
  XNOR U9259 ( .A(n8849), .B(n8850), .Z(n7958) );
  XOR U9260 ( .A(n8851), .B(n8852), .Z(n8850) );
  XNOR U9261 ( .A(n8853), .B(n8854), .Z(n8849) );
  XOR U9262 ( .A(n8855), .B(n8856), .Z(n8854) );
  ANDN U9263 ( .B(n8857), .A(n8858), .Z(n8856) );
  XNOR U9264 ( .A(n7953), .B(n8859), .Z(n8837) );
  XNOR U9265 ( .A(key[941]), .B(n7330), .Z(n8859) );
  XOR U9266 ( .A(n8829), .B(n8818), .Z(n7330) );
  XNOR U9267 ( .A(n8860), .B(n8861), .Z(n8818) );
  XNOR U9268 ( .A(n8862), .B(n8863), .Z(n8861) );
  ANDN U9269 ( .B(n8864), .A(n8865), .Z(n8862) );
  XNOR U9270 ( .A(n8866), .B(n8867), .Z(n7953) );
  XOR U9271 ( .A(n8868), .B(n8869), .Z(n8807) );
  XNOR U9272 ( .A(n8822), .B(n8820), .Z(n8869) );
  XNOR U9273 ( .A(n8870), .B(n8871), .Z(n8820) );
  XNOR U9274 ( .A(n7955), .B(n7342), .Z(n8871) );
  XNOR U9275 ( .A(n8826), .B(n7950), .Z(n7342) );
  XNOR U9276 ( .A(n8872), .B(n8873), .Z(n7950) );
  XNOR U9277 ( .A(n8874), .B(n8842), .Z(n8873) );
  XNOR U9278 ( .A(n8875), .B(n8876), .Z(n8842) );
  XNOR U9279 ( .A(n8877), .B(n8878), .Z(n8876) );
  NANDN U9280 ( .A(n8879), .B(n8880), .Z(n8878) );
  XOR U9281 ( .A(n8881), .B(n8833), .Z(n8872) );
  IV U9282 ( .A(n7967), .Z(n8826) );
  XNOR U9283 ( .A(n8882), .B(n8883), .Z(n7967) );
  XNOR U9284 ( .A(n8866), .B(n8884), .Z(n8883) );
  XNOR U9285 ( .A(n8885), .B(n8886), .Z(n8882) );
  XNOR U9286 ( .A(n8887), .B(n8888), .Z(n7955) );
  XOR U9287 ( .A(n8889), .B(n8852), .Z(n8888) );
  XNOR U9288 ( .A(n8890), .B(n8891), .Z(n8852) );
  XNOR U9289 ( .A(n8892), .B(n8893), .Z(n8891) );
  NANDN U9290 ( .A(n8894), .B(n8895), .Z(n8893) );
  XOR U9291 ( .A(n8896), .B(n8835), .Z(n8887) );
  XNOR U9292 ( .A(key[943]), .B(n7364), .Z(n8870) );
  XNOR U9293 ( .A(n6567), .B(n6590), .Z(n7364) );
  XNOR U9294 ( .A(n8897), .B(n8898), .Z(n8822) );
  XNOR U9295 ( .A(n7346), .B(n6570), .Z(n8898) );
  XOR U9296 ( .A(n8825), .B(n7959), .Z(n6570) );
  XOR U9297 ( .A(n8899), .B(n8900), .Z(n7959) );
  XNOR U9298 ( .A(n8901), .B(n8884), .Z(n8900) );
  XNOR U9299 ( .A(n8902), .B(n8903), .Z(n8884) );
  XNOR U9300 ( .A(n8904), .B(n8905), .Z(n8903) );
  NANDN U9301 ( .A(n8906), .B(n8907), .Z(n8905) );
  XNOR U9302 ( .A(n8908), .B(n8909), .Z(n8899) );
  XNOR U9303 ( .A(n8910), .B(n8911), .Z(n8909) );
  ANDN U9304 ( .B(n8912), .A(n8913), .Z(n8911) );
  XNOR U9305 ( .A(n7973), .B(n6572), .Z(n7346) );
  XNOR U9306 ( .A(n8843), .B(n6544), .Z(n6572) );
  IV U9307 ( .A(n8813), .Z(n6544) );
  XNOR U9308 ( .A(n8914), .B(n8874), .Z(n8813) );
  XNOR U9309 ( .A(n7348), .B(n8915), .Z(n8897) );
  XNOR U9310 ( .A(key[940]), .B(n7971), .Z(n8915) );
  XNOR U9311 ( .A(n7943), .B(n8851), .Z(n7971) );
  IV U9312 ( .A(n7979), .Z(n7943) );
  XOR U9313 ( .A(n8916), .B(n8889), .Z(n7979) );
  XOR U9314 ( .A(n6590), .B(n7336), .Z(n7348) );
  XNOR U9315 ( .A(n8917), .B(n8918), .Z(n7336) );
  XOR U9316 ( .A(n8919), .B(n8830), .Z(n8918) );
  XNOR U9317 ( .A(n8920), .B(n8921), .Z(n8830) );
  XNOR U9318 ( .A(n8922), .B(n8923), .Z(n8921) );
  OR U9319 ( .A(n8924), .B(n8925), .Z(n8923) );
  XNOR U9320 ( .A(n8926), .B(n8927), .Z(n8917) );
  XOR U9321 ( .A(n8863), .B(n8928), .Z(n8927) );
  ANDN U9322 ( .B(n8929), .A(n8930), .Z(n8928) );
  ANDN U9323 ( .B(n8931), .A(n8932), .Z(n8863) );
  XNOR U9324 ( .A(n8586), .B(n8801), .Z(n8868) );
  XOR U9325 ( .A(n8933), .B(n8934), .Z(n8801) );
  XNOR U9326 ( .A(n8805), .B(n8935), .Z(n8934) );
  XOR U9327 ( .A(n7941), .B(n6577), .Z(n8935) );
  XOR U9328 ( .A(n8825), .B(n7973), .Z(n6577) );
  XOR U9329 ( .A(n8908), .B(n7940), .Z(n7973) );
  XNOR U9330 ( .A(n8936), .B(n8937), .Z(n7941) );
  XOR U9331 ( .A(n8889), .B(n8836), .Z(n8937) );
  XNOR U9332 ( .A(n8938), .B(n8939), .Z(n8836) );
  XNOR U9333 ( .A(n8940), .B(n8855), .Z(n8939) );
  NOR U9334 ( .A(n8941), .B(n8942), .Z(n8855) );
  ANDN U9335 ( .B(n8943), .A(n8944), .Z(n8940) );
  XOR U9336 ( .A(n8896), .B(n8945), .Z(n8936) );
  XOR U9337 ( .A(n8946), .B(n8947), .Z(n8805) );
  XOR U9338 ( .A(n6588), .B(n7940), .Z(n8947) );
  XOR U9339 ( .A(n8948), .B(n8885), .Z(n7940) );
  XOR U9340 ( .A(n7980), .B(n7987), .Z(n6588) );
  IV U9341 ( .A(n6580), .Z(n7987) );
  XNOR U9342 ( .A(n8881), .B(n8833), .Z(n8949) );
  XOR U9343 ( .A(n8950), .B(n8951), .Z(n8833) );
  XNOR U9344 ( .A(n8952), .B(n8953), .Z(n8946) );
  XNOR U9345 ( .A(key[937]), .B(n7982), .Z(n8953) );
  XOR U9346 ( .A(n8889), .B(n8954), .Z(n7982) );
  XNOR U9347 ( .A(n8896), .B(n8835), .Z(n8954) );
  XOR U9348 ( .A(n8955), .B(n8945), .Z(n8835) );
  XOR U9349 ( .A(n8853), .B(n8956), .Z(n8945) );
  XNOR U9350 ( .A(n8957), .B(n8958), .Z(n8956) );
  NANDN U9351 ( .A(n8959), .B(n8960), .Z(n8958) );
  XNOR U9352 ( .A(n8957), .B(n8962), .Z(n8961) );
  NAND U9353 ( .A(n8963), .B(n8895), .Z(n8962) );
  OR U9354 ( .A(n8964), .B(n8965), .Z(n8957) );
  XNOR U9355 ( .A(n8853), .B(n8966), .Z(n8938) );
  XNOR U9356 ( .A(n8967), .B(n8968), .Z(n8966) );
  OR U9357 ( .A(n8969), .B(n8970), .Z(n8968) );
  XOR U9358 ( .A(n8971), .B(n8967), .Z(n8853) );
  OR U9359 ( .A(n8972), .B(n8973), .Z(n8967) );
  ANDN U9360 ( .B(n8974), .A(n8975), .Z(n8971) );
  XOR U9361 ( .A(n8976), .B(n8977), .Z(n8889) );
  XOR U9362 ( .A(n8978), .B(n8979), .Z(n8977) );
  NANDN U9363 ( .A(n8980), .B(n8857), .Z(n8979) );
  XOR U9364 ( .A(n7355), .B(n8981), .Z(n8933) );
  XNOR U9365 ( .A(key[939]), .B(n7361), .Z(n8981) );
  XNOR U9366 ( .A(n6590), .B(n7350), .Z(n7361) );
  XOR U9367 ( .A(n8926), .B(n7321), .Z(n7350) );
  IV U9368 ( .A(n8952), .Z(n7321) );
  XOR U9369 ( .A(n8982), .B(n8831), .Z(n8952) );
  XOR U9370 ( .A(n8983), .B(n8926), .Z(n6590) );
  XNOR U9371 ( .A(n8920), .B(n8984), .Z(n8926) );
  XNOR U9372 ( .A(n8985), .B(n8986), .Z(n8984) );
  ANDN U9373 ( .B(n8864), .A(n8987), .Z(n8985) );
  XNOR U9374 ( .A(n8988), .B(n8989), .Z(n8920) );
  XNOR U9375 ( .A(n8990), .B(n8991), .Z(n8989) );
  NAND U9376 ( .A(n8992), .B(n8993), .Z(n8991) );
  IV U9377 ( .A(n6543), .Z(n7355) );
  XOR U9378 ( .A(n7984), .B(n6585), .Z(n6543) );
  XNOR U9379 ( .A(n8994), .B(n8995), .Z(n6585) );
  XNOR U9380 ( .A(n8874), .B(n8834), .Z(n8995) );
  XNOR U9381 ( .A(n8996), .B(n8997), .Z(n8834) );
  XNOR U9382 ( .A(n8998), .B(n8845), .Z(n8997) );
  ANDN U9383 ( .B(n8999), .A(n9000), .Z(n8845) );
  ANDN U9384 ( .B(n9001), .A(n9002), .Z(n8998) );
  XOR U9385 ( .A(n9003), .B(n9004), .Z(n8874) );
  XNOR U9386 ( .A(n9005), .B(n9006), .Z(n9004) );
  NANDN U9387 ( .A(n9007), .B(n8847), .Z(n9006) );
  XNOR U9388 ( .A(n8881), .B(n8951), .Z(n8994) );
  XNOR U9389 ( .A(n8841), .B(n9008), .Z(n8951) );
  XNOR U9390 ( .A(n9009), .B(n9010), .Z(n9008) );
  NANDN U9391 ( .A(n9011), .B(n9012), .Z(n9010) );
  XNOR U9392 ( .A(n9009), .B(n9014), .Z(n9013) );
  NANDN U9393 ( .A(n9015), .B(n8880), .Z(n9014) );
  OR U9394 ( .A(n9016), .B(n9017), .Z(n9009) );
  XNOR U9395 ( .A(n8841), .B(n9018), .Z(n8996) );
  XNOR U9396 ( .A(n9019), .B(n9020), .Z(n9018) );
  NANDN U9397 ( .A(n9021), .B(n9022), .Z(n9020) );
  XOR U9398 ( .A(n9023), .B(n9019), .Z(n8841) );
  NANDN U9399 ( .A(n9024), .B(n9025), .Z(n9019) );
  ANDN U9400 ( .B(n9026), .A(n9027), .Z(n9023) );
  XOR U9401 ( .A(n9028), .B(n9029), .Z(n7984) );
  XNOR U9402 ( .A(n9030), .B(n8867), .Z(n9029) );
  XNOR U9403 ( .A(n9031), .B(n9032), .Z(n8867) );
  XOR U9404 ( .A(n9033), .B(n8910), .Z(n9032) );
  NANDN U9405 ( .A(n9034), .B(n9035), .Z(n8910) );
  ANDN U9406 ( .B(n9036), .A(n9037), .Z(n9033) );
  XOR U9407 ( .A(n8885), .B(n9038), .Z(n9028) );
  XNOR U9408 ( .A(n9039), .B(n9040), .Z(n8586) );
  XOR U9409 ( .A(n7980), .B(n6589), .Z(n9040) );
  XOR U9410 ( .A(n7365), .B(n7954), .Z(n6589) );
  XOR U9411 ( .A(n8955), .B(n8851), .Z(n7954) );
  XOR U9412 ( .A(n8890), .B(n9041), .Z(n8851) );
  XNOR U9413 ( .A(n9042), .B(n8978), .Z(n9041) );
  NOR U9414 ( .A(n8941), .B(n9043), .Z(n8978) );
  XNOR U9415 ( .A(n8943), .B(n8857), .Z(n8941) );
  XNOR U9416 ( .A(n8976), .B(n9045), .Z(n8890) );
  XNOR U9417 ( .A(n9046), .B(n9047), .Z(n9045) );
  NANDN U9418 ( .A(n8969), .B(n9048), .Z(n9047) );
  IV U9419 ( .A(n8916), .Z(n8955) );
  XNOR U9420 ( .A(n8976), .B(n9049), .Z(n8916) );
  XOR U9421 ( .A(n9050), .B(n8892), .Z(n9049) );
  OR U9422 ( .A(n9051), .B(n8964), .Z(n8892) );
  XNOR U9423 ( .A(n8895), .B(n8960), .Z(n8964) );
  ANDN U9424 ( .B(n8960), .A(n9052), .Z(n9050) );
  XOR U9425 ( .A(n9053), .B(n9046), .Z(n8976) );
  OR U9426 ( .A(n8972), .B(n9054), .Z(n9046) );
  XOR U9427 ( .A(n8974), .B(n8969), .Z(n8972) );
  XNOR U9428 ( .A(n8960), .B(n8857), .Z(n8969) );
  XNOR U9429 ( .A(n9055), .B(n9056), .Z(n8857) );
  NANDN U9430 ( .A(n9057), .B(n9058), .Z(n9056) );
  XOR U9431 ( .A(n9059), .B(n9060), .Z(n8960) );
  NANDN U9432 ( .A(n9057), .B(n9061), .Z(n9060) );
  XOR U9433 ( .A(n8943), .B(n8895), .Z(n8974) );
  XNOR U9434 ( .A(n9063), .B(n9059), .Z(n8895) );
  NANDN U9435 ( .A(n9064), .B(n9065), .Z(n9059) );
  XOR U9436 ( .A(n9061), .B(n9066), .Z(n9065) );
  ANDN U9437 ( .B(n9066), .A(n9067), .Z(n9063) );
  XOR U9438 ( .A(n9068), .B(n9055), .Z(n8943) );
  ANDN U9439 ( .B(n9069), .A(n9064), .Z(n9055) );
  XNOR U9440 ( .A(n9070), .B(n9071), .Z(n9057) );
  XOR U9441 ( .A(n9072), .B(n9073), .Z(n9071) );
  XNOR U9442 ( .A(n9074), .B(n9075), .Z(n9070) );
  XNOR U9443 ( .A(n9076), .B(n9077), .Z(n9075) );
  ANDN U9444 ( .B(n9078), .A(n9073), .Z(n9076) );
  XOR U9445 ( .A(n9078), .B(n9058), .Z(n9069) );
  ANDN U9446 ( .B(n9078), .A(n9067), .Z(n9068) );
  XNOR U9447 ( .A(n9072), .B(n9079), .Z(n9067) );
  XOR U9448 ( .A(n9080), .B(n9077), .Z(n9079) );
  NAND U9449 ( .A(n9081), .B(n9082), .Z(n9077) );
  XNOR U9450 ( .A(n9074), .B(n9058), .Z(n9082) );
  IV U9451 ( .A(n9078), .Z(n9074) );
  XNOR U9452 ( .A(n9061), .B(n9073), .Z(n9081) );
  IV U9453 ( .A(n9066), .Z(n9073) );
  XOR U9454 ( .A(n9083), .B(n9084), .Z(n9066) );
  XNOR U9455 ( .A(n9085), .B(n9086), .Z(n9084) );
  XNOR U9456 ( .A(n9087), .B(n9088), .Z(n9083) );
  ANDN U9457 ( .B(n9044), .A(n8944), .Z(n9087) );
  AND U9458 ( .A(n9058), .B(n9061), .Z(n9080) );
  XNOR U9459 ( .A(n9058), .B(n9061), .Z(n9072) );
  XNOR U9460 ( .A(n9089), .B(n9090), .Z(n9061) );
  XNOR U9461 ( .A(n9091), .B(n9086), .Z(n9090) );
  XOR U9462 ( .A(n9092), .B(n9093), .Z(n9089) );
  XNOR U9463 ( .A(n9094), .B(n9088), .Z(n9093) );
  OR U9464 ( .A(n8942), .B(n9043), .Z(n9088) );
  XNOR U9465 ( .A(n9044), .B(n9125), .Z(n9043) );
  XNOR U9466 ( .A(n8944), .B(n8858), .Z(n8942) );
  ANDN U9467 ( .B(n9095), .A(n8980), .Z(n9094) );
  XNOR U9468 ( .A(n9096), .B(n9097), .Z(n9058) );
  XNOR U9469 ( .A(n9086), .B(n9098), .Z(n9097) );
  XNOR U9470 ( .A(n8963), .B(n9092), .Z(n9098) );
  XNOR U9471 ( .A(n8944), .B(n9044), .Z(n9086) );
  XOR U9472 ( .A(n8894), .B(n9099), .Z(n9096) );
  XNOR U9473 ( .A(n9100), .B(n9101), .Z(n9099) );
  ANDN U9474 ( .B(n9102), .A(n9052), .Z(n9100) );
  XNOR U9475 ( .A(n9103), .B(n9104), .Z(n9078) );
  XNOR U9476 ( .A(n9091), .B(n9105), .Z(n9104) );
  XNOR U9477 ( .A(n9106), .B(n9085), .Z(n9105) );
  XOR U9478 ( .A(n9092), .B(n9107), .Z(n9085) );
  XNOR U9479 ( .A(n9108), .B(n9109), .Z(n9107) );
  NANDN U9480 ( .A(n8970), .B(n9048), .Z(n9109) );
  XNOR U9481 ( .A(n9110), .B(n9108), .Z(n9092) );
  OR U9482 ( .A(n9054), .B(n8973), .Z(n9108) );
  XOR U9483 ( .A(n9111), .B(n8970), .Z(n8973) );
  XNOR U9484 ( .A(n9095), .B(n9102), .Z(n8970) );
  IV U9485 ( .A(n8858), .Z(n9095) );
  XNOR U9486 ( .A(n9062), .B(n9048), .Z(n9054) );
  XNOR U9487 ( .A(n9052), .B(n9125), .Z(n9048) );
  ANDN U9488 ( .B(n9062), .A(n8975), .Z(n9110) );
  IV U9489 ( .A(n9111), .Z(n8975) );
  XOR U9490 ( .A(n9112), .B(n8963), .Z(n9111) );
  XOR U9491 ( .A(n8858), .B(n8980), .Z(n9091) );
  XOR U9492 ( .A(n9113), .B(n9114), .Z(n8980) );
  XOR U9493 ( .A(n9115), .B(n9116), .Z(n8858) );
  XOR U9494 ( .A(n9117), .B(n9114), .Z(n9116) );
  XNOR U9495 ( .A(n8959), .B(n9118), .Z(n9103) );
  XNOR U9496 ( .A(n9119), .B(n9101), .Z(n9118) );
  OR U9497 ( .A(n8965), .B(n9051), .Z(n9101) );
  XNOR U9498 ( .A(n8894), .B(n9052), .Z(n9051) );
  IV U9499 ( .A(n9106), .Z(n9052) );
  XOR U9500 ( .A(n9120), .B(n9121), .Z(n9106) );
  XNOR U9501 ( .A(n9122), .B(n9123), .Z(n9121) );
  XNOR U9502 ( .A(n8894), .B(n9124), .Z(n9120) );
  XNOR U9503 ( .A(n8963), .B(n9102), .Z(n8965) );
  IV U9504 ( .A(n8959), .Z(n9102) );
  ANDN U9505 ( .B(n8963), .A(n8894), .Z(n9119) );
  XOR U9506 ( .A(n9122), .B(n9125), .Z(n8963) );
  XOR U9507 ( .A(n9126), .B(n9127), .Z(n9122) );
  XNOR U9508 ( .A(n9128), .B(n9129), .Z(n9127) );
  XNOR U9509 ( .A(key[788]), .B(n9130), .Z(n9126) );
  XNOR U9510 ( .A(n9131), .B(n9132), .Z(n8959) );
  XOR U9511 ( .A(n8944), .B(n9115), .Z(n9132) );
  IV U9512 ( .A(n9112), .Z(n8944) );
  XOR U9513 ( .A(n9124), .B(n9125), .Z(n9112) );
  XNOR U9514 ( .A(n9113), .B(n9114), .Z(n9125) );
  IV U9515 ( .A(n9117), .Z(n9113) );
  XNOR U9516 ( .A(n9133), .B(n9134), .Z(n9117) );
  XNOR U9517 ( .A(n9135), .B(n9136), .Z(n9134) );
  XNOR U9518 ( .A(key[789]), .B(n9137), .Z(n9133) );
  XOR U9519 ( .A(n9138), .B(n9139), .Z(n9124) );
  XOR U9520 ( .A(n9140), .B(n9141), .Z(n9139) );
  XOR U9521 ( .A(key[791]), .B(n9142), .Z(n9138) );
  XNOR U9522 ( .A(n8894), .B(n9044), .Z(n9062) );
  XNOR U9523 ( .A(n9123), .B(n9143), .Z(n9044) );
  XNOR U9524 ( .A(n9114), .B(n9131), .Z(n9143) );
  XOR U9525 ( .A(n9144), .B(n9145), .Z(n9131) );
  XOR U9526 ( .A(n9146), .B(n9147), .Z(n9145) );
  XNOR U9527 ( .A(key[786]), .B(n9148), .Z(n9144) );
  XOR U9528 ( .A(n9149), .B(n9150), .Z(n9114) );
  XNOR U9529 ( .A(n8894), .B(n9151), .Z(n9150) );
  XNOR U9530 ( .A(n9152), .B(n9153), .Z(n9149) );
  XNOR U9531 ( .A(key[790]), .B(n9154), .Z(n9153) );
  XOR U9532 ( .A(n9155), .B(n9156), .Z(n9123) );
  XNOR U9533 ( .A(n9157), .B(n9158), .Z(n9156) );
  XOR U9534 ( .A(n9159), .B(n9160), .Z(n9158) );
  XNOR U9535 ( .A(n9161), .B(n9162), .Z(n9155) );
  XOR U9536 ( .A(key[787]), .B(n9115), .Z(n9162) );
  XNOR U9537 ( .A(n9163), .B(n9164), .Z(n9115) );
  XOR U9538 ( .A(n9165), .B(n9166), .Z(n9164) );
  XNOR U9539 ( .A(key[785]), .B(n9167), .Z(n9163) );
  XNOR U9540 ( .A(n9168), .B(n9169), .Z(n8894) );
  XOR U9541 ( .A(n9170), .B(n9171), .Z(n9169) );
  XNOR U9542 ( .A(key[784]), .B(n9172), .Z(n9168) );
  XOR U9543 ( .A(n8843), .B(n8950), .Z(n7365) );
  IV U9544 ( .A(n8914), .Z(n8950) );
  XOR U9545 ( .A(n9174), .B(n8877), .Z(n9173) );
  OR U9546 ( .A(n9016), .B(n9175), .Z(n8877) );
  XNOR U9547 ( .A(n8880), .B(n9012), .Z(n9016) );
  ANDN U9548 ( .B(n9012), .A(n9176), .Z(n9174) );
  XNOR U9549 ( .A(n8875), .B(n9177), .Z(n8843) );
  XOR U9550 ( .A(n9178), .B(n9005), .Z(n9177) );
  XOR U9551 ( .A(n9180), .B(n8847), .Z(n8999) );
  ANDN U9552 ( .B(n9181), .A(n9002), .Z(n9178) );
  IV U9553 ( .A(n9180), .Z(n9002) );
  XOR U9554 ( .A(n9003), .B(n9182), .Z(n8875) );
  XNOR U9555 ( .A(n9183), .B(n9184), .Z(n9182) );
  NANDN U9556 ( .A(n9021), .B(n9185), .Z(n9184) );
  XNOR U9557 ( .A(n9186), .B(n9183), .Z(n9003) );
  OR U9558 ( .A(n9024), .B(n9187), .Z(n9183) );
  XNOR U9559 ( .A(n9027), .B(n9021), .Z(n9024) );
  XNOR U9560 ( .A(n9012), .B(n8847), .Z(n9021) );
  XOR U9561 ( .A(n9188), .B(n9189), .Z(n8847) );
  NANDN U9562 ( .A(n9190), .B(n9191), .Z(n9189) );
  XOR U9563 ( .A(n9192), .B(n9193), .Z(n9012) );
  NANDN U9564 ( .A(n9190), .B(n9194), .Z(n9193) );
  NOR U9565 ( .A(n9027), .B(n9195), .Z(n9186) );
  XNOR U9566 ( .A(n9180), .B(n8880), .Z(n9027) );
  XNOR U9567 ( .A(n9196), .B(n9192), .Z(n8880) );
  NANDN U9568 ( .A(n9197), .B(n9198), .Z(n9192) );
  XOR U9569 ( .A(n9194), .B(n9199), .Z(n9198) );
  ANDN U9570 ( .B(n9199), .A(n9200), .Z(n9196) );
  XNOR U9571 ( .A(n9201), .B(n9188), .Z(n9180) );
  NANDN U9572 ( .A(n9197), .B(n9202), .Z(n9188) );
  XOR U9573 ( .A(n9203), .B(n9191), .Z(n9202) );
  XNOR U9574 ( .A(n9204), .B(n9205), .Z(n9190) );
  XOR U9575 ( .A(n9206), .B(n9207), .Z(n9205) );
  XNOR U9576 ( .A(n9208), .B(n9209), .Z(n9204) );
  XNOR U9577 ( .A(n9210), .B(n9211), .Z(n9209) );
  ANDN U9578 ( .B(n9203), .A(n9207), .Z(n9210) );
  ANDN U9579 ( .B(n9203), .A(n9200), .Z(n9201) );
  XNOR U9580 ( .A(n9206), .B(n9212), .Z(n9200) );
  XOR U9581 ( .A(n9213), .B(n9211), .Z(n9212) );
  NAND U9582 ( .A(n9214), .B(n9215), .Z(n9211) );
  XNOR U9583 ( .A(n9208), .B(n9191), .Z(n9215) );
  IV U9584 ( .A(n9203), .Z(n9208) );
  XNOR U9585 ( .A(n9194), .B(n9207), .Z(n9214) );
  IV U9586 ( .A(n9199), .Z(n9207) );
  XOR U9587 ( .A(n9216), .B(n9217), .Z(n9199) );
  XNOR U9588 ( .A(n9218), .B(n9219), .Z(n9217) );
  XNOR U9589 ( .A(n9220), .B(n9221), .Z(n9216) );
  ANDN U9590 ( .B(n9181), .A(n9222), .Z(n9220) );
  AND U9591 ( .A(n9191), .B(n9194), .Z(n9213) );
  XNOR U9592 ( .A(n9191), .B(n9194), .Z(n9206) );
  XNOR U9593 ( .A(n9223), .B(n9224), .Z(n9194) );
  XNOR U9594 ( .A(n9225), .B(n9219), .Z(n9224) );
  XOR U9595 ( .A(n9226), .B(n9227), .Z(n9223) );
  XNOR U9596 ( .A(n9228), .B(n9221), .Z(n9227) );
  OR U9597 ( .A(n9000), .B(n9179), .Z(n9221) );
  XNOR U9598 ( .A(n9181), .B(n9229), .Z(n9179) );
  XNOR U9599 ( .A(n9222), .B(n8848), .Z(n9000) );
  ANDN U9600 ( .B(n9230), .A(n9007), .Z(n9228) );
  XNOR U9601 ( .A(n9231), .B(n9232), .Z(n9191) );
  XNOR U9602 ( .A(n9219), .B(n9233), .Z(n9232) );
  XOR U9603 ( .A(n9015), .B(n9226), .Z(n9233) );
  XNOR U9604 ( .A(n9181), .B(n9222), .Z(n9219) );
  XOR U9605 ( .A(n8879), .B(n9234), .Z(n9231) );
  XNOR U9606 ( .A(n9235), .B(n9236), .Z(n9234) );
  ANDN U9607 ( .B(n9237), .A(n9176), .Z(n9235) );
  XNOR U9608 ( .A(n9238), .B(n9239), .Z(n9203) );
  XNOR U9609 ( .A(n9225), .B(n9240), .Z(n9239) );
  XNOR U9610 ( .A(n9011), .B(n9218), .Z(n9240) );
  XOR U9611 ( .A(n9226), .B(n9241), .Z(n9218) );
  XNOR U9612 ( .A(n9242), .B(n9243), .Z(n9241) );
  NAND U9613 ( .A(n9185), .B(n9022), .Z(n9243) );
  XNOR U9614 ( .A(n9244), .B(n9242), .Z(n9226) );
  NANDN U9615 ( .A(n9187), .B(n9025), .Z(n9242) );
  XOR U9616 ( .A(n9026), .B(n9022), .Z(n9025) );
  XNOR U9617 ( .A(n9237), .B(n8848), .Z(n9022) );
  XOR U9618 ( .A(n9195), .B(n9185), .Z(n9187) );
  XNOR U9619 ( .A(n9176), .B(n9229), .Z(n9185) );
  ANDN U9620 ( .B(n9026), .A(n9195), .Z(n9244) );
  XOR U9621 ( .A(n8879), .B(n9181), .Z(n9195) );
  XNOR U9622 ( .A(n9245), .B(n9246), .Z(n9181) );
  XNOR U9623 ( .A(n9247), .B(n9248), .Z(n9246) );
  XOR U9624 ( .A(n9229), .B(n9230), .Z(n9225) );
  IV U9625 ( .A(n8848), .Z(n9230) );
  XOR U9626 ( .A(n9249), .B(n9250), .Z(n8848) );
  XNOR U9627 ( .A(n9251), .B(n9248), .Z(n9250) );
  IV U9628 ( .A(n9007), .Z(n9229) );
  XOR U9629 ( .A(n9248), .B(n9252), .Z(n9007) );
  XNOR U9630 ( .A(n9253), .B(n9254), .Z(n9238) );
  XNOR U9631 ( .A(n9255), .B(n9236), .Z(n9254) );
  OR U9632 ( .A(n9017), .B(n9175), .Z(n9236) );
  XNOR U9633 ( .A(n8879), .B(n9176), .Z(n9175) );
  IV U9634 ( .A(n9253), .Z(n9176) );
  XOR U9635 ( .A(n9015), .B(n9237), .Z(n9017) );
  IV U9636 ( .A(n9011), .Z(n9237) );
  XOR U9637 ( .A(n9001), .B(n9256), .Z(n9011) );
  XNOR U9638 ( .A(n9251), .B(n9245), .Z(n9256) );
  XOR U9639 ( .A(n9257), .B(n9258), .Z(n9245) );
  XOR U9640 ( .A(n9259), .B(n9260), .Z(n9258) );
  XOR U9641 ( .A(n9261), .B(n9262), .Z(n9257) );
  XNOR U9642 ( .A(key[826]), .B(n9263), .Z(n9262) );
  IV U9643 ( .A(n9222), .Z(n9001) );
  XOR U9644 ( .A(n9249), .B(n9264), .Z(n9222) );
  XOR U9645 ( .A(n9248), .B(n9265), .Z(n9264) );
  NOR U9646 ( .A(n9015), .B(n8879), .Z(n9255) );
  XOR U9647 ( .A(n9249), .B(n9266), .Z(n9015) );
  XOR U9648 ( .A(n9248), .B(n9267), .Z(n9266) );
  XOR U9649 ( .A(n9268), .B(n9269), .Z(n9248) );
  XOR U9650 ( .A(n9270), .B(n9271), .Z(n9269) );
  XNOR U9651 ( .A(n9272), .B(n9273), .Z(n9268) );
  XOR U9652 ( .A(key[830]), .B(n8879), .Z(n9273) );
  IV U9653 ( .A(n9252), .Z(n9249) );
  XOR U9654 ( .A(n9274), .B(n9275), .Z(n9252) );
  XNOR U9655 ( .A(n9276), .B(n9277), .Z(n9275) );
  XNOR U9656 ( .A(n9278), .B(n9279), .Z(n9274) );
  XNOR U9657 ( .A(key[829]), .B(n9280), .Z(n9279) );
  XOR U9658 ( .A(n9281), .B(n9282), .Z(n9253) );
  XNOR U9659 ( .A(n9267), .B(n9265), .Z(n9282) );
  XNOR U9660 ( .A(n9283), .B(n9284), .Z(n9265) );
  XNOR U9661 ( .A(n9285), .B(n9286), .Z(n9284) );
  XNOR U9662 ( .A(key[831]), .B(n9287), .Z(n9283) );
  XNOR U9663 ( .A(n9288), .B(n9289), .Z(n9267) );
  XNOR U9664 ( .A(n9290), .B(n9291), .Z(n9289) );
  XNOR U9665 ( .A(n9292), .B(n9293), .Z(n9288) );
  XNOR U9666 ( .A(key[828]), .B(n9294), .Z(n9293) );
  XNOR U9667 ( .A(n8879), .B(n9247), .Z(n9281) );
  XOR U9668 ( .A(n9295), .B(n9296), .Z(n9247) );
  XNOR U9669 ( .A(n9297), .B(n9298), .Z(n9296) );
  XNOR U9670 ( .A(n9251), .B(n9299), .Z(n9298) );
  XOR U9671 ( .A(n9300), .B(n9301), .Z(n9251) );
  XNOR U9672 ( .A(n9302), .B(n9303), .Z(n9301) );
  XOR U9673 ( .A(n9304), .B(n9305), .Z(n9300) );
  XNOR U9674 ( .A(key[825]), .B(n9306), .Z(n9305) );
  XNOR U9675 ( .A(n9307), .B(n9308), .Z(n9295) );
  XNOR U9676 ( .A(key[827]), .B(n9309), .Z(n9308) );
  XNOR U9677 ( .A(n9310), .B(n9311), .Z(n8879) );
  XOR U9678 ( .A(n9312), .B(n9313), .Z(n9311) );
  XNOR U9679 ( .A(n9314), .B(n9315), .Z(n9310) );
  XOR U9680 ( .A(key[824]), .B(n9316), .Z(n9315) );
  XNOR U9681 ( .A(n8866), .B(n9317), .Z(n7980) );
  XOR U9682 ( .A(n8885), .B(n8886), .Z(n9317) );
  IV U9683 ( .A(n9038), .Z(n8886) );
  XOR U9684 ( .A(n9031), .B(n9318), .Z(n9038) );
  XNOR U9685 ( .A(n9319), .B(n9320), .Z(n9318) );
  NANDN U9686 ( .A(n9321), .B(n8907), .Z(n9320) );
  XNOR U9687 ( .A(n8901), .B(n9322), .Z(n9031) );
  XNOR U9688 ( .A(n9323), .B(n9324), .Z(n9322) );
  NANDN U9689 ( .A(n9325), .B(n9326), .Z(n9324) );
  XOR U9690 ( .A(n9327), .B(n9328), .Z(n8885) );
  XNOR U9691 ( .A(n9329), .B(n9330), .Z(n9328) );
  NANDN U9692 ( .A(n9331), .B(n8912), .Z(n9330) );
  XOR U9693 ( .A(n8948), .B(n9030), .Z(n8866) );
  XNOR U9694 ( .A(n8901), .B(n9332), .Z(n9030) );
  XNOR U9695 ( .A(n9319), .B(n9333), .Z(n9332) );
  NANDN U9696 ( .A(n9334), .B(n9335), .Z(n9333) );
  OR U9697 ( .A(n9336), .B(n9337), .Z(n9319) );
  XOR U9698 ( .A(n9338), .B(n9323), .Z(n8901) );
  NANDN U9699 ( .A(n9339), .B(n9340), .Z(n9323) );
  ANDN U9700 ( .B(n9341), .A(n9342), .Z(n9338) );
  XNOR U9701 ( .A(n7358), .B(n9343), .Z(n9039) );
  XOR U9702 ( .A(key[936]), .B(n8825), .Z(n9343) );
  IV U9703 ( .A(n6567), .Z(n8825) );
  XOR U9704 ( .A(n8908), .B(n8948), .Z(n6567) );
  XOR U9705 ( .A(n9327), .B(n9344), .Z(n8948) );
  XOR U9706 ( .A(n9345), .B(n8904), .Z(n9344) );
  OR U9707 ( .A(n9346), .B(n9336), .Z(n8904) );
  XNOR U9708 ( .A(n8907), .B(n9335), .Z(n9336) );
  ANDN U9709 ( .B(n9335), .A(n9347), .Z(n9345) );
  XNOR U9710 ( .A(n8902), .B(n9348), .Z(n8908) );
  XOR U9711 ( .A(n9349), .B(n9329), .Z(n9348) );
  NANDN U9712 ( .A(n9350), .B(n9035), .Z(n9329) );
  XNOR U9713 ( .A(n9037), .B(n8912), .Z(n9035) );
  ANDN U9714 ( .B(n9351), .A(n9037), .Z(n9349) );
  XNOR U9715 ( .A(n9327), .B(n9352), .Z(n8902) );
  XNOR U9716 ( .A(n9353), .B(n9354), .Z(n9352) );
  NANDN U9717 ( .A(n9325), .B(n9355), .Z(n9354) );
  XOR U9718 ( .A(n9356), .B(n9353), .Z(n9327) );
  OR U9719 ( .A(n9339), .B(n9357), .Z(n9353) );
  XNOR U9720 ( .A(n9342), .B(n9325), .Z(n9339) );
  XNOR U9721 ( .A(n9335), .B(n8912), .Z(n9325) );
  XOR U9722 ( .A(n9358), .B(n9359), .Z(n8912) );
  NANDN U9723 ( .A(n9360), .B(n9361), .Z(n9359) );
  XOR U9724 ( .A(n9362), .B(n9363), .Z(n9335) );
  NANDN U9725 ( .A(n9360), .B(n9364), .Z(n9363) );
  NOR U9726 ( .A(n9342), .B(n9365), .Z(n9356) );
  XOR U9727 ( .A(n9037), .B(n8907), .Z(n9342) );
  XNOR U9728 ( .A(n9366), .B(n9362), .Z(n8907) );
  NANDN U9729 ( .A(n9367), .B(n9368), .Z(n9362) );
  XOR U9730 ( .A(n9364), .B(n9369), .Z(n9368) );
  ANDN U9731 ( .B(n9369), .A(n9370), .Z(n9366) );
  XOR U9732 ( .A(n9371), .B(n9358), .Z(n9037) );
  NANDN U9733 ( .A(n9367), .B(n9372), .Z(n9358) );
  XOR U9734 ( .A(n9373), .B(n9361), .Z(n9372) );
  XNOR U9735 ( .A(n9374), .B(n9375), .Z(n9360) );
  XOR U9736 ( .A(n9376), .B(n9377), .Z(n9375) );
  XNOR U9737 ( .A(n9378), .B(n9379), .Z(n9374) );
  XNOR U9738 ( .A(n9380), .B(n9381), .Z(n9379) );
  ANDN U9739 ( .B(n9373), .A(n9377), .Z(n9380) );
  ANDN U9740 ( .B(n9373), .A(n9370), .Z(n9371) );
  XNOR U9741 ( .A(n9376), .B(n9382), .Z(n9370) );
  XOR U9742 ( .A(n9383), .B(n9381), .Z(n9382) );
  NAND U9743 ( .A(n9384), .B(n9385), .Z(n9381) );
  XNOR U9744 ( .A(n9378), .B(n9361), .Z(n9385) );
  IV U9745 ( .A(n9373), .Z(n9378) );
  XNOR U9746 ( .A(n9364), .B(n9377), .Z(n9384) );
  IV U9747 ( .A(n9369), .Z(n9377) );
  XOR U9748 ( .A(n9386), .B(n9387), .Z(n9369) );
  XNOR U9749 ( .A(n9388), .B(n9389), .Z(n9387) );
  XNOR U9750 ( .A(n9390), .B(n9391), .Z(n9386) );
  ANDN U9751 ( .B(n9351), .A(n9392), .Z(n9390) );
  AND U9752 ( .A(n9361), .B(n9364), .Z(n9383) );
  XNOR U9753 ( .A(n9361), .B(n9364), .Z(n9376) );
  XNOR U9754 ( .A(n9393), .B(n9394), .Z(n9364) );
  XNOR U9755 ( .A(n9395), .B(n9389), .Z(n9394) );
  XOR U9756 ( .A(n9396), .B(n9397), .Z(n9393) );
  XNOR U9757 ( .A(n9398), .B(n9391), .Z(n9397) );
  OR U9758 ( .A(n9034), .B(n9350), .Z(n9391) );
  XNOR U9759 ( .A(n9351), .B(n9399), .Z(n9350) );
  XNOR U9760 ( .A(n9392), .B(n8913), .Z(n9034) );
  ANDN U9761 ( .B(n9400), .A(n9331), .Z(n9398) );
  XNOR U9762 ( .A(n9401), .B(n9402), .Z(n9361) );
  XNOR U9763 ( .A(n9389), .B(n9403), .Z(n9402) );
  XOR U9764 ( .A(n9321), .B(n9396), .Z(n9403) );
  XNOR U9765 ( .A(n9351), .B(n9392), .Z(n9389) );
  XOR U9766 ( .A(n8906), .B(n9404), .Z(n9401) );
  XNOR U9767 ( .A(n9405), .B(n9406), .Z(n9404) );
  ANDN U9768 ( .B(n9407), .A(n9347), .Z(n9405) );
  XNOR U9769 ( .A(n9408), .B(n9409), .Z(n9373) );
  XNOR U9770 ( .A(n9395), .B(n9410), .Z(n9409) );
  XNOR U9771 ( .A(n9334), .B(n9388), .Z(n9410) );
  XOR U9772 ( .A(n9396), .B(n9411), .Z(n9388) );
  XNOR U9773 ( .A(n9412), .B(n9413), .Z(n9411) );
  NAND U9774 ( .A(n9355), .B(n9326), .Z(n9413) );
  XNOR U9775 ( .A(n9414), .B(n9412), .Z(n9396) );
  NANDN U9776 ( .A(n9357), .B(n9340), .Z(n9412) );
  XOR U9777 ( .A(n9341), .B(n9326), .Z(n9340) );
  XNOR U9778 ( .A(n9407), .B(n8913), .Z(n9326) );
  XOR U9779 ( .A(n9365), .B(n9355), .Z(n9357) );
  XNOR U9780 ( .A(n9347), .B(n9399), .Z(n9355) );
  ANDN U9781 ( .B(n9341), .A(n9365), .Z(n9414) );
  XOR U9782 ( .A(n8906), .B(n9351), .Z(n9365) );
  XNOR U9783 ( .A(n9415), .B(n9416), .Z(n9351) );
  XNOR U9784 ( .A(n9417), .B(n9418), .Z(n9416) );
  XOR U9785 ( .A(n9399), .B(n9400), .Z(n9395) );
  IV U9786 ( .A(n8913), .Z(n9400) );
  XOR U9787 ( .A(n9419), .B(n9420), .Z(n8913) );
  XNOR U9788 ( .A(n9421), .B(n9418), .Z(n9420) );
  IV U9789 ( .A(n9331), .Z(n9399) );
  XOR U9790 ( .A(n9418), .B(n9422), .Z(n9331) );
  XNOR U9791 ( .A(n9423), .B(n9424), .Z(n9408) );
  XNOR U9792 ( .A(n9425), .B(n9406), .Z(n9424) );
  OR U9793 ( .A(n9337), .B(n9346), .Z(n9406) );
  XNOR U9794 ( .A(n8906), .B(n9347), .Z(n9346) );
  IV U9795 ( .A(n9423), .Z(n9347) );
  XOR U9796 ( .A(n9321), .B(n9407), .Z(n9337) );
  IV U9797 ( .A(n9334), .Z(n9407) );
  XOR U9798 ( .A(n9036), .B(n9426), .Z(n9334) );
  XNOR U9799 ( .A(n9421), .B(n9415), .Z(n9426) );
  XOR U9800 ( .A(n9427), .B(n9428), .Z(n9415) );
  XNOR U9801 ( .A(n9429), .B(n9430), .Z(n9428) );
  XNOR U9802 ( .A(key[834]), .B(n9431), .Z(n9427) );
  IV U9803 ( .A(n9392), .Z(n9036) );
  XOR U9804 ( .A(n9419), .B(n9432), .Z(n9392) );
  XOR U9805 ( .A(n9418), .B(n9433), .Z(n9432) );
  NOR U9806 ( .A(n9321), .B(n8906), .Z(n9425) );
  XOR U9807 ( .A(n9419), .B(n9434), .Z(n9321) );
  XOR U9808 ( .A(n9418), .B(n9435), .Z(n9434) );
  XOR U9809 ( .A(n9436), .B(n9437), .Z(n9418) );
  XOR U9810 ( .A(n9438), .B(n9439), .Z(n9437) );
  XOR U9811 ( .A(n9440), .B(n9441), .Z(n9436) );
  XOR U9812 ( .A(key[838]), .B(n8906), .Z(n9441) );
  IV U9813 ( .A(n9422), .Z(n9419) );
  XOR U9814 ( .A(n9442), .B(n9443), .Z(n9422) );
  XOR U9815 ( .A(n9444), .B(n9445), .Z(n9443) );
  XOR U9816 ( .A(key[837]), .B(n9446), .Z(n9442) );
  XOR U9817 ( .A(n9447), .B(n9448), .Z(n9423) );
  XNOR U9818 ( .A(n9435), .B(n9433), .Z(n9448) );
  XNOR U9819 ( .A(n9449), .B(n9450), .Z(n9433) );
  XOR U9820 ( .A(n9451), .B(n9452), .Z(n9450) );
  XNOR U9821 ( .A(key[839]), .B(n9453), .Z(n9449) );
  XNOR U9822 ( .A(n9454), .B(n9455), .Z(n9435) );
  XOR U9823 ( .A(n9456), .B(n9457), .Z(n9455) );
  XNOR U9824 ( .A(n9458), .B(n9459), .Z(n9454) );
  XNOR U9825 ( .A(key[836]), .B(n9460), .Z(n9459) );
  XNOR U9826 ( .A(n8906), .B(n9417), .Z(n9447) );
  XOR U9827 ( .A(n9461), .B(n9462), .Z(n9417) );
  XNOR U9828 ( .A(n9463), .B(n9464), .Z(n9462) );
  XNOR U9829 ( .A(n9421), .B(n9465), .Z(n9464) );
  XOR U9830 ( .A(n9466), .B(n9467), .Z(n9421) );
  XOR U9831 ( .A(n9468), .B(n9469), .Z(n9467) );
  XNOR U9832 ( .A(key[833]), .B(n9470), .Z(n9466) );
  XNOR U9833 ( .A(n9471), .B(n9472), .Z(n9461) );
  XNOR U9834 ( .A(key[835]), .B(n9473), .Z(n9472) );
  XNOR U9835 ( .A(n9474), .B(n9475), .Z(n8906) );
  XOR U9836 ( .A(n9476), .B(n9477), .Z(n9475) );
  XNOR U9837 ( .A(key[832]), .B(n9478), .Z(n9474) );
  XOR U9838 ( .A(n8829), .B(n9479), .Z(n7358) );
  XNOR U9839 ( .A(n8831), .B(n8832), .Z(n9479) );
  XNOR U9840 ( .A(n9481), .B(n9482), .Z(n9480) );
  OR U9841 ( .A(n8924), .B(n9483), .Z(n9482) );
  XOR U9842 ( .A(n8919), .B(n9484), .Z(n8860) );
  XNOR U9843 ( .A(n9485), .B(n9486), .Z(n9484) );
  NAND U9844 ( .A(n9487), .B(n8992), .Z(n9486) );
  XOR U9845 ( .A(n8988), .B(n9488), .Z(n8831) );
  XOR U9846 ( .A(n8986), .B(n9489), .Z(n9488) );
  NAND U9847 ( .A(n9490), .B(n8929), .Z(n9489) );
  XOR U9848 ( .A(n8864), .B(n8929), .Z(n8931) );
  XOR U9849 ( .A(n8983), .B(n8817), .Z(n8829) );
  XNOR U9850 ( .A(n8919), .B(n9492), .Z(n8817) );
  XNOR U9851 ( .A(n9481), .B(n9493), .Z(n9492) );
  NANDN U9852 ( .A(n9494), .B(n9495), .Z(n9493) );
  OR U9853 ( .A(n9496), .B(n9497), .Z(n9481) );
  XNOR U9854 ( .A(n9498), .B(n9485), .Z(n8919) );
  NANDN U9855 ( .A(n9499), .B(n9500), .Z(n9485) );
  ANDN U9856 ( .B(n9501), .A(n9502), .Z(n9498) );
  IV U9857 ( .A(n8982), .Z(n8983) );
  XNOR U9858 ( .A(n8988), .B(n9503), .Z(n8982) );
  XOR U9859 ( .A(n9504), .B(n8922), .Z(n9503) );
  OR U9860 ( .A(n9505), .B(n9496), .Z(n8922) );
  XNOR U9861 ( .A(n8924), .B(n9494), .Z(n9496) );
  NOR U9862 ( .A(n9506), .B(n9494), .Z(n9504) );
  XOR U9863 ( .A(n9507), .B(n8990), .Z(n8988) );
  OR U9864 ( .A(n9499), .B(n9508), .Z(n8990) );
  XNOR U9865 ( .A(n9509), .B(n8992), .Z(n9499) );
  XNOR U9866 ( .A(n9494), .B(n8929), .Z(n8992) );
  XOR U9867 ( .A(n9510), .B(n9511), .Z(n8929) );
  NANDN U9868 ( .A(n9512), .B(n9513), .Z(n9511) );
  XNOR U9869 ( .A(n9514), .B(n9515), .Z(n9494) );
  OR U9870 ( .A(n9512), .B(n9516), .Z(n9515) );
  ANDN U9871 ( .B(n9509), .A(n9517), .Z(n9507) );
  IV U9872 ( .A(n9502), .Z(n9509) );
  XOR U9873 ( .A(n8924), .B(n8864), .Z(n9502) );
  XNOR U9874 ( .A(n9518), .B(n9510), .Z(n8864) );
  NANDN U9875 ( .A(n9519), .B(n9520), .Z(n9510) );
  ANDN U9876 ( .B(n9521), .A(n9522), .Z(n9518) );
  NANDN U9877 ( .A(n9519), .B(n9524), .Z(n9514) );
  XOR U9878 ( .A(n9525), .B(n9512), .Z(n9519) );
  XNOR U9879 ( .A(n9526), .B(n9527), .Z(n9512) );
  XOR U9880 ( .A(n9528), .B(n9521), .Z(n9527) );
  XNOR U9881 ( .A(n9529), .B(n9530), .Z(n9526) );
  XNOR U9882 ( .A(n9531), .B(n9532), .Z(n9530) );
  ANDN U9883 ( .B(n9521), .A(n9533), .Z(n9531) );
  IV U9884 ( .A(n9534), .Z(n9521) );
  ANDN U9885 ( .B(n9525), .A(n9533), .Z(n9523) );
  IV U9886 ( .A(n9529), .Z(n9533) );
  IV U9887 ( .A(n9522), .Z(n9525) );
  XNOR U9888 ( .A(n9528), .B(n9535), .Z(n9522) );
  XOR U9889 ( .A(n9536), .B(n9532), .Z(n9535) );
  NAND U9890 ( .A(n9524), .B(n9520), .Z(n9532) );
  XNOR U9891 ( .A(n9513), .B(n9534), .Z(n9520) );
  XOR U9892 ( .A(n9537), .B(n9538), .Z(n9534) );
  XOR U9893 ( .A(n9539), .B(n9540), .Z(n9538) );
  XNOR U9894 ( .A(n9495), .B(n9541), .Z(n9540) );
  XNOR U9895 ( .A(n9542), .B(n9543), .Z(n9537) );
  XNOR U9896 ( .A(n9544), .B(n9545), .Z(n9543) );
  ANDN U9897 ( .B(n9546), .A(n8925), .Z(n9544) );
  XNOR U9898 ( .A(n9529), .B(n9516), .Z(n9524) );
  XOR U9899 ( .A(n9547), .B(n9548), .Z(n9529) );
  XNOR U9900 ( .A(n9549), .B(n9541), .Z(n9548) );
  XOR U9901 ( .A(n9550), .B(n9551), .Z(n9541) );
  XNOR U9902 ( .A(n9552), .B(n9553), .Z(n9551) );
  NAND U9903 ( .A(n8993), .B(n9487), .Z(n9553) );
  XNOR U9904 ( .A(n9554), .B(n9555), .Z(n9547) );
  ANDN U9905 ( .B(n9556), .A(n8987), .Z(n9554) );
  ANDN U9906 ( .B(n9513), .A(n9516), .Z(n9536) );
  XOR U9907 ( .A(n9516), .B(n9513), .Z(n9528) );
  XNOR U9908 ( .A(n9557), .B(n9558), .Z(n9513) );
  XNOR U9909 ( .A(n9550), .B(n9559), .Z(n9558) );
  XOR U9910 ( .A(n9549), .B(n9483), .Z(n9559) );
  XOR U9911 ( .A(n8925), .B(n9560), .Z(n9557) );
  XNOR U9912 ( .A(n9561), .B(n9545), .Z(n9560) );
  OR U9913 ( .A(n9497), .B(n9505), .Z(n9545) );
  XNOR U9914 ( .A(n8925), .B(n9506), .Z(n9505) );
  XOR U9915 ( .A(n9483), .B(n9495), .Z(n9497) );
  ANDN U9916 ( .B(n9495), .A(n9506), .Z(n9561) );
  XOR U9917 ( .A(n9562), .B(n9563), .Z(n9516) );
  XOR U9918 ( .A(n9550), .B(n9539), .Z(n9563) );
  XOR U9919 ( .A(n9490), .B(n8930), .Z(n9539) );
  XOR U9920 ( .A(n9564), .B(n9552), .Z(n9550) );
  NANDN U9921 ( .A(n9508), .B(n9500), .Z(n9552) );
  XOR U9922 ( .A(n9501), .B(n9487), .Z(n9500) );
  XNOR U9923 ( .A(n9556), .B(n9565), .Z(n9495) );
  XNOR U9924 ( .A(n9566), .B(n9567), .Z(n9565) );
  XOR U9925 ( .A(n9517), .B(n8993), .Z(n9508) );
  XNOR U9926 ( .A(n9506), .B(n9490), .Z(n8993) );
  IV U9927 ( .A(n9542), .Z(n9506) );
  XOR U9928 ( .A(n9568), .B(n9569), .Z(n9542) );
  XOR U9929 ( .A(n9570), .B(n9571), .Z(n9569) );
  XNOR U9930 ( .A(n8925), .B(n9572), .Z(n9568) );
  ANDN U9931 ( .B(n9501), .A(n9517), .Z(n9564) );
  XNOR U9932 ( .A(n8925), .B(n8987), .Z(n9517) );
  XOR U9933 ( .A(n9556), .B(n9546), .Z(n9501) );
  IV U9934 ( .A(n9483), .Z(n9546) );
  XOR U9935 ( .A(n9573), .B(n9574), .Z(n9483) );
  XOR U9936 ( .A(n9575), .B(n9571), .Z(n9574) );
  XNOR U9937 ( .A(n9576), .B(n9577), .Z(n9571) );
  XNOR U9938 ( .A(n9578), .B(n9579), .Z(n9577) );
  XOR U9939 ( .A(n9580), .B(n9581), .Z(n9576) );
  XNOR U9940 ( .A(key[876]), .B(n9582), .Z(n9581) );
  IV U9941 ( .A(n8865), .Z(n9556) );
  XOR U9942 ( .A(n9549), .B(n9583), .Z(n9562) );
  XNOR U9943 ( .A(n9584), .B(n9555), .Z(n9583) );
  OR U9944 ( .A(n8932), .B(n9491), .Z(n9555) );
  XNOR U9945 ( .A(n9585), .B(n9490), .Z(n9491) );
  XNOR U9946 ( .A(n8865), .B(n8930), .Z(n8932) );
  ANDN U9947 ( .B(n9490), .A(n8930), .Z(n9584) );
  XOR U9948 ( .A(n9573), .B(n9586), .Z(n8930) );
  XOR U9949 ( .A(n9566), .B(n9587), .Z(n9586) );
  XOR U9950 ( .A(n9575), .B(n9573), .Z(n9490) );
  XNOR U9951 ( .A(n8987), .B(n8865), .Z(n9549) );
  XOR U9952 ( .A(n9573), .B(n9588), .Z(n8865) );
  XNOR U9953 ( .A(n9575), .B(n9570), .Z(n9588) );
  XOR U9954 ( .A(n9589), .B(n9590), .Z(n9570) );
  XNOR U9955 ( .A(n9591), .B(n9592), .Z(n9590) );
  XOR U9956 ( .A(key[879]), .B(n9593), .Z(n9589) );
  XNOR U9957 ( .A(n9594), .B(n9595), .Z(n9573) );
  XNOR U9958 ( .A(n9596), .B(n9597), .Z(n9595) );
  XOR U9959 ( .A(n9598), .B(n9599), .Z(n9594) );
  XNOR U9960 ( .A(key[877]), .B(n9600), .Z(n9599) );
  IV U9961 ( .A(n9585), .Z(n8987) );
  XNOR U9962 ( .A(n9567), .B(n9601), .Z(n9585) );
  XOR U9963 ( .A(n9572), .B(n9587), .Z(n9601) );
  IV U9964 ( .A(n9575), .Z(n9587) );
  XOR U9965 ( .A(n9602), .B(n9603), .Z(n9575) );
  XNOR U9966 ( .A(n9604), .B(n9605), .Z(n9603) );
  XNOR U9967 ( .A(n9606), .B(n9607), .Z(n9602) );
  XOR U9968 ( .A(key[878]), .B(n8925), .Z(n9607) );
  XNOR U9969 ( .A(n9608), .B(n9609), .Z(n8925) );
  XOR U9970 ( .A(n9610), .B(n9611), .Z(n9609) );
  XOR U9971 ( .A(n9612), .B(n9613), .Z(n9608) );
  XNOR U9972 ( .A(key[872]), .B(n9614), .Z(n9613) );
  XOR U9973 ( .A(n9615), .B(n9616), .Z(n9572) );
  XNOR U9974 ( .A(n9617), .B(n9618), .Z(n9616) );
  XOR U9975 ( .A(n9566), .B(n9619), .Z(n9618) );
  XOR U9976 ( .A(n9620), .B(n9621), .Z(n9566) );
  XOR U9977 ( .A(n9622), .B(n9623), .Z(n9621) );
  XOR U9978 ( .A(n9624), .B(n9625), .Z(n9620) );
  XNOR U9979 ( .A(key[873]), .B(n9626), .Z(n9625) );
  XNOR U9980 ( .A(n9627), .B(n9628), .Z(n9615) );
  XNOR U9981 ( .A(key[875]), .B(n9629), .Z(n9628) );
  XOR U9982 ( .A(n9630), .B(n9631), .Z(n9567) );
  XOR U9983 ( .A(n9632), .B(n9633), .Z(n9631) );
  XOR U9984 ( .A(n9634), .B(n9635), .Z(n9630) );
  XOR U9985 ( .A(key[874]), .B(n9636), .Z(n9635) );
  XNOR U9986 ( .A(n8660), .B(n8661), .Z(n2992) );
  XNOR U9987 ( .A(n8702), .B(n9637), .Z(n8661) );
  XOR U9988 ( .A(n9638), .B(n8598), .Z(n9637) );
  OR U9989 ( .A(n9639), .B(n9640), .Z(n8598) );
  ANDN U9990 ( .B(n9641), .A(n9642), .Z(n9638) );
  XNOR U9991 ( .A(n8579), .B(n8495), .Z(n3012) );
  XNOR U9992 ( .A(n8573), .B(n9643), .Z(n8495) );
  XNOR U9993 ( .A(n8570), .B(n9644), .Z(n9643) );
  NANDN U9994 ( .A(n9645), .B(n8527), .Z(n9644) );
  XNOR U9995 ( .A(n8572), .B(n8527), .Z(n8675) );
  XNOR U9996 ( .A(n8573), .B(n9647), .Z(n8579) );
  XOR U9997 ( .A(n9648), .B(n8519), .Z(n9647) );
  OR U9998 ( .A(n8690), .B(n9649), .Z(n8519) );
  XNOR U9999 ( .A(n8522), .B(n8689), .Z(n8690) );
  ANDN U10000 ( .B(n8689), .A(n9650), .Z(n9648) );
  XOR U10001 ( .A(n9651), .B(n8575), .Z(n8573) );
  OR U10002 ( .A(n8693), .B(n9652), .Z(n8575) );
  XOR U10003 ( .A(n8696), .B(n8577), .Z(n8693) );
  XOR U10004 ( .A(n8689), .B(n8527), .Z(n8577) );
  XOR U10005 ( .A(n9653), .B(n9654), .Z(n8527) );
  NANDN U10006 ( .A(n9655), .B(n9656), .Z(n9654) );
  XOR U10007 ( .A(n9657), .B(n9658), .Z(n8689) );
  NANDN U10008 ( .A(n9655), .B(n9659), .Z(n9658) );
  NOR U10009 ( .A(n8696), .B(n9660), .Z(n9651) );
  XOR U10010 ( .A(n8572), .B(n8522), .Z(n8696) );
  XNOR U10011 ( .A(n9661), .B(n9657), .Z(n8522) );
  NANDN U10012 ( .A(n9662), .B(n9663), .Z(n9657) );
  XOR U10013 ( .A(n9659), .B(n9664), .Z(n9663) );
  ANDN U10014 ( .B(n9664), .A(n9665), .Z(n9661) );
  XOR U10015 ( .A(n9666), .B(n9653), .Z(n8572) );
  NANDN U10016 ( .A(n9662), .B(n9667), .Z(n9653) );
  XOR U10017 ( .A(n9668), .B(n9656), .Z(n9667) );
  XNOR U10018 ( .A(n9669), .B(n9670), .Z(n9655) );
  XOR U10019 ( .A(n9671), .B(n9672), .Z(n9670) );
  XNOR U10020 ( .A(n9673), .B(n9674), .Z(n9669) );
  XNOR U10021 ( .A(n9675), .B(n9676), .Z(n9674) );
  ANDN U10022 ( .B(n9668), .A(n9672), .Z(n9675) );
  ANDN U10023 ( .B(n9668), .A(n9665), .Z(n9666) );
  XNOR U10024 ( .A(n9671), .B(n9677), .Z(n9665) );
  XOR U10025 ( .A(n9678), .B(n9676), .Z(n9677) );
  NAND U10026 ( .A(n9679), .B(n9680), .Z(n9676) );
  XNOR U10027 ( .A(n9673), .B(n9656), .Z(n9680) );
  IV U10028 ( .A(n9668), .Z(n9673) );
  XNOR U10029 ( .A(n9659), .B(n9672), .Z(n9679) );
  IV U10030 ( .A(n9664), .Z(n9672) );
  XOR U10031 ( .A(n9681), .B(n9682), .Z(n9664) );
  XNOR U10032 ( .A(n9683), .B(n9684), .Z(n9682) );
  XNOR U10033 ( .A(n9685), .B(n9686), .Z(n9681) );
  ANDN U10034 ( .B(n8571), .A(n8677), .Z(n9685) );
  AND U10035 ( .A(n9656), .B(n9659), .Z(n9678) );
  XNOR U10036 ( .A(n9656), .B(n9659), .Z(n9671) );
  XNOR U10037 ( .A(n9687), .B(n9688), .Z(n9659) );
  XNOR U10038 ( .A(n9689), .B(n9684), .Z(n9688) );
  XOR U10039 ( .A(n9690), .B(n9691), .Z(n9687) );
  XNOR U10040 ( .A(n9692), .B(n9686), .Z(n9691) );
  OR U10041 ( .A(n8676), .B(n9646), .Z(n9686) );
  XNOR U10042 ( .A(n8571), .B(n9693), .Z(n9646) );
  XNOR U10043 ( .A(n8677), .B(n8528), .Z(n8676) );
  ANDN U10044 ( .B(n9694), .A(n9645), .Z(n9692) );
  XNOR U10045 ( .A(n9695), .B(n9696), .Z(n9656) );
  XNOR U10046 ( .A(n9684), .B(n9697), .Z(n9696) );
  XOR U10047 ( .A(n8681), .B(n9690), .Z(n9697) );
  XNOR U10048 ( .A(n8571), .B(n8677), .Z(n9684) );
  XOR U10049 ( .A(n8521), .B(n9698), .Z(n9695) );
  XNOR U10050 ( .A(n9699), .B(n9700), .Z(n9698) );
  ANDN U10051 ( .B(n9701), .A(n9650), .Z(n9699) );
  XNOR U10052 ( .A(n9702), .B(n9703), .Z(n9668) );
  XNOR U10053 ( .A(n9689), .B(n9704), .Z(n9703) );
  XNOR U10054 ( .A(n8688), .B(n9683), .Z(n9704) );
  XOR U10055 ( .A(n9690), .B(n9705), .Z(n9683) );
  XNOR U10056 ( .A(n9706), .B(n9707), .Z(n9705) );
  NAND U10057 ( .A(n8578), .B(n8685), .Z(n9707) );
  XNOR U10058 ( .A(n9708), .B(n9706), .Z(n9690) );
  NANDN U10059 ( .A(n9652), .B(n8694), .Z(n9706) );
  XOR U10060 ( .A(n8695), .B(n8685), .Z(n8694) );
  XNOR U10061 ( .A(n9701), .B(n8528), .Z(n8685) );
  XOR U10062 ( .A(n9660), .B(n8578), .Z(n9652) );
  XNOR U10063 ( .A(n9650), .B(n9693), .Z(n8578) );
  ANDN U10064 ( .B(n8695), .A(n9660), .Z(n9708) );
  XOR U10065 ( .A(n8521), .B(n8571), .Z(n9660) );
  XNOR U10066 ( .A(n9709), .B(n9710), .Z(n8571) );
  XNOR U10067 ( .A(n9711), .B(n9712), .Z(n9710) );
  XOR U10068 ( .A(n9693), .B(n9694), .Z(n9689) );
  IV U10069 ( .A(n8528), .Z(n9694) );
  XOR U10070 ( .A(n9713), .B(n9714), .Z(n8528) );
  XNOR U10071 ( .A(n9715), .B(n9712), .Z(n9714) );
  IV U10072 ( .A(n9645), .Z(n9693) );
  XOR U10073 ( .A(n9712), .B(n9716), .Z(n9645) );
  XNOR U10074 ( .A(n9717), .B(n9718), .Z(n9702) );
  XNOR U10075 ( .A(n9719), .B(n9700), .Z(n9718) );
  OR U10076 ( .A(n8691), .B(n9649), .Z(n9700) );
  XNOR U10077 ( .A(n8521), .B(n9650), .Z(n9649) );
  IV U10078 ( .A(n9717), .Z(n9650) );
  XOR U10079 ( .A(n8681), .B(n9701), .Z(n8691) );
  IV U10080 ( .A(n8688), .Z(n9701) );
  XNOR U10081 ( .A(n9715), .B(n9709), .Z(n9720) );
  XOR U10082 ( .A(n9721), .B(n9722), .Z(n9709) );
  XOR U10083 ( .A(n8250), .B(n9723), .Z(n9722) );
  XNOR U10084 ( .A(n7042), .B(n9724), .Z(n9721) );
  XNOR U10085 ( .A(key[1018]), .B(n6142), .Z(n9724) );
  IV U10086 ( .A(n7046), .Z(n6142) );
  XOR U10087 ( .A(n8251), .B(n8259), .Z(n7046) );
  XOR U10088 ( .A(n9725), .B(n9726), .Z(n7042) );
  XOR U10089 ( .A(n9727), .B(n9728), .Z(n9726) );
  XOR U10090 ( .A(n9713), .B(n9729), .Z(n8677) );
  XOR U10091 ( .A(n9712), .B(n9730), .Z(n9729) );
  NOR U10092 ( .A(n8681), .B(n8521), .Z(n9719) );
  XOR U10093 ( .A(n9713), .B(n9731), .Z(n8681) );
  XOR U10094 ( .A(n9712), .B(n9732), .Z(n9731) );
  XOR U10095 ( .A(n9733), .B(n9734), .Z(n9712) );
  XOR U10096 ( .A(n8521), .B(n6115), .Z(n9734) );
  XOR U10097 ( .A(n9735), .B(n9736), .Z(n6115) );
  XNOR U10098 ( .A(n8230), .B(n9737), .Z(n9733) );
  XNOR U10099 ( .A(key[1022]), .B(n7063), .Z(n9737) );
  XOR U10100 ( .A(n6122), .B(n7058), .Z(n7063) );
  XNOR U10101 ( .A(n9725), .B(n9738), .Z(n8225) );
  XOR U10102 ( .A(n9739), .B(n9740), .Z(n9738) );
  XOR U10103 ( .A(n9741), .B(n9742), .Z(n9725) );
  XOR U10104 ( .A(n8243), .B(n8233), .Z(n6122) );
  IV U10105 ( .A(n6117), .Z(n8233) );
  XOR U10106 ( .A(n9743), .B(n9744), .Z(n6117) );
  XOR U10107 ( .A(n9745), .B(n9746), .Z(n8230) );
  IV U10108 ( .A(n9716), .Z(n9713) );
  XOR U10109 ( .A(n9747), .B(n9748), .Z(n9716) );
  XNOR U10110 ( .A(n8217), .B(n7073), .Z(n9748) );
  XNOR U10111 ( .A(n8231), .B(n6120), .Z(n7073) );
  XNOR U10112 ( .A(n9749), .B(n9750), .Z(n6120) );
  XNOR U10113 ( .A(n9751), .B(n9752), .Z(n9750) );
  XNOR U10114 ( .A(n9753), .B(n9754), .Z(n9749) );
  XOR U10115 ( .A(n9755), .B(n9756), .Z(n9754) );
  ANDN U10116 ( .B(n9757), .A(n9758), .Z(n9756) );
  XNOR U10117 ( .A(n9759), .B(n9760), .Z(n8217) );
  XOR U10118 ( .A(n9761), .B(n9762), .Z(n9760) );
  XNOR U10119 ( .A(n9763), .B(n9764), .Z(n9759) );
  XOR U10120 ( .A(n9765), .B(n9766), .Z(n9764) );
  ANDN U10121 ( .B(n9767), .A(n9768), .Z(n9766) );
  XNOR U10122 ( .A(n8243), .B(n9769), .Z(n9747) );
  XNOR U10123 ( .A(key[1021]), .B(n7065), .Z(n9769) );
  XOR U10124 ( .A(n9739), .B(n9728), .Z(n7065) );
  XNOR U10125 ( .A(n9770), .B(n9771), .Z(n9728) );
  XNOR U10126 ( .A(n9772), .B(n9773), .Z(n9771) );
  ANDN U10127 ( .B(n9774), .A(n9775), .Z(n9772) );
  XNOR U10128 ( .A(n9776), .B(n9777), .Z(n8243) );
  XOR U10129 ( .A(n9778), .B(n9779), .Z(n9717) );
  XNOR U10130 ( .A(n9732), .B(n9730), .Z(n9779) );
  XNOR U10131 ( .A(n9780), .B(n9781), .Z(n9730) );
  XNOR U10132 ( .A(n8226), .B(n7059), .Z(n9781) );
  XNOR U10133 ( .A(n9736), .B(n8241), .Z(n7059) );
  XNOR U10134 ( .A(n9782), .B(n9783), .Z(n8241) );
  XOR U10135 ( .A(n9743), .B(n9752), .Z(n9783) );
  XNOR U10136 ( .A(n9784), .B(n9785), .Z(n9752) );
  XNOR U10137 ( .A(n9786), .B(n9787), .Z(n9785) );
  NANDN U10138 ( .A(n9788), .B(n9789), .Z(n9787) );
  XOR U10139 ( .A(n9790), .B(n9791), .Z(n9782) );
  IV U10140 ( .A(n8227), .Z(n9736) );
  XNOR U10141 ( .A(n9792), .B(n9793), .Z(n8227) );
  XNOR U10142 ( .A(n9776), .B(n9794), .Z(n9793) );
  XNOR U10143 ( .A(n9795), .B(n9796), .Z(n9792) );
  XNOR U10144 ( .A(n9797), .B(n9798), .Z(n8226) );
  XNOR U10145 ( .A(n9799), .B(n9762), .Z(n9798) );
  XNOR U10146 ( .A(n9800), .B(n9801), .Z(n9762) );
  XNOR U10147 ( .A(n9802), .B(n9803), .Z(n9801) );
  NANDN U10148 ( .A(n9804), .B(n9805), .Z(n9803) );
  XOR U10149 ( .A(n9806), .B(n9745), .Z(n9797) );
  XNOR U10150 ( .A(key[1023]), .B(n7069), .Z(n9780) );
  XNOR U10151 ( .A(n6129), .B(n6152), .Z(n7069) );
  XNOR U10152 ( .A(n9807), .B(n9808), .Z(n9732) );
  XNOR U10153 ( .A(n7050), .B(n6132), .Z(n9808) );
  XOR U10154 ( .A(n9735), .B(n8231), .Z(n6132) );
  XOR U10155 ( .A(n9809), .B(n9810), .Z(n8231) );
  XNOR U10156 ( .A(n9811), .B(n9794), .Z(n9810) );
  XNOR U10157 ( .A(n9812), .B(n9813), .Z(n9794) );
  XNOR U10158 ( .A(n9814), .B(n9815), .Z(n9813) );
  NANDN U10159 ( .A(n9816), .B(n9817), .Z(n9815) );
  XNOR U10160 ( .A(n9818), .B(n9819), .Z(n9809) );
  XNOR U10161 ( .A(n9820), .B(n9821), .Z(n9819) );
  ANDN U10162 ( .B(n9822), .A(n9823), .Z(n9821) );
  XOR U10163 ( .A(n9753), .B(n8251), .Z(n6134) );
  IV U10164 ( .A(n6107), .Z(n8251) );
  XNOR U10165 ( .A(n9824), .B(n9790), .Z(n6107) );
  XNOR U10166 ( .A(n7052), .B(n9825), .Z(n9807) );
  XNOR U10167 ( .A(key[1020]), .B(n8212), .Z(n9825) );
  XOR U10168 ( .A(n8250), .B(n9761), .Z(n8212) );
  XOR U10169 ( .A(n9826), .B(n9827), .Z(n8250) );
  XOR U10170 ( .A(n6152), .B(n7075), .Z(n7052) );
  XNOR U10171 ( .A(n9828), .B(n9829), .Z(n7075) );
  XOR U10172 ( .A(n9830), .B(n9740), .Z(n9829) );
  XNOR U10173 ( .A(n9831), .B(n9832), .Z(n9740) );
  XNOR U10174 ( .A(n9833), .B(n9834), .Z(n9832) );
  OR U10175 ( .A(n9835), .B(n9836), .Z(n9834) );
  XNOR U10176 ( .A(n9837), .B(n9838), .Z(n9828) );
  XOR U10177 ( .A(n9773), .B(n9839), .Z(n9838) );
  ANDN U10178 ( .B(n9840), .A(n9841), .Z(n9839) );
  ANDN U10179 ( .B(n9842), .A(n9843), .Z(n9773) );
  XNOR U10180 ( .A(n8521), .B(n9711), .Z(n9778) );
  XOR U10181 ( .A(n9844), .B(n9845), .Z(n9711) );
  XNOR U10182 ( .A(n9715), .B(n9846), .Z(n9845) );
  XOR U10183 ( .A(n9735), .B(n8215), .Z(n6139) );
  XOR U10184 ( .A(n9818), .B(n8259), .Z(n8215) );
  XOR U10185 ( .A(n9723), .B(n6145), .Z(n6106) );
  XNOR U10186 ( .A(n9847), .B(n9848), .Z(n6145) );
  XNOR U10187 ( .A(n9849), .B(n9744), .Z(n9848) );
  XNOR U10188 ( .A(n9850), .B(n9851), .Z(n9744) );
  XNOR U10189 ( .A(n9852), .B(n9755), .Z(n9851) );
  ANDN U10190 ( .B(n9853), .A(n9854), .Z(n9755) );
  ANDN U10191 ( .B(n9855), .A(n9856), .Z(n9852) );
  XNOR U10192 ( .A(n9790), .B(n9857), .Z(n9847) );
  IV U10193 ( .A(n8253), .Z(n9723) );
  XOR U10194 ( .A(n9858), .B(n9859), .Z(n8253) );
  XNOR U10195 ( .A(n9860), .B(n9777), .Z(n9859) );
  XNOR U10196 ( .A(n9861), .B(n9862), .Z(n9777) );
  XOR U10197 ( .A(n9863), .B(n9820), .Z(n9862) );
  NANDN U10198 ( .A(n9864), .B(n9865), .Z(n9820) );
  ANDN U10199 ( .B(n9866), .A(n9867), .Z(n9863) );
  XOR U10200 ( .A(n9795), .B(n9868), .Z(n9858) );
  XOR U10201 ( .A(n9869), .B(n9870), .Z(n9715) );
  XNOR U10202 ( .A(n7045), .B(n6150), .Z(n9870) );
  XNOR U10203 ( .A(n8249), .B(n6143), .Z(n6150) );
  XNOR U10204 ( .A(n9743), .B(n9871), .Z(n6143) );
  XOR U10205 ( .A(n9790), .B(n9857), .Z(n9871) );
  IV U10206 ( .A(n9791), .Z(n9857) );
  XOR U10207 ( .A(n9850), .B(n9872), .Z(n9791) );
  XNOR U10208 ( .A(n9873), .B(n9874), .Z(n9872) );
  NANDN U10209 ( .A(n9875), .B(n9789), .Z(n9874) );
  XNOR U10210 ( .A(n9751), .B(n9876), .Z(n9850) );
  XNOR U10211 ( .A(n9877), .B(n9878), .Z(n9876) );
  NANDN U10212 ( .A(n9879), .B(n9880), .Z(n9878) );
  XOR U10213 ( .A(n9881), .B(n9882), .Z(n9790) );
  XNOR U10214 ( .A(n9883), .B(n9884), .Z(n9882) );
  NANDN U10215 ( .A(n9885), .B(n9757), .Z(n9884) );
  XNOR U10216 ( .A(n9824), .B(n9849), .Z(n9743) );
  XNOR U10217 ( .A(n9751), .B(n9886), .Z(n9849) );
  XNOR U10218 ( .A(n9873), .B(n9887), .Z(n9886) );
  NANDN U10219 ( .A(n9888), .B(n9889), .Z(n9887) );
  OR U10220 ( .A(n9890), .B(n9891), .Z(n9873) );
  XOR U10221 ( .A(n9892), .B(n9877), .Z(n9751) );
  NANDN U10222 ( .A(n9893), .B(n9894), .Z(n9877) );
  ANDN U10223 ( .B(n9895), .A(n9896), .Z(n9892) );
  XOR U10224 ( .A(n8259), .B(n9897), .Z(n9869) );
  XNOR U10225 ( .A(key[1017]), .B(n8239), .Z(n9897) );
  XOR U10226 ( .A(n9827), .B(n9898), .Z(n8239) );
  XNOR U10227 ( .A(n9806), .B(n9745), .Z(n9898) );
  XOR U10228 ( .A(n9899), .B(n9900), .Z(n9745) );
  XOR U10229 ( .A(n9901), .B(n9795), .Z(n8259) );
  XNOR U10230 ( .A(n7040), .B(n9902), .Z(n9844) );
  XNOR U10231 ( .A(n9903), .B(n9904), .Z(n8255) );
  XNOR U10232 ( .A(n9799), .B(n9746), .Z(n9904) );
  XNOR U10233 ( .A(n9905), .B(n9906), .Z(n9746) );
  XNOR U10234 ( .A(n9907), .B(n9765), .Z(n9906) );
  NOR U10235 ( .A(n9908), .B(n9909), .Z(n9765) );
  ANDN U10236 ( .B(n9910), .A(n9911), .Z(n9907) );
  IV U10237 ( .A(n9827), .Z(n9799) );
  XOR U10238 ( .A(n9912), .B(n9913), .Z(n9827) );
  XOR U10239 ( .A(n9914), .B(n9915), .Z(n9913) );
  NANDN U10240 ( .A(n9916), .B(n9767), .Z(n9915) );
  XOR U10241 ( .A(n9806), .B(n9900), .Z(n9903) );
  XOR U10242 ( .A(n9763), .B(n9917), .Z(n9900) );
  XNOR U10243 ( .A(n9918), .B(n9919), .Z(n9917) );
  NANDN U10244 ( .A(n9920), .B(n9921), .Z(n9919) );
  XNOR U10245 ( .A(n9918), .B(n9923), .Z(n9922) );
  NAND U10246 ( .A(n9924), .B(n9805), .Z(n9923) );
  OR U10247 ( .A(n9925), .B(n9926), .Z(n9918) );
  XNOR U10248 ( .A(n9763), .B(n9927), .Z(n9905) );
  XNOR U10249 ( .A(n9928), .B(n9929), .Z(n9927) );
  OR U10250 ( .A(n9930), .B(n9931), .Z(n9929) );
  XOR U10251 ( .A(n9932), .B(n9928), .Z(n9763) );
  OR U10252 ( .A(n9933), .B(n9934), .Z(n9928) );
  ANDN U10253 ( .B(n9935), .A(n9936), .Z(n9932) );
  XNOR U10254 ( .A(n6152), .B(n7054), .Z(n7040) );
  XOR U10255 ( .A(n9837), .B(n7045), .Z(n7054) );
  XNOR U10256 ( .A(n9937), .B(n9741), .Z(n7045) );
  XNOR U10257 ( .A(n9937), .B(n9837), .Z(n6152) );
  XNOR U10258 ( .A(n9831), .B(n9938), .Z(n9837) );
  XNOR U10259 ( .A(n9939), .B(n9940), .Z(n9938) );
  ANDN U10260 ( .B(n9774), .A(n9941), .Z(n9939) );
  XNOR U10261 ( .A(n9942), .B(n9943), .Z(n9831) );
  XNOR U10262 ( .A(n9944), .B(n9945), .Z(n9943) );
  NAND U10263 ( .A(n9946), .B(n9947), .Z(n9945) );
  XNOR U10264 ( .A(n9948), .B(n9949), .Z(n8521) );
  XOR U10265 ( .A(n8249), .B(n6151), .Z(n9949) );
  XOR U10266 ( .A(n7070), .B(n8216), .Z(n6151) );
  XOR U10267 ( .A(n9899), .B(n9761), .Z(n8216) );
  XOR U10268 ( .A(n9800), .B(n9950), .Z(n9761) );
  XNOR U10269 ( .A(n9951), .B(n9914), .Z(n9950) );
  NOR U10270 ( .A(n9908), .B(n9952), .Z(n9914) );
  XNOR U10271 ( .A(n9910), .B(n9767), .Z(n9908) );
  XNOR U10272 ( .A(n9912), .B(n9954), .Z(n9800) );
  XNOR U10273 ( .A(n9955), .B(n9956), .Z(n9954) );
  NANDN U10274 ( .A(n9930), .B(n9957), .Z(n9956) );
  IV U10275 ( .A(n9826), .Z(n9899) );
  XNOR U10276 ( .A(n9912), .B(n9958), .Z(n9826) );
  XOR U10277 ( .A(n9959), .B(n9802), .Z(n9958) );
  OR U10278 ( .A(n9960), .B(n9925), .Z(n9802) );
  XNOR U10279 ( .A(n9805), .B(n9921), .Z(n9925) );
  ANDN U10280 ( .B(n9921), .A(n9961), .Z(n9959) );
  XOR U10281 ( .A(n9962), .B(n9955), .Z(n9912) );
  OR U10282 ( .A(n9933), .B(n9963), .Z(n9955) );
  XOR U10283 ( .A(n9935), .B(n9930), .Z(n9933) );
  XNOR U10284 ( .A(n9921), .B(n9767), .Z(n9930) );
  XNOR U10285 ( .A(n9964), .B(n9965), .Z(n9767) );
  NANDN U10286 ( .A(n9966), .B(n9967), .Z(n9965) );
  XOR U10287 ( .A(n9968), .B(n9969), .Z(n9921) );
  NANDN U10288 ( .A(n9966), .B(n9970), .Z(n9969) );
  XOR U10289 ( .A(n9910), .B(n9805), .Z(n9935) );
  XNOR U10290 ( .A(n9972), .B(n9968), .Z(n9805) );
  NANDN U10291 ( .A(n9973), .B(n9974), .Z(n9968) );
  XOR U10292 ( .A(n9970), .B(n9975), .Z(n9974) );
  ANDN U10293 ( .B(n9975), .A(n9976), .Z(n9972) );
  XOR U10294 ( .A(n9977), .B(n9964), .Z(n9910) );
  ANDN U10295 ( .B(n9978), .A(n9973), .Z(n9964) );
  XNOR U10296 ( .A(n9979), .B(n9980), .Z(n9966) );
  XOR U10297 ( .A(n9981), .B(n9982), .Z(n9980) );
  XNOR U10298 ( .A(n9983), .B(n9984), .Z(n9979) );
  XNOR U10299 ( .A(n9985), .B(n9986), .Z(n9984) );
  ANDN U10300 ( .B(n9987), .A(n9982), .Z(n9985) );
  XOR U10301 ( .A(n9987), .B(n9967), .Z(n9978) );
  ANDN U10302 ( .B(n9987), .A(n9976), .Z(n9977) );
  XNOR U10303 ( .A(n9981), .B(n9988), .Z(n9976) );
  XOR U10304 ( .A(n9989), .B(n9986), .Z(n9988) );
  NAND U10305 ( .A(n9990), .B(n9991), .Z(n9986) );
  XNOR U10306 ( .A(n9983), .B(n9967), .Z(n9991) );
  IV U10307 ( .A(n9987), .Z(n9983) );
  XNOR U10308 ( .A(n9970), .B(n9982), .Z(n9990) );
  IV U10309 ( .A(n9975), .Z(n9982) );
  XOR U10310 ( .A(n9992), .B(n9993), .Z(n9975) );
  XNOR U10311 ( .A(n9994), .B(n9995), .Z(n9993) );
  XNOR U10312 ( .A(n9996), .B(n9997), .Z(n9992) );
  ANDN U10313 ( .B(n9953), .A(n9911), .Z(n9996) );
  AND U10314 ( .A(n9967), .B(n9970), .Z(n9989) );
  XNOR U10315 ( .A(n9967), .B(n9970), .Z(n9981) );
  XNOR U10316 ( .A(n9998), .B(n9999), .Z(n9970) );
  XNOR U10317 ( .A(n10000), .B(n9995), .Z(n9999) );
  XOR U10318 ( .A(n10001), .B(n10002), .Z(n9998) );
  XNOR U10319 ( .A(n10003), .B(n9997), .Z(n10002) );
  OR U10320 ( .A(n9909), .B(n9952), .Z(n9997) );
  XNOR U10321 ( .A(n9953), .B(n10034), .Z(n9952) );
  XNOR U10322 ( .A(n9911), .B(n9768), .Z(n9909) );
  ANDN U10323 ( .B(n10004), .A(n9916), .Z(n10003) );
  XNOR U10324 ( .A(n10005), .B(n10006), .Z(n9967) );
  XNOR U10325 ( .A(n9995), .B(n10007), .Z(n10006) );
  XNOR U10326 ( .A(n9924), .B(n10001), .Z(n10007) );
  XNOR U10327 ( .A(n9911), .B(n9953), .Z(n9995) );
  XOR U10328 ( .A(n9804), .B(n10008), .Z(n10005) );
  XNOR U10329 ( .A(n10009), .B(n10010), .Z(n10008) );
  ANDN U10330 ( .B(n10011), .A(n9961), .Z(n10009) );
  XNOR U10331 ( .A(n10012), .B(n10013), .Z(n9987) );
  XNOR U10332 ( .A(n10000), .B(n10014), .Z(n10013) );
  XNOR U10333 ( .A(n10015), .B(n9994), .Z(n10014) );
  XOR U10334 ( .A(n10001), .B(n10016), .Z(n9994) );
  XNOR U10335 ( .A(n10017), .B(n10018), .Z(n10016) );
  NANDN U10336 ( .A(n9931), .B(n9957), .Z(n10018) );
  XNOR U10337 ( .A(n10019), .B(n10017), .Z(n10001) );
  OR U10338 ( .A(n9963), .B(n9934), .Z(n10017) );
  XOR U10339 ( .A(n10020), .B(n9931), .Z(n9934) );
  XNOR U10340 ( .A(n10004), .B(n10011), .Z(n9931) );
  IV U10341 ( .A(n9768), .Z(n10004) );
  XNOR U10342 ( .A(n9971), .B(n9957), .Z(n9963) );
  XNOR U10343 ( .A(n9961), .B(n10034), .Z(n9957) );
  ANDN U10344 ( .B(n9971), .A(n9936), .Z(n10019) );
  IV U10345 ( .A(n10020), .Z(n9936) );
  XOR U10346 ( .A(n10021), .B(n9924), .Z(n10020) );
  XOR U10347 ( .A(n9768), .B(n9916), .Z(n10000) );
  XOR U10348 ( .A(n10022), .B(n10023), .Z(n9916) );
  XOR U10349 ( .A(n10024), .B(n10025), .Z(n9768) );
  XOR U10350 ( .A(n10026), .B(n10023), .Z(n10025) );
  XNOR U10351 ( .A(n9920), .B(n10027), .Z(n10012) );
  XNOR U10352 ( .A(n10028), .B(n10010), .Z(n10027) );
  OR U10353 ( .A(n9926), .B(n9960), .Z(n10010) );
  XNOR U10354 ( .A(n9804), .B(n9961), .Z(n9960) );
  IV U10355 ( .A(n10015), .Z(n9961) );
  XOR U10356 ( .A(n10029), .B(n10030), .Z(n10015) );
  XNOR U10357 ( .A(n10031), .B(n10032), .Z(n10030) );
  XNOR U10358 ( .A(n9804), .B(n10033), .Z(n10029) );
  XNOR U10359 ( .A(n9924), .B(n10011), .Z(n9926) );
  IV U10360 ( .A(n9920), .Z(n10011) );
  ANDN U10361 ( .B(n9924), .A(n9804), .Z(n10028) );
  XOR U10362 ( .A(n10031), .B(n10034), .Z(n9924) );
  XOR U10363 ( .A(n10035), .B(n10036), .Z(n10031) );
  XNOR U10364 ( .A(n10037), .B(n10038), .Z(n10035) );
  XNOR U10365 ( .A(key[772]), .B(n10039), .Z(n10038) );
  XNOR U10366 ( .A(n10040), .B(n10041), .Z(n9920) );
  XOR U10367 ( .A(n9911), .B(n10024), .Z(n10041) );
  IV U10368 ( .A(n10021), .Z(n9911) );
  XOR U10369 ( .A(n10033), .B(n10034), .Z(n10021) );
  XNOR U10370 ( .A(n10022), .B(n10023), .Z(n10034) );
  IV U10371 ( .A(n10026), .Z(n10022) );
  XNOR U10372 ( .A(n10042), .B(n10043), .Z(n10026) );
  XOR U10373 ( .A(n10044), .B(n10045), .Z(n10043) );
  XOR U10374 ( .A(key[773]), .B(n10046), .Z(n10042) );
  XOR U10375 ( .A(n10047), .B(n10048), .Z(n10033) );
  XNOR U10376 ( .A(n10049), .B(n10050), .Z(n10048) );
  XNOR U10377 ( .A(key[775]), .B(n10051), .Z(n10047) );
  XNOR U10378 ( .A(n9804), .B(n9953), .Z(n9971) );
  XNOR U10379 ( .A(n10032), .B(n10052), .Z(n9953) );
  XNOR U10380 ( .A(n10023), .B(n10040), .Z(n10052) );
  XOR U10381 ( .A(n10053), .B(n10054), .Z(n10040) );
  XOR U10382 ( .A(n9166), .B(n9159), .Z(n10054) );
  XNOR U10383 ( .A(key[770]), .B(n10055), .Z(n10053) );
  XOR U10384 ( .A(n10056), .B(n10057), .Z(n10023) );
  XOR U10385 ( .A(n9804), .B(n10058), .Z(n10057) );
  XNOR U10386 ( .A(n10059), .B(n10060), .Z(n10056) );
  XOR U10387 ( .A(key[774]), .B(n10061), .Z(n10060) );
  XOR U10388 ( .A(n10062), .B(n10063), .Z(n10032) );
  XNOR U10389 ( .A(n10064), .B(n10065), .Z(n10063) );
  XNOR U10390 ( .A(n10024), .B(n10066), .Z(n10065) );
  XNOR U10391 ( .A(n10067), .B(n10068), .Z(n10024) );
  XOR U10392 ( .A(n10069), .B(n9147), .Z(n10068) );
  XOR U10393 ( .A(n10070), .B(n10071), .Z(n10062) );
  XOR U10394 ( .A(key[771]), .B(n9146), .Z(n10071) );
  XNOR U10395 ( .A(n10072), .B(n10073), .Z(n9804) );
  XNOR U10396 ( .A(n9165), .B(n10074), .Z(n10073) );
  IV U10397 ( .A(n10075), .Z(n9165) );
  XOR U10398 ( .A(key[768]), .B(n10076), .Z(n10072) );
  IV U10399 ( .A(n8213), .Z(n7070) );
  XOR U10400 ( .A(n9753), .B(n9824), .Z(n8213) );
  XOR U10401 ( .A(n9881), .B(n10077), .Z(n9824) );
  XOR U10402 ( .A(n10078), .B(n9786), .Z(n10077) );
  OR U10403 ( .A(n10079), .B(n9890), .Z(n9786) );
  XNOR U10404 ( .A(n9789), .B(n9889), .Z(n9890) );
  ANDN U10405 ( .B(n9889), .A(n10080), .Z(n10078) );
  XNOR U10406 ( .A(n9784), .B(n10081), .Z(n9753) );
  XOR U10407 ( .A(n10082), .B(n9883), .Z(n10081) );
  XOR U10408 ( .A(n10084), .B(n9757), .Z(n9853) );
  ANDN U10409 ( .B(n10085), .A(n9856), .Z(n10082) );
  IV U10410 ( .A(n10084), .Z(n9856) );
  XNOR U10411 ( .A(n9881), .B(n10086), .Z(n9784) );
  XNOR U10412 ( .A(n10087), .B(n10088), .Z(n10086) );
  NANDN U10413 ( .A(n9879), .B(n10089), .Z(n10088) );
  XOR U10414 ( .A(n10090), .B(n10087), .Z(n9881) );
  OR U10415 ( .A(n9893), .B(n10091), .Z(n10087) );
  XNOR U10416 ( .A(n9896), .B(n9879), .Z(n9893) );
  XNOR U10417 ( .A(n9889), .B(n9757), .Z(n9879) );
  XOR U10418 ( .A(n10092), .B(n10093), .Z(n9757) );
  NANDN U10419 ( .A(n10094), .B(n10095), .Z(n10093) );
  XOR U10420 ( .A(n10096), .B(n10097), .Z(n9889) );
  NANDN U10421 ( .A(n10094), .B(n10098), .Z(n10097) );
  NOR U10422 ( .A(n9896), .B(n10099), .Z(n10090) );
  XNOR U10423 ( .A(n10084), .B(n9789), .Z(n9896) );
  XNOR U10424 ( .A(n10100), .B(n10096), .Z(n9789) );
  NANDN U10425 ( .A(n10101), .B(n10102), .Z(n10096) );
  XOR U10426 ( .A(n10098), .B(n10103), .Z(n10102) );
  ANDN U10427 ( .B(n10103), .A(n10104), .Z(n10100) );
  XNOR U10428 ( .A(n10105), .B(n10092), .Z(n10084) );
  NANDN U10429 ( .A(n10101), .B(n10106), .Z(n10092) );
  XOR U10430 ( .A(n10107), .B(n10095), .Z(n10106) );
  XNOR U10431 ( .A(n10108), .B(n10109), .Z(n10094) );
  XOR U10432 ( .A(n10110), .B(n10111), .Z(n10109) );
  XNOR U10433 ( .A(n10112), .B(n10113), .Z(n10108) );
  XNOR U10434 ( .A(n10114), .B(n10115), .Z(n10113) );
  ANDN U10435 ( .B(n10107), .A(n10111), .Z(n10114) );
  ANDN U10436 ( .B(n10107), .A(n10104), .Z(n10105) );
  XNOR U10437 ( .A(n10110), .B(n10116), .Z(n10104) );
  XOR U10438 ( .A(n10117), .B(n10115), .Z(n10116) );
  NAND U10439 ( .A(n10118), .B(n10119), .Z(n10115) );
  XNOR U10440 ( .A(n10112), .B(n10095), .Z(n10119) );
  IV U10441 ( .A(n10107), .Z(n10112) );
  XNOR U10442 ( .A(n10098), .B(n10111), .Z(n10118) );
  IV U10443 ( .A(n10103), .Z(n10111) );
  XOR U10444 ( .A(n10120), .B(n10121), .Z(n10103) );
  XNOR U10445 ( .A(n10122), .B(n10123), .Z(n10121) );
  XNOR U10446 ( .A(n10124), .B(n10125), .Z(n10120) );
  ANDN U10447 ( .B(n10085), .A(n10126), .Z(n10124) );
  AND U10448 ( .A(n10095), .B(n10098), .Z(n10117) );
  XNOR U10449 ( .A(n10095), .B(n10098), .Z(n10110) );
  XNOR U10450 ( .A(n10127), .B(n10128), .Z(n10098) );
  XNOR U10451 ( .A(n10129), .B(n10123), .Z(n10128) );
  XOR U10452 ( .A(n10130), .B(n10131), .Z(n10127) );
  XNOR U10453 ( .A(n10132), .B(n10125), .Z(n10131) );
  OR U10454 ( .A(n9854), .B(n10083), .Z(n10125) );
  XNOR U10455 ( .A(n10085), .B(n10133), .Z(n10083) );
  XNOR U10456 ( .A(n10126), .B(n9758), .Z(n9854) );
  ANDN U10457 ( .B(n10134), .A(n9885), .Z(n10132) );
  XNOR U10458 ( .A(n10135), .B(n10136), .Z(n10095) );
  XNOR U10459 ( .A(n10123), .B(n10137), .Z(n10136) );
  XOR U10460 ( .A(n9875), .B(n10130), .Z(n10137) );
  XNOR U10461 ( .A(n10085), .B(n10126), .Z(n10123) );
  XOR U10462 ( .A(n9788), .B(n10138), .Z(n10135) );
  XNOR U10463 ( .A(n10139), .B(n10140), .Z(n10138) );
  ANDN U10464 ( .B(n10141), .A(n10080), .Z(n10139) );
  XNOR U10465 ( .A(n10142), .B(n10143), .Z(n10107) );
  XNOR U10466 ( .A(n10129), .B(n10144), .Z(n10143) );
  XNOR U10467 ( .A(n9888), .B(n10122), .Z(n10144) );
  XOR U10468 ( .A(n10130), .B(n10145), .Z(n10122) );
  XNOR U10469 ( .A(n10146), .B(n10147), .Z(n10145) );
  NAND U10470 ( .A(n10089), .B(n9880), .Z(n10147) );
  XNOR U10471 ( .A(n10148), .B(n10146), .Z(n10130) );
  NANDN U10472 ( .A(n10091), .B(n9894), .Z(n10146) );
  XOR U10473 ( .A(n9895), .B(n9880), .Z(n9894) );
  XNOR U10474 ( .A(n10141), .B(n9758), .Z(n9880) );
  XOR U10475 ( .A(n10099), .B(n10089), .Z(n10091) );
  XNOR U10476 ( .A(n10080), .B(n10133), .Z(n10089) );
  ANDN U10477 ( .B(n9895), .A(n10099), .Z(n10148) );
  XOR U10478 ( .A(n9788), .B(n10085), .Z(n10099) );
  XNOR U10479 ( .A(n10149), .B(n10150), .Z(n10085) );
  XNOR U10480 ( .A(n10151), .B(n10152), .Z(n10150) );
  XOR U10481 ( .A(n10133), .B(n10134), .Z(n10129) );
  IV U10482 ( .A(n9758), .Z(n10134) );
  XOR U10483 ( .A(n10153), .B(n10154), .Z(n9758) );
  XOR U10484 ( .A(n10155), .B(n10152), .Z(n10154) );
  IV U10485 ( .A(n9885), .Z(n10133) );
  XOR U10486 ( .A(n10152), .B(n10156), .Z(n9885) );
  XNOR U10487 ( .A(n10157), .B(n10158), .Z(n10142) );
  XNOR U10488 ( .A(n10159), .B(n10140), .Z(n10158) );
  OR U10489 ( .A(n9891), .B(n10079), .Z(n10140) );
  XNOR U10490 ( .A(n9788), .B(n10080), .Z(n10079) );
  IV U10491 ( .A(n10157), .Z(n10080) );
  XOR U10492 ( .A(n9875), .B(n10141), .Z(n9891) );
  IV U10493 ( .A(n9888), .Z(n10141) );
  XOR U10494 ( .A(n9855), .B(n10160), .Z(n9888) );
  XNOR U10495 ( .A(n10161), .B(n10149), .Z(n10160) );
  XOR U10496 ( .A(n10162), .B(n10163), .Z(n10149) );
  XNOR U10497 ( .A(n10164), .B(n10165), .Z(n10163) );
  XNOR U10498 ( .A(n9302), .B(n10166), .Z(n10162) );
  XOR U10499 ( .A(key[810]), .B(n10167), .Z(n10166) );
  IV U10500 ( .A(n10126), .Z(n9855) );
  XOR U10501 ( .A(n10153), .B(n10168), .Z(n10126) );
  XOR U10502 ( .A(n10152), .B(n10169), .Z(n10168) );
  NOR U10503 ( .A(n9875), .B(n9788), .Z(n10159) );
  XOR U10504 ( .A(n10153), .B(n10170), .Z(n9875) );
  XOR U10505 ( .A(n10152), .B(n10171), .Z(n10170) );
  XOR U10506 ( .A(n10172), .B(n10173), .Z(n10152) );
  XOR U10507 ( .A(n10174), .B(n10175), .Z(n10173) );
  XOR U10508 ( .A(n9788), .B(n10176), .Z(n10172) );
  XOR U10509 ( .A(key[814]), .B(n10177), .Z(n10176) );
  IV U10510 ( .A(n10156), .Z(n10153) );
  XOR U10511 ( .A(n10178), .B(n10179), .Z(n10156) );
  XNOR U10512 ( .A(n10180), .B(n10181), .Z(n10179) );
  XOR U10513 ( .A(n10182), .B(n10183), .Z(n10178) );
  XNOR U10514 ( .A(key[813]), .B(n10184), .Z(n10183) );
  XOR U10515 ( .A(n10185), .B(n10186), .Z(n10157) );
  XNOR U10516 ( .A(n10171), .B(n10169), .Z(n10186) );
  XNOR U10517 ( .A(n10187), .B(n10188), .Z(n10169) );
  XNOR U10518 ( .A(n10189), .B(n10190), .Z(n10188) );
  XOR U10519 ( .A(key[815]), .B(n9313), .Z(n10187) );
  IV U10520 ( .A(n10191), .Z(n9313) );
  XNOR U10521 ( .A(n10192), .B(n10193), .Z(n10171) );
  XOR U10522 ( .A(n10194), .B(n10195), .Z(n10193) );
  XNOR U10523 ( .A(n10196), .B(n10197), .Z(n10192) );
  XOR U10524 ( .A(key[812]), .B(n10198), .Z(n10197) );
  XNOR U10525 ( .A(n9788), .B(n10151), .Z(n10185) );
  XOR U10526 ( .A(n10199), .B(n10200), .Z(n10151) );
  XNOR U10527 ( .A(n10201), .B(n10202), .Z(n10200) );
  XOR U10528 ( .A(n10203), .B(n10161), .Z(n10202) );
  IV U10529 ( .A(n10155), .Z(n10161) );
  XNOR U10530 ( .A(n10204), .B(n10205), .Z(n10155) );
  XNOR U10531 ( .A(n10206), .B(n10207), .Z(n10205) );
  XNOR U10532 ( .A(n9259), .B(n10208), .Z(n10204) );
  XOR U10533 ( .A(key[809]), .B(n10209), .Z(n10208) );
  XNOR U10534 ( .A(n10210), .B(n10211), .Z(n10199) );
  XNOR U10535 ( .A(key[811]), .B(n9263), .Z(n10211) );
  XNOR U10536 ( .A(n10212), .B(n10213), .Z(n9788) );
  XOR U10537 ( .A(n9304), .B(n10215), .Z(n10212) );
  XOR U10538 ( .A(key[808]), .B(n10216), .Z(n10215) );
  XNOR U10539 ( .A(n9776), .B(n10217), .Z(n8249) );
  XOR U10540 ( .A(n9795), .B(n9796), .Z(n10217) );
  IV U10541 ( .A(n9868), .Z(n9796) );
  XOR U10542 ( .A(n9861), .B(n10218), .Z(n9868) );
  XNOR U10543 ( .A(n10219), .B(n10220), .Z(n10218) );
  NANDN U10544 ( .A(n10221), .B(n9817), .Z(n10220) );
  XNOR U10545 ( .A(n9811), .B(n10222), .Z(n9861) );
  XNOR U10546 ( .A(n10223), .B(n10224), .Z(n10222) );
  NANDN U10547 ( .A(n10225), .B(n10226), .Z(n10224) );
  XOR U10548 ( .A(n10227), .B(n10228), .Z(n9795) );
  XNOR U10549 ( .A(n10229), .B(n10230), .Z(n10228) );
  NANDN U10550 ( .A(n10231), .B(n9822), .Z(n10230) );
  XOR U10551 ( .A(n9901), .B(n9860), .Z(n9776) );
  XNOR U10552 ( .A(n9811), .B(n10232), .Z(n9860) );
  XNOR U10553 ( .A(n10219), .B(n10233), .Z(n10232) );
  NANDN U10554 ( .A(n10234), .B(n10235), .Z(n10233) );
  OR U10555 ( .A(n10236), .B(n10237), .Z(n10219) );
  XOR U10556 ( .A(n10238), .B(n10223), .Z(n9811) );
  NANDN U10557 ( .A(n10239), .B(n10240), .Z(n10223) );
  ANDN U10558 ( .B(n10241), .A(n10242), .Z(n10238) );
  XNOR U10559 ( .A(n7039), .B(n10243), .Z(n9948) );
  XOR U10560 ( .A(key[1016]), .B(n9735), .Z(n10243) );
  IV U10561 ( .A(n6129), .Z(n9735) );
  XOR U10562 ( .A(n9818), .B(n9901), .Z(n6129) );
  XOR U10563 ( .A(n10227), .B(n10244), .Z(n9901) );
  XOR U10564 ( .A(n10245), .B(n9814), .Z(n10244) );
  OR U10565 ( .A(n10246), .B(n10236), .Z(n9814) );
  XNOR U10566 ( .A(n9817), .B(n10235), .Z(n10236) );
  ANDN U10567 ( .B(n10235), .A(n10247), .Z(n10245) );
  XNOR U10568 ( .A(n9812), .B(n10248), .Z(n9818) );
  XOR U10569 ( .A(n10249), .B(n10229), .Z(n10248) );
  NANDN U10570 ( .A(n10250), .B(n9865), .Z(n10229) );
  XNOR U10571 ( .A(n9867), .B(n9822), .Z(n9865) );
  ANDN U10572 ( .B(n10251), .A(n9867), .Z(n10249) );
  XNOR U10573 ( .A(n10227), .B(n10252), .Z(n9812) );
  XNOR U10574 ( .A(n10253), .B(n10254), .Z(n10252) );
  NANDN U10575 ( .A(n10225), .B(n10255), .Z(n10254) );
  XOR U10576 ( .A(n10256), .B(n10253), .Z(n10227) );
  OR U10577 ( .A(n10239), .B(n10257), .Z(n10253) );
  XNOR U10578 ( .A(n10242), .B(n10225), .Z(n10239) );
  XNOR U10579 ( .A(n10235), .B(n9822), .Z(n10225) );
  XOR U10580 ( .A(n10258), .B(n10259), .Z(n9822) );
  NANDN U10581 ( .A(n10260), .B(n10261), .Z(n10259) );
  XOR U10582 ( .A(n10262), .B(n10263), .Z(n10235) );
  NANDN U10583 ( .A(n10260), .B(n10264), .Z(n10263) );
  NOR U10584 ( .A(n10242), .B(n10265), .Z(n10256) );
  XOR U10585 ( .A(n9867), .B(n9817), .Z(n10242) );
  XNOR U10586 ( .A(n10266), .B(n10262), .Z(n9817) );
  NANDN U10587 ( .A(n10267), .B(n10268), .Z(n10262) );
  XOR U10588 ( .A(n10264), .B(n10269), .Z(n10268) );
  ANDN U10589 ( .B(n10269), .A(n10270), .Z(n10266) );
  XOR U10590 ( .A(n10271), .B(n10258), .Z(n9867) );
  NANDN U10591 ( .A(n10267), .B(n10272), .Z(n10258) );
  XOR U10592 ( .A(n10273), .B(n10261), .Z(n10272) );
  XNOR U10593 ( .A(n10274), .B(n10275), .Z(n10260) );
  XOR U10594 ( .A(n10276), .B(n10277), .Z(n10275) );
  XNOR U10595 ( .A(n10278), .B(n10279), .Z(n10274) );
  XNOR U10596 ( .A(n10280), .B(n10281), .Z(n10279) );
  ANDN U10597 ( .B(n10273), .A(n10277), .Z(n10280) );
  ANDN U10598 ( .B(n10273), .A(n10270), .Z(n10271) );
  XNOR U10599 ( .A(n10276), .B(n10282), .Z(n10270) );
  XOR U10600 ( .A(n10283), .B(n10281), .Z(n10282) );
  NAND U10601 ( .A(n10284), .B(n10285), .Z(n10281) );
  XNOR U10602 ( .A(n10278), .B(n10261), .Z(n10285) );
  IV U10603 ( .A(n10273), .Z(n10278) );
  XNOR U10604 ( .A(n10264), .B(n10277), .Z(n10284) );
  IV U10605 ( .A(n10269), .Z(n10277) );
  XOR U10606 ( .A(n10286), .B(n10287), .Z(n10269) );
  XNOR U10607 ( .A(n10288), .B(n10289), .Z(n10287) );
  XNOR U10608 ( .A(n10290), .B(n10291), .Z(n10286) );
  ANDN U10609 ( .B(n10251), .A(n10292), .Z(n10290) );
  AND U10610 ( .A(n10261), .B(n10264), .Z(n10283) );
  XNOR U10611 ( .A(n10261), .B(n10264), .Z(n10276) );
  XNOR U10612 ( .A(n10293), .B(n10294), .Z(n10264) );
  XNOR U10613 ( .A(n10295), .B(n10289), .Z(n10294) );
  XOR U10614 ( .A(n10296), .B(n10297), .Z(n10293) );
  XNOR U10615 ( .A(n10298), .B(n10291), .Z(n10297) );
  OR U10616 ( .A(n9864), .B(n10250), .Z(n10291) );
  XNOR U10617 ( .A(n10251), .B(n10299), .Z(n10250) );
  XNOR U10618 ( .A(n10292), .B(n9823), .Z(n9864) );
  ANDN U10619 ( .B(n10300), .A(n10231), .Z(n10298) );
  XNOR U10620 ( .A(n10301), .B(n10302), .Z(n10261) );
  XNOR U10621 ( .A(n10289), .B(n10303), .Z(n10302) );
  XOR U10622 ( .A(n10221), .B(n10296), .Z(n10303) );
  XNOR U10623 ( .A(n10251), .B(n10292), .Z(n10289) );
  XOR U10624 ( .A(n9816), .B(n10304), .Z(n10301) );
  XNOR U10625 ( .A(n10305), .B(n10306), .Z(n10304) );
  ANDN U10626 ( .B(n10307), .A(n10247), .Z(n10305) );
  XNOR U10627 ( .A(n10308), .B(n10309), .Z(n10273) );
  XNOR U10628 ( .A(n10295), .B(n10310), .Z(n10309) );
  XNOR U10629 ( .A(n10234), .B(n10288), .Z(n10310) );
  XOR U10630 ( .A(n10296), .B(n10311), .Z(n10288) );
  XNOR U10631 ( .A(n10312), .B(n10313), .Z(n10311) );
  NAND U10632 ( .A(n10255), .B(n10226), .Z(n10313) );
  XNOR U10633 ( .A(n10314), .B(n10312), .Z(n10296) );
  NANDN U10634 ( .A(n10257), .B(n10240), .Z(n10312) );
  XOR U10635 ( .A(n10241), .B(n10226), .Z(n10240) );
  XNOR U10636 ( .A(n10307), .B(n9823), .Z(n10226) );
  XOR U10637 ( .A(n10265), .B(n10255), .Z(n10257) );
  XNOR U10638 ( .A(n10247), .B(n10299), .Z(n10255) );
  ANDN U10639 ( .B(n10241), .A(n10265), .Z(n10314) );
  XOR U10640 ( .A(n9816), .B(n10251), .Z(n10265) );
  XNOR U10641 ( .A(n10315), .B(n10316), .Z(n10251) );
  XNOR U10642 ( .A(n10317), .B(n10318), .Z(n10316) );
  XOR U10643 ( .A(n10299), .B(n10300), .Z(n10295) );
  IV U10644 ( .A(n9823), .Z(n10300) );
  XOR U10645 ( .A(n10319), .B(n10320), .Z(n9823) );
  XNOR U10646 ( .A(n10321), .B(n10318), .Z(n10320) );
  IV U10647 ( .A(n10231), .Z(n10299) );
  XOR U10648 ( .A(n10318), .B(n10322), .Z(n10231) );
  XNOR U10649 ( .A(n10323), .B(n10324), .Z(n10308) );
  XNOR U10650 ( .A(n10325), .B(n10306), .Z(n10324) );
  OR U10651 ( .A(n10237), .B(n10246), .Z(n10306) );
  XNOR U10652 ( .A(n9816), .B(n10247), .Z(n10246) );
  IV U10653 ( .A(n10323), .Z(n10247) );
  XOR U10654 ( .A(n10221), .B(n10307), .Z(n10237) );
  IV U10655 ( .A(n10234), .Z(n10307) );
  XOR U10656 ( .A(n9866), .B(n10326), .Z(n10234) );
  XNOR U10657 ( .A(n10321), .B(n10315), .Z(n10326) );
  XOR U10658 ( .A(n10327), .B(n10328), .Z(n10315) );
  XOR U10659 ( .A(n9469), .B(n10329), .Z(n10328) );
  IV U10660 ( .A(n10292), .Z(n9866) );
  XOR U10661 ( .A(n10319), .B(n10330), .Z(n10292) );
  XOR U10662 ( .A(n10318), .B(n10331), .Z(n10330) );
  NOR U10663 ( .A(n10221), .B(n9816), .Z(n10325) );
  XOR U10664 ( .A(n10319), .B(n10332), .Z(n10221) );
  XOR U10665 ( .A(n10318), .B(n10333), .Z(n10332) );
  XOR U10666 ( .A(n10334), .B(n10335), .Z(n10318) );
  XNOR U10667 ( .A(n10336), .B(n10337), .Z(n10335) );
  XOR U10668 ( .A(n9816), .B(n10338), .Z(n10334) );
  XNOR U10669 ( .A(key[854]), .B(n10339), .Z(n10338) );
  IV U10670 ( .A(n10322), .Z(n10319) );
  XOR U10671 ( .A(n10340), .B(n10341), .Z(n10322) );
  XNOR U10672 ( .A(n10342), .B(n10343), .Z(n10341) );
  XNOR U10673 ( .A(key[853]), .B(n10344), .Z(n10340) );
  XOR U10674 ( .A(n10345), .B(n10346), .Z(n10323) );
  XNOR U10675 ( .A(n10333), .B(n10331), .Z(n10346) );
  XNOR U10676 ( .A(n10347), .B(n10348), .Z(n10331) );
  XOR U10677 ( .A(n10349), .B(n10350), .Z(n10348) );
  XOR U10678 ( .A(key[855]), .B(n10351), .Z(n10347) );
  XNOR U10679 ( .A(n10352), .B(n10353), .Z(n10333) );
  XNOR U10680 ( .A(n10354), .B(n10355), .Z(n10353) );
  XNOR U10681 ( .A(n10356), .B(n10357), .Z(n10352) );
  XOR U10682 ( .A(key[852]), .B(n10358), .Z(n10357) );
  XNOR U10683 ( .A(n9816), .B(n10317), .Z(n10345) );
  XOR U10684 ( .A(n10359), .B(n10360), .Z(n10317) );
  XOR U10685 ( .A(n10361), .B(n10362), .Z(n10360) );
  XOR U10686 ( .A(n10321), .B(n10363), .Z(n10362) );
  XOR U10687 ( .A(n10364), .B(n10365), .Z(n10321) );
  XNOR U10688 ( .A(n10366), .B(n9430), .Z(n10365) );
  XOR U10689 ( .A(key[849]), .B(n10367), .Z(n10364) );
  IV U10690 ( .A(n9476), .Z(n10367) );
  XOR U10691 ( .A(n9429), .B(n10368), .Z(n10359) );
  XOR U10692 ( .A(key[851]), .B(n10369), .Z(n10368) );
  XNOR U10693 ( .A(n10370), .B(n10371), .Z(n9816) );
  XOR U10694 ( .A(key[848]), .B(n10373), .Z(n10370) );
  XOR U10695 ( .A(n9739), .B(n10374), .Z(n7039) );
  XNOR U10696 ( .A(n9741), .B(n9742), .Z(n10374) );
  XNOR U10697 ( .A(n10376), .B(n10377), .Z(n10375) );
  OR U10698 ( .A(n9835), .B(n10378), .Z(n10377) );
  XOR U10699 ( .A(n9830), .B(n10379), .Z(n9770) );
  XNOR U10700 ( .A(n10380), .B(n10381), .Z(n10379) );
  NAND U10701 ( .A(n10382), .B(n9946), .Z(n10381) );
  XOR U10702 ( .A(n9942), .B(n10383), .Z(n9741) );
  XOR U10703 ( .A(n9940), .B(n10384), .Z(n10383) );
  NAND U10704 ( .A(n10385), .B(n9840), .Z(n10384) );
  XOR U10705 ( .A(n9774), .B(n9840), .Z(n9842) );
  XNOR U10706 ( .A(n9937), .B(n9727), .Z(n9739) );
  XNOR U10707 ( .A(n9830), .B(n10387), .Z(n9727) );
  XNOR U10708 ( .A(n10376), .B(n10388), .Z(n10387) );
  NANDN U10709 ( .A(n10389), .B(n10390), .Z(n10388) );
  OR U10710 ( .A(n10391), .B(n10392), .Z(n10376) );
  XNOR U10711 ( .A(n10393), .B(n10380), .Z(n9830) );
  NANDN U10712 ( .A(n10394), .B(n10395), .Z(n10380) );
  ANDN U10713 ( .B(n10396), .A(n10397), .Z(n10393) );
  XNOR U10714 ( .A(n9942), .B(n10398), .Z(n9937) );
  XOR U10715 ( .A(n10399), .B(n9833), .Z(n10398) );
  OR U10716 ( .A(n10400), .B(n10391), .Z(n9833) );
  XNOR U10717 ( .A(n9835), .B(n10389), .Z(n10391) );
  NOR U10718 ( .A(n10401), .B(n10389), .Z(n10399) );
  XOR U10719 ( .A(n10402), .B(n9944), .Z(n9942) );
  OR U10720 ( .A(n10394), .B(n10403), .Z(n9944) );
  XNOR U10721 ( .A(n10404), .B(n9946), .Z(n10394) );
  XNOR U10722 ( .A(n10389), .B(n9840), .Z(n9946) );
  XOR U10723 ( .A(n10405), .B(n10406), .Z(n9840) );
  NANDN U10724 ( .A(n10407), .B(n10408), .Z(n10406) );
  XNOR U10725 ( .A(n10409), .B(n10410), .Z(n10389) );
  OR U10726 ( .A(n10407), .B(n10411), .Z(n10410) );
  ANDN U10727 ( .B(n10404), .A(n10412), .Z(n10402) );
  IV U10728 ( .A(n10397), .Z(n10404) );
  XOR U10729 ( .A(n9835), .B(n9774), .Z(n10397) );
  XNOR U10730 ( .A(n10413), .B(n10405), .Z(n9774) );
  NANDN U10731 ( .A(n10414), .B(n10415), .Z(n10405) );
  ANDN U10732 ( .B(n10416), .A(n10417), .Z(n10413) );
  NANDN U10733 ( .A(n10414), .B(n10419), .Z(n10409) );
  XOR U10734 ( .A(n10420), .B(n10407), .Z(n10414) );
  XNOR U10735 ( .A(n10421), .B(n10422), .Z(n10407) );
  XOR U10736 ( .A(n10423), .B(n10416), .Z(n10422) );
  XNOR U10737 ( .A(n10424), .B(n10425), .Z(n10421) );
  XNOR U10738 ( .A(n10426), .B(n10427), .Z(n10425) );
  ANDN U10739 ( .B(n10416), .A(n10428), .Z(n10426) );
  IV U10740 ( .A(n10429), .Z(n10416) );
  ANDN U10741 ( .B(n10420), .A(n10428), .Z(n10418) );
  IV U10742 ( .A(n10424), .Z(n10428) );
  IV U10743 ( .A(n10417), .Z(n10420) );
  XNOR U10744 ( .A(n10423), .B(n10430), .Z(n10417) );
  XOR U10745 ( .A(n10431), .B(n10427), .Z(n10430) );
  NAND U10746 ( .A(n10419), .B(n10415), .Z(n10427) );
  XNOR U10747 ( .A(n10408), .B(n10429), .Z(n10415) );
  XOR U10748 ( .A(n10432), .B(n10433), .Z(n10429) );
  XOR U10749 ( .A(n10434), .B(n10435), .Z(n10433) );
  XNOR U10750 ( .A(n10390), .B(n10436), .Z(n10435) );
  XNOR U10751 ( .A(n10437), .B(n10438), .Z(n10432) );
  XNOR U10752 ( .A(n10439), .B(n10440), .Z(n10438) );
  ANDN U10753 ( .B(n10441), .A(n9836), .Z(n10439) );
  XNOR U10754 ( .A(n10424), .B(n10411), .Z(n10419) );
  XOR U10755 ( .A(n10442), .B(n10443), .Z(n10424) );
  XNOR U10756 ( .A(n10444), .B(n10436), .Z(n10443) );
  XOR U10757 ( .A(n10445), .B(n10446), .Z(n10436) );
  XNOR U10758 ( .A(n10447), .B(n10448), .Z(n10446) );
  NAND U10759 ( .A(n9947), .B(n10382), .Z(n10448) );
  XNOR U10760 ( .A(n10449), .B(n10450), .Z(n10442) );
  ANDN U10761 ( .B(n10451), .A(n9941), .Z(n10449) );
  ANDN U10762 ( .B(n10408), .A(n10411), .Z(n10431) );
  XOR U10763 ( .A(n10411), .B(n10408), .Z(n10423) );
  XNOR U10764 ( .A(n10452), .B(n10453), .Z(n10408) );
  XNOR U10765 ( .A(n10445), .B(n10454), .Z(n10453) );
  XOR U10766 ( .A(n10444), .B(n10378), .Z(n10454) );
  XOR U10767 ( .A(n9836), .B(n10455), .Z(n10452) );
  XNOR U10768 ( .A(n10456), .B(n10440), .Z(n10455) );
  OR U10769 ( .A(n10392), .B(n10400), .Z(n10440) );
  XNOR U10770 ( .A(n9836), .B(n10401), .Z(n10400) );
  XOR U10771 ( .A(n10378), .B(n10390), .Z(n10392) );
  ANDN U10772 ( .B(n10390), .A(n10401), .Z(n10456) );
  XOR U10773 ( .A(n10457), .B(n10458), .Z(n10411) );
  XOR U10774 ( .A(n10445), .B(n10434), .Z(n10458) );
  XOR U10775 ( .A(n10385), .B(n9841), .Z(n10434) );
  XOR U10776 ( .A(n10459), .B(n10447), .Z(n10445) );
  NANDN U10777 ( .A(n10403), .B(n10395), .Z(n10447) );
  XOR U10778 ( .A(n10396), .B(n10382), .Z(n10395) );
  XNOR U10779 ( .A(n10451), .B(n10460), .Z(n10390) );
  XOR U10780 ( .A(n10461), .B(n10462), .Z(n10460) );
  XOR U10781 ( .A(n10412), .B(n9947), .Z(n10403) );
  XNOR U10782 ( .A(n10401), .B(n10385), .Z(n9947) );
  IV U10783 ( .A(n10437), .Z(n10401) );
  XOR U10784 ( .A(n10463), .B(n10464), .Z(n10437) );
  XOR U10785 ( .A(n10465), .B(n10466), .Z(n10464) );
  XNOR U10786 ( .A(n9836), .B(n10467), .Z(n10463) );
  ANDN U10787 ( .B(n10396), .A(n10412), .Z(n10459) );
  XNOR U10788 ( .A(n9836), .B(n9941), .Z(n10412) );
  XOR U10789 ( .A(n10451), .B(n10441), .Z(n10396) );
  IV U10790 ( .A(n10378), .Z(n10441) );
  XOR U10791 ( .A(n10468), .B(n10469), .Z(n10378) );
  XOR U10792 ( .A(n10470), .B(n10466), .Z(n10469) );
  XNOR U10793 ( .A(n10471), .B(n10472), .Z(n10466) );
  XOR U10794 ( .A(n10473), .B(n10474), .Z(n10471) );
  XOR U10795 ( .A(key[892]), .B(n10475), .Z(n10474) );
  IV U10796 ( .A(n9775), .Z(n10451) );
  XOR U10797 ( .A(n10444), .B(n10476), .Z(n10457) );
  XNOR U10798 ( .A(n10477), .B(n10450), .Z(n10476) );
  OR U10799 ( .A(n9843), .B(n10386), .Z(n10450) );
  XNOR U10800 ( .A(n10478), .B(n10385), .Z(n10386) );
  XNOR U10801 ( .A(n9775), .B(n9841), .Z(n9843) );
  ANDN U10802 ( .B(n10385), .A(n9841), .Z(n10477) );
  XOR U10803 ( .A(n10468), .B(n10479), .Z(n9841) );
  XNOR U10804 ( .A(n10480), .B(n10470), .Z(n10479) );
  XOR U10805 ( .A(n10470), .B(n10468), .Z(n10385) );
  XNOR U10806 ( .A(n9941), .B(n9775), .Z(n10444) );
  XOR U10807 ( .A(n10468), .B(n10481), .Z(n9775) );
  XNOR U10808 ( .A(n10470), .B(n10465), .Z(n10481) );
  XOR U10809 ( .A(n10482), .B(n10483), .Z(n10465) );
  XNOR U10810 ( .A(n10484), .B(n10485), .Z(n10483) );
  XOR U10811 ( .A(key[895]), .B(n9611), .Z(n10482) );
  IV U10812 ( .A(n10486), .Z(n9611) );
  XNOR U10813 ( .A(n10487), .B(n10488), .Z(n10468) );
  XNOR U10814 ( .A(n10489), .B(n10490), .Z(n10488) );
  XOR U10815 ( .A(n10491), .B(n10492), .Z(n10487) );
  XNOR U10816 ( .A(key[893]), .B(n10493), .Z(n10492) );
  IV U10817 ( .A(n10478), .Z(n9941) );
  XNOR U10818 ( .A(n10462), .B(n10494), .Z(n10478) );
  XOR U10819 ( .A(n10495), .B(n10496), .Z(n10470) );
  XOR U10820 ( .A(n10497), .B(n10498), .Z(n10496) );
  XOR U10821 ( .A(n9836), .B(n10499), .Z(n10495) );
  XNOR U10822 ( .A(key[894]), .B(n9600), .Z(n10499) );
  XNOR U10823 ( .A(n10500), .B(n10501), .Z(n9836) );
  XOR U10824 ( .A(n10502), .B(n9593), .Z(n10501) );
  XOR U10825 ( .A(n9624), .B(n10503), .Z(n10500) );
  XOR U10826 ( .A(key[888]), .B(n10504), .Z(n10503) );
  XOR U10827 ( .A(n10505), .B(n10506), .Z(n10467) );
  XNOR U10828 ( .A(n10507), .B(n10508), .Z(n10506) );
  XOR U10829 ( .A(n10509), .B(n10480), .Z(n10508) );
  IV U10830 ( .A(n10461), .Z(n10480) );
  XNOR U10831 ( .A(n10510), .B(n10511), .Z(n10461) );
  XOR U10832 ( .A(n10512), .B(n10513), .Z(n10511) );
  XOR U10833 ( .A(n9634), .B(n10514), .Z(n10510) );
  XOR U10834 ( .A(key[889]), .B(n10515), .Z(n10514) );
  XNOR U10835 ( .A(n10516), .B(n10517), .Z(n10505) );
  XOR U10836 ( .A(key[891]), .B(n9636), .Z(n10517) );
  XOR U10837 ( .A(n10518), .B(n10519), .Z(n10462) );
  XNOR U10838 ( .A(n10520), .B(n10521), .Z(n10519) );
  XOR U10839 ( .A(n9622), .B(n10522), .Z(n10518) );
  XOR U10840 ( .A(key[890]), .B(n10523), .Z(n10522) );
  XOR U10841 ( .A(n3010), .B(n10524), .Z(n8708) );
  XNOR U10842 ( .A(key[1130]), .B(n3017), .Z(n10524) );
  XOR U10843 ( .A(n10525), .B(n10526), .Z(n3017) );
  XNOR U10844 ( .A(n8662), .B(n8591), .Z(n10526) );
  XNOR U10845 ( .A(n10527), .B(n10528), .Z(n8591) );
  XNOR U10846 ( .A(n10529), .B(n8511), .Z(n10528) );
  ANDN U10847 ( .B(n10530), .A(n10531), .Z(n8511) );
  ANDN U10848 ( .B(n10532), .A(n8701), .Z(n10529) );
  IV U10849 ( .A(n10533), .Z(n8701) );
  XNOR U10850 ( .A(n8509), .B(n10534), .Z(n8662) );
  XNOR U10851 ( .A(n10535), .B(n10536), .Z(n10534) );
  NANDN U10852 ( .A(n10537), .B(n9641), .Z(n10536) );
  XOR U10853 ( .A(n8660), .B(n8604), .Z(n10525) );
  XNOR U10854 ( .A(n10535), .B(n10539), .Z(n10538) );
  NANDN U10855 ( .A(n10540), .B(n8601), .Z(n10539) );
  OR U10856 ( .A(n9640), .B(n10541), .Z(n10535) );
  XNOR U10857 ( .A(n8601), .B(n9641), .Z(n9640) );
  XNOR U10858 ( .A(n8509), .B(n10542), .Z(n10527) );
  XNOR U10859 ( .A(n10543), .B(n10544), .Z(n10542) );
  NANDN U10860 ( .A(n8706), .B(n10545), .Z(n10544) );
  XOR U10861 ( .A(n10546), .B(n10543), .Z(n8509) );
  NANDN U10862 ( .A(n10547), .B(n10548), .Z(n10543) );
  ANDN U10863 ( .B(n10549), .A(n10550), .Z(n10546) );
  XOR U10864 ( .A(n8702), .B(n10551), .Z(n8660) );
  XOR U10865 ( .A(n8699), .B(n10552), .Z(n10551) );
  NANDN U10866 ( .A(n10553), .B(n8513), .Z(n10552) );
  XOR U10867 ( .A(n10533), .B(n8513), .Z(n10530) );
  XOR U10868 ( .A(n10555), .B(n8704), .Z(n8702) );
  OR U10869 ( .A(n10547), .B(n10556), .Z(n8704) );
  XNOR U10870 ( .A(n10550), .B(n8706), .Z(n10547) );
  XNOR U10871 ( .A(n9641), .B(n8513), .Z(n8706) );
  XOR U10872 ( .A(n10557), .B(n10558), .Z(n8513) );
  NANDN U10873 ( .A(n10559), .B(n10560), .Z(n10558) );
  XOR U10874 ( .A(n10561), .B(n10562), .Z(n9641) );
  NANDN U10875 ( .A(n10559), .B(n10563), .Z(n10562) );
  NOR U10876 ( .A(n10550), .B(n10564), .Z(n10555) );
  XNOR U10877 ( .A(n10533), .B(n8601), .Z(n10550) );
  XNOR U10878 ( .A(n10565), .B(n10561), .Z(n8601) );
  NANDN U10879 ( .A(n10566), .B(n10567), .Z(n10561) );
  XOR U10880 ( .A(n10563), .B(n10568), .Z(n10567) );
  ANDN U10881 ( .B(n10568), .A(n10569), .Z(n10565) );
  XNOR U10882 ( .A(n10570), .B(n10557), .Z(n10533) );
  NANDN U10883 ( .A(n10566), .B(n10571), .Z(n10557) );
  XOR U10884 ( .A(n10572), .B(n10560), .Z(n10571) );
  XNOR U10885 ( .A(n10573), .B(n10574), .Z(n10559) );
  XOR U10886 ( .A(n10575), .B(n10576), .Z(n10574) );
  XNOR U10887 ( .A(n10577), .B(n10578), .Z(n10573) );
  XNOR U10888 ( .A(n10579), .B(n10580), .Z(n10578) );
  ANDN U10889 ( .B(n10572), .A(n10576), .Z(n10579) );
  ANDN U10890 ( .B(n10572), .A(n10569), .Z(n10570) );
  XNOR U10891 ( .A(n10575), .B(n10581), .Z(n10569) );
  XOR U10892 ( .A(n10582), .B(n10580), .Z(n10581) );
  NAND U10893 ( .A(n10583), .B(n10584), .Z(n10580) );
  XNOR U10894 ( .A(n10577), .B(n10560), .Z(n10584) );
  IV U10895 ( .A(n10572), .Z(n10577) );
  XNOR U10896 ( .A(n10563), .B(n10576), .Z(n10583) );
  IV U10897 ( .A(n10568), .Z(n10576) );
  XOR U10898 ( .A(n10585), .B(n10586), .Z(n10568) );
  XNOR U10899 ( .A(n10587), .B(n10588), .Z(n10586) );
  XNOR U10900 ( .A(n10589), .B(n10590), .Z(n10585) );
  ANDN U10901 ( .B(n8700), .A(n10591), .Z(n10589) );
  AND U10902 ( .A(n10560), .B(n10563), .Z(n10582) );
  XNOR U10903 ( .A(n10560), .B(n10563), .Z(n10575) );
  XNOR U10904 ( .A(n10592), .B(n10593), .Z(n10563) );
  XNOR U10905 ( .A(n10594), .B(n10588), .Z(n10593) );
  XOR U10906 ( .A(n10595), .B(n10596), .Z(n10592) );
  XNOR U10907 ( .A(n10597), .B(n10590), .Z(n10596) );
  OR U10908 ( .A(n10531), .B(n10554), .Z(n10590) );
  XNOR U10909 ( .A(n8700), .B(n10598), .Z(n10554) );
  XNOR U10910 ( .A(n10591), .B(n8514), .Z(n10531) );
  ANDN U10911 ( .B(n10599), .A(n10553), .Z(n10597) );
  XNOR U10912 ( .A(n10600), .B(n10601), .Z(n10560) );
  XNOR U10913 ( .A(n10588), .B(n10602), .Z(n10601) );
  XOR U10914 ( .A(n10540), .B(n10595), .Z(n10602) );
  XNOR U10915 ( .A(n8700), .B(n10591), .Z(n10588) );
  XOR U10916 ( .A(n8600), .B(n10603), .Z(n10600) );
  XNOR U10917 ( .A(n10604), .B(n10605), .Z(n10603) );
  ANDN U10918 ( .B(n10606), .A(n9642), .Z(n10604) );
  XNOR U10919 ( .A(n10607), .B(n10608), .Z(n10572) );
  XNOR U10920 ( .A(n10594), .B(n10609), .Z(n10608) );
  XNOR U10921 ( .A(n10537), .B(n10587), .Z(n10609) );
  XOR U10922 ( .A(n10595), .B(n10610), .Z(n10587) );
  XNOR U10923 ( .A(n10611), .B(n10612), .Z(n10610) );
  NAND U10924 ( .A(n8707), .B(n10545), .Z(n10612) );
  XNOR U10925 ( .A(n10613), .B(n10611), .Z(n10595) );
  NANDN U10926 ( .A(n10556), .B(n10548), .Z(n10611) );
  XOR U10927 ( .A(n10549), .B(n10545), .Z(n10548) );
  XNOR U10928 ( .A(n10606), .B(n8514), .Z(n10545) );
  XOR U10929 ( .A(n10564), .B(n8707), .Z(n10556) );
  XNOR U10930 ( .A(n9642), .B(n10598), .Z(n8707) );
  ANDN U10931 ( .B(n10549), .A(n10564), .Z(n10613) );
  XOR U10932 ( .A(n8600), .B(n8700), .Z(n10564) );
  XNOR U10933 ( .A(n10614), .B(n10615), .Z(n8700) );
  XNOR U10934 ( .A(n10616), .B(n10617), .Z(n10615) );
  XOR U10935 ( .A(n10598), .B(n10599), .Z(n10594) );
  IV U10936 ( .A(n8514), .Z(n10599) );
  XOR U10937 ( .A(n10618), .B(n10619), .Z(n8514) );
  XNOR U10938 ( .A(n10620), .B(n10617), .Z(n10619) );
  IV U10939 ( .A(n10553), .Z(n10598) );
  XOR U10940 ( .A(n10617), .B(n10621), .Z(n10553) );
  XNOR U10941 ( .A(n10622), .B(n10623), .Z(n10607) );
  XNOR U10942 ( .A(n10624), .B(n10605), .Z(n10623) );
  OR U10943 ( .A(n10541), .B(n9639), .Z(n10605) );
  XNOR U10944 ( .A(n8600), .B(n9642), .Z(n9639) );
  IV U10945 ( .A(n10622), .Z(n9642) );
  XOR U10946 ( .A(n10540), .B(n10606), .Z(n10541) );
  IV U10947 ( .A(n10537), .Z(n10606) );
  XOR U10948 ( .A(n10532), .B(n10625), .Z(n10537) );
  XNOR U10949 ( .A(n10620), .B(n10614), .Z(n10625) );
  XOR U10950 ( .A(n10626), .B(n10627), .Z(n10614) );
  XOR U10951 ( .A(n7478), .B(n6403), .Z(n10627) );
  XNOR U10952 ( .A(n6447), .B(n7476), .Z(n6403) );
  XOR U10953 ( .A(n6452), .B(n6404), .Z(n7478) );
  IV U10954 ( .A(n7485), .Z(n6452) );
  XNOR U10955 ( .A(n10628), .B(n10629), .Z(n7485) );
  XOR U10956 ( .A(n10630), .B(n10631), .Z(n10629) );
  XNOR U10957 ( .A(n10632), .B(n10633), .Z(n10628) );
  XNOR U10958 ( .A(key[898]), .B(n6445), .Z(n10626) );
  IV U10959 ( .A(n10591), .Z(n10532) );
  XOR U10960 ( .A(n10618), .B(n10634), .Z(n10591) );
  XOR U10961 ( .A(n10617), .B(n10635), .Z(n10634) );
  NOR U10962 ( .A(n10540), .B(n8600), .Z(n10624) );
  XOR U10963 ( .A(n10618), .B(n10636), .Z(n10540) );
  XOR U10964 ( .A(n10617), .B(n10637), .Z(n10636) );
  XOR U10965 ( .A(n10638), .B(n10639), .Z(n10617) );
  XOR U10966 ( .A(n8600), .B(n6414), .Z(n10639) );
  XNOR U10967 ( .A(n8125), .B(n10640), .Z(n6414) );
  XOR U10968 ( .A(n6423), .B(n7464), .Z(n8125) );
  XOR U10969 ( .A(n10641), .B(n10642), .Z(n7464) );
  XOR U10970 ( .A(n10643), .B(n10644), .Z(n6423) );
  XNOR U10971 ( .A(n6421), .B(n10645), .Z(n10638) );
  XNOR U10972 ( .A(key[902]), .B(n7490), .Z(n10645) );
  XOR U10973 ( .A(n7494), .B(n6428), .Z(n7490) );
  XNOR U10974 ( .A(n10646), .B(n10647), .Z(n6428) );
  XOR U10975 ( .A(n10648), .B(n10649), .Z(n10647) );
  XOR U10976 ( .A(n10650), .B(n10633), .Z(n10646) );
  IV U10977 ( .A(n10621), .Z(n10618) );
  XOR U10978 ( .A(n10651), .B(n10652), .Z(n10621) );
  XOR U10979 ( .A(n8126), .B(n6420), .Z(n10652) );
  XOR U10980 ( .A(n8109), .B(n7466), .Z(n6420) );
  XNOR U10981 ( .A(n10653), .B(n10654), .Z(n7466) );
  XNOR U10982 ( .A(n10655), .B(n10656), .Z(n10654) );
  XOR U10983 ( .A(n10657), .B(n10658), .Z(n10653) );
  XOR U10984 ( .A(n10659), .B(n10660), .Z(n10658) );
  ANDN U10985 ( .B(n10661), .A(n10662), .Z(n10660) );
  XNOR U10986 ( .A(n10663), .B(n10664), .Z(n8109) );
  XOR U10987 ( .A(n10665), .B(n10666), .Z(n10664) );
  XNOR U10988 ( .A(n10667), .B(n10668), .Z(n10663) );
  XOR U10989 ( .A(n10669), .B(n10670), .Z(n10668) );
  ANDN U10990 ( .B(n10671), .A(n10672), .Z(n10670) );
  XNOR U10991 ( .A(key[901]), .B(n8121), .Z(n10651) );
  XOR U10992 ( .A(n6421), .B(n6416), .Z(n8121) );
  XNOR U10993 ( .A(n10673), .B(n10674), .Z(n10631) );
  XNOR U10994 ( .A(n10675), .B(n10676), .Z(n10674) );
  ANDN U10995 ( .B(n10677), .A(n10678), .Z(n10675) );
  XNOR U10996 ( .A(n10679), .B(n10680), .Z(n6421) );
  XOR U10997 ( .A(n10681), .B(n10682), .Z(n10622) );
  XNOR U10998 ( .A(n10637), .B(n10635), .Z(n10682) );
  XNOR U10999 ( .A(n10683), .B(n10684), .Z(n10635) );
  XNOR U11000 ( .A(n10640), .B(n6429), .Z(n10684) );
  XNOR U11001 ( .A(n8122), .B(n7461), .Z(n6429) );
  XNOR U11002 ( .A(n10685), .B(n10686), .Z(n7461) );
  XNOR U11003 ( .A(n10643), .B(n10656), .Z(n10686) );
  XNOR U11004 ( .A(n10687), .B(n10688), .Z(n10656) );
  XNOR U11005 ( .A(n10689), .B(n10690), .Z(n10688) );
  NANDN U11006 ( .A(n10691), .B(n10692), .Z(n10690) );
  XOR U11007 ( .A(n10693), .B(n10694), .Z(n10685) );
  XNOR U11008 ( .A(n10695), .B(n10696), .Z(n8122) );
  XNOR U11009 ( .A(n10697), .B(n10666), .Z(n10696) );
  XNOR U11010 ( .A(n10698), .B(n10699), .Z(n10666) );
  XNOR U11011 ( .A(n10700), .B(n10701), .Z(n10699) );
  NANDN U11012 ( .A(n10702), .B(n10703), .Z(n10701) );
  XOR U11013 ( .A(n10704), .B(n10641), .Z(n10695) );
  XNOR U11014 ( .A(n10705), .B(n8114), .Z(n10640) );
  XNOR U11015 ( .A(n10706), .B(n10707), .Z(n8114) );
  XNOR U11016 ( .A(n10680), .B(n10708), .Z(n10707) );
  XNOR U11017 ( .A(n10709), .B(n10710), .Z(n10706) );
  XNOR U11018 ( .A(key[903]), .B(n7494), .Z(n10683) );
  XNOR U11019 ( .A(n10711), .B(n10712), .Z(n10637) );
  XNOR U11020 ( .A(n6435), .B(n6433), .Z(n10712) );
  XOR U11021 ( .A(n8095), .B(n7449), .Z(n6433) );
  XNOR U11022 ( .A(n10713), .B(n6447), .Z(n7449) );
  XNOR U11023 ( .A(n10714), .B(n10693), .Z(n6447) );
  XOR U11024 ( .A(n7476), .B(n10665), .Z(n8095) );
  XOR U11025 ( .A(n10715), .B(n10716), .Z(n7476) );
  XNOR U11026 ( .A(n8119), .B(n8126), .Z(n6435) );
  XOR U11027 ( .A(n10717), .B(n10718), .Z(n8126) );
  XNOR U11028 ( .A(n10719), .B(n10708), .Z(n10718) );
  XNOR U11029 ( .A(n10720), .B(n10721), .Z(n10708) );
  XNOR U11030 ( .A(n10722), .B(n10723), .Z(n10721) );
  OR U11031 ( .A(n10724), .B(n10725), .Z(n10723) );
  XNOR U11032 ( .A(n10726), .B(n10727), .Z(n10717) );
  XNOR U11033 ( .A(n10728), .B(n10729), .Z(n10727) );
  ANDN U11034 ( .B(n10730), .A(n10731), .Z(n10729) );
  XNOR U11035 ( .A(n8108), .B(n10732), .Z(n10711) );
  XNOR U11036 ( .A(key[900]), .B(n7451), .Z(n10732) );
  XOR U11037 ( .A(n7494), .B(n6419), .Z(n7451) );
  XNOR U11038 ( .A(n10733), .B(n10734), .Z(n6419) );
  XNOR U11039 ( .A(n10735), .B(n10649), .Z(n10734) );
  XNOR U11040 ( .A(n10736), .B(n10737), .Z(n10649) );
  XNOR U11041 ( .A(n10738), .B(n10739), .Z(n10737) );
  OR U11042 ( .A(n10740), .B(n10741), .Z(n10739) );
  XOR U11043 ( .A(n10742), .B(n10743), .Z(n10733) );
  XOR U11044 ( .A(n10676), .B(n10744), .Z(n10743) );
  ANDN U11045 ( .B(n10745), .A(n10746), .Z(n10744) );
  ANDN U11046 ( .B(n10747), .A(n10748), .Z(n10676) );
  XNOR U11047 ( .A(n8600), .B(n10616), .Z(n10681) );
  XOR U11048 ( .A(n10749), .B(n10750), .Z(n10616) );
  XNOR U11049 ( .A(n10620), .B(n6450), .Z(n10751) );
  XOR U11050 ( .A(n10705), .B(n8108), .Z(n6450) );
  XNOR U11051 ( .A(n10726), .B(n6445), .Z(n8108) );
  IV U11052 ( .A(n8119), .Z(n10705) );
  XOR U11053 ( .A(n10752), .B(n10753), .Z(n10620) );
  XNOR U11054 ( .A(n6457), .B(n6446), .Z(n10753) );
  XOR U11055 ( .A(n7495), .B(n6455), .Z(n6446) );
  XOR U11056 ( .A(n10643), .B(n10754), .Z(n6455) );
  XOR U11057 ( .A(n10693), .B(n10755), .Z(n10754) );
  XOR U11058 ( .A(n10714), .B(n10756), .Z(n10643) );
  IV U11059 ( .A(n8098), .Z(n7495) );
  XOR U11060 ( .A(n10716), .B(n10757), .Z(n8098) );
  XNOR U11061 ( .A(n10704), .B(n10641), .Z(n10757) );
  XOR U11062 ( .A(n10758), .B(n10759), .Z(n10641) );
  XOR U11063 ( .A(key[897]), .B(n7484), .Z(n10752) );
  XNOR U11064 ( .A(n6445), .B(n6406), .Z(n7484) );
  XOR U11065 ( .A(n10760), .B(n10709), .Z(n6445) );
  XOR U11066 ( .A(n7483), .B(n6402), .Z(n6442) );
  XNOR U11067 ( .A(n10761), .B(n10762), .Z(n6402) );
  XOR U11068 ( .A(n10756), .B(n10644), .Z(n10762) );
  XNOR U11069 ( .A(n10763), .B(n10764), .Z(n10644) );
  XNOR U11070 ( .A(n10765), .B(n10659), .Z(n10764) );
  ANDN U11071 ( .B(n10766), .A(n10767), .Z(n10659) );
  ANDN U11072 ( .B(n10768), .A(n10769), .Z(n10765) );
  XOR U11073 ( .A(n10655), .B(n10770), .Z(n10756) );
  XNOR U11074 ( .A(n10771), .B(n10772), .Z(n10770) );
  NANDN U11075 ( .A(n10773), .B(n10774), .Z(n10772) );
  XNOR U11076 ( .A(n10693), .B(n10755), .Z(n10761) );
  IV U11077 ( .A(n10694), .Z(n10755) );
  XOR U11078 ( .A(n10763), .B(n10775), .Z(n10694) );
  XNOR U11079 ( .A(n10771), .B(n10776), .Z(n10775) );
  NANDN U11080 ( .A(n10777), .B(n10692), .Z(n10776) );
  OR U11081 ( .A(n10778), .B(n10779), .Z(n10771) );
  XNOR U11082 ( .A(n10655), .B(n10780), .Z(n10763) );
  XNOR U11083 ( .A(n10781), .B(n10782), .Z(n10780) );
  NANDN U11084 ( .A(n10783), .B(n10784), .Z(n10782) );
  XOR U11085 ( .A(n10785), .B(n10781), .Z(n10655) );
  NANDN U11086 ( .A(n10786), .B(n10787), .Z(n10781) );
  ANDN U11087 ( .B(n10788), .A(n10789), .Z(n10785) );
  XOR U11088 ( .A(n10790), .B(n10791), .Z(n10693) );
  XOR U11089 ( .A(n10792), .B(n10793), .Z(n10791) );
  NANDN U11090 ( .A(n10794), .B(n10661), .Z(n10793) );
  XOR U11091 ( .A(n10795), .B(n10796), .Z(n7483) );
  XNOR U11092 ( .A(n10697), .B(n10642), .Z(n10796) );
  XNOR U11093 ( .A(n10797), .B(n10798), .Z(n10642) );
  XNOR U11094 ( .A(n10799), .B(n10669), .Z(n10798) );
  NOR U11095 ( .A(n10800), .B(n10801), .Z(n10669) );
  ANDN U11096 ( .B(n10802), .A(n10803), .Z(n10799) );
  IV U11097 ( .A(n10716), .Z(n10697) );
  XOR U11098 ( .A(n10804), .B(n10805), .Z(n10716) );
  XOR U11099 ( .A(n10806), .B(n10807), .Z(n10805) );
  NANDN U11100 ( .A(n10808), .B(n10809), .Z(n10807) );
  XOR U11101 ( .A(n10704), .B(n10759), .Z(n10795) );
  XOR U11102 ( .A(n10667), .B(n10810), .Z(n10759) );
  XNOR U11103 ( .A(n10811), .B(n10812), .Z(n10810) );
  NANDN U11104 ( .A(n10813), .B(n10814), .Z(n10812) );
  XNOR U11105 ( .A(n10811), .B(n10816), .Z(n10815) );
  NAND U11106 ( .A(n10817), .B(n10703), .Z(n10816) );
  OR U11107 ( .A(n10818), .B(n10819), .Z(n10811) );
  XNOR U11108 ( .A(n10667), .B(n10820), .Z(n10797) );
  XNOR U11109 ( .A(n10821), .B(n10822), .Z(n10820) );
  OR U11110 ( .A(n10823), .B(n10824), .Z(n10822) );
  XOR U11111 ( .A(n10825), .B(n10821), .Z(n10667) );
  OR U11112 ( .A(n10826), .B(n10827), .Z(n10821) );
  ANDN U11113 ( .B(n10828), .A(n10829), .Z(n10825) );
  XOR U11114 ( .A(n6404), .B(n10830), .Z(n10749) );
  XNOR U11115 ( .A(key[899]), .B(n7480), .Z(n10830) );
  XOR U11116 ( .A(n7494), .B(n6437), .Z(n7480) );
  XNOR U11117 ( .A(n10735), .B(n6406), .Z(n6437) );
  XOR U11118 ( .A(n10650), .B(n10831), .Z(n6406) );
  XOR U11119 ( .A(n10831), .B(n10735), .Z(n7494) );
  XNOR U11120 ( .A(n10736), .B(n10832), .Z(n10735) );
  XNOR U11121 ( .A(n10833), .B(n10834), .Z(n10832) );
  ANDN U11122 ( .B(n10677), .A(n10835), .Z(n10833) );
  XNOR U11123 ( .A(n10836), .B(n10837), .Z(n10736) );
  XNOR U11124 ( .A(n10838), .B(n10839), .Z(n10837) );
  NAND U11125 ( .A(n10840), .B(n10841), .Z(n10839) );
  XNOR U11126 ( .A(n10842), .B(n10843), .Z(n6404) );
  XNOR U11127 ( .A(n10844), .B(n10679), .Z(n10843) );
  XNOR U11128 ( .A(n10845), .B(n10846), .Z(n10679) );
  XOR U11129 ( .A(n10847), .B(n10728), .Z(n10846) );
  NANDN U11130 ( .A(n10848), .B(n10849), .Z(n10728) );
  ANDN U11131 ( .B(n10850), .A(n10851), .Z(n10847) );
  XOR U11132 ( .A(n10709), .B(n10852), .Z(n10842) );
  XNOR U11133 ( .A(n10853), .B(n10854), .Z(n8600) );
  XOR U11134 ( .A(n10758), .B(n10665), .Z(n8094) );
  XOR U11135 ( .A(n10698), .B(n10855), .Z(n10665) );
  XNOR U11136 ( .A(n10856), .B(n10806), .Z(n10855) );
  NOR U11137 ( .A(n10800), .B(n10857), .Z(n10806) );
  XNOR U11138 ( .A(n10802), .B(n10809), .Z(n10800) );
  ANDN U11139 ( .B(n10802), .A(n10858), .Z(n10856) );
  XNOR U11140 ( .A(n10804), .B(n10859), .Z(n10698) );
  XNOR U11141 ( .A(n10860), .B(n10861), .Z(n10859) );
  NANDN U11142 ( .A(n10823), .B(n10862), .Z(n10861) );
  IV U11143 ( .A(n10715), .Z(n10758) );
  XNOR U11144 ( .A(n10804), .B(n10863), .Z(n10715) );
  XOR U11145 ( .A(n10864), .B(n10700), .Z(n10863) );
  OR U11146 ( .A(n10865), .B(n10818), .Z(n10700) );
  XNOR U11147 ( .A(n10703), .B(n10814), .Z(n10818) );
  ANDN U11148 ( .B(n10814), .A(n10866), .Z(n10864) );
  XOR U11149 ( .A(n10867), .B(n10860), .Z(n10804) );
  OR U11150 ( .A(n10826), .B(n10868), .Z(n10860) );
  XOR U11151 ( .A(n10828), .B(n10823), .Z(n10826) );
  XOR U11152 ( .A(n10814), .B(n10672), .Z(n10823) );
  IV U11153 ( .A(n10809), .Z(n10672) );
  XOR U11154 ( .A(n10869), .B(n10870), .Z(n10809) );
  NANDN U11155 ( .A(n10871), .B(n10872), .Z(n10870) );
  XOR U11156 ( .A(n10873), .B(n10874), .Z(n10814) );
  NANDN U11157 ( .A(n10871), .B(n10875), .Z(n10874) );
  AND U11158 ( .A(n10876), .B(n10828), .Z(n10867) );
  XOR U11159 ( .A(n10802), .B(n10703), .Z(n10828) );
  XNOR U11160 ( .A(n10877), .B(n10873), .Z(n10703) );
  NANDN U11161 ( .A(n10878), .B(n10879), .Z(n10873) );
  XOR U11162 ( .A(n10875), .B(n10880), .Z(n10879) );
  ANDN U11163 ( .B(n10880), .A(n10881), .Z(n10877) );
  NANDN U11164 ( .A(n10878), .B(n10883), .Z(n10869) );
  XOR U11165 ( .A(n10884), .B(n10872), .Z(n10883) );
  XNOR U11166 ( .A(n10885), .B(n10886), .Z(n10871) );
  XOR U11167 ( .A(n10887), .B(n10888), .Z(n10886) );
  XNOR U11168 ( .A(n10889), .B(n10890), .Z(n10885) );
  XNOR U11169 ( .A(n10891), .B(n10892), .Z(n10890) );
  ANDN U11170 ( .B(n10884), .A(n10888), .Z(n10891) );
  ANDN U11171 ( .B(n10884), .A(n10881), .Z(n10882) );
  XNOR U11172 ( .A(n10887), .B(n10893), .Z(n10881) );
  XOR U11173 ( .A(n10894), .B(n10892), .Z(n10893) );
  NAND U11174 ( .A(n10895), .B(n10896), .Z(n10892) );
  XNOR U11175 ( .A(n10889), .B(n10872), .Z(n10896) );
  IV U11176 ( .A(n10884), .Z(n10889) );
  XNOR U11177 ( .A(n10875), .B(n10888), .Z(n10895) );
  IV U11178 ( .A(n10880), .Z(n10888) );
  XOR U11179 ( .A(n10897), .B(n10898), .Z(n10880) );
  XNOR U11180 ( .A(n10899), .B(n10900), .Z(n10898) );
  XNOR U11181 ( .A(n10901), .B(n10902), .Z(n10897) );
  ANDN U11182 ( .B(n10903), .A(n10858), .Z(n10901) );
  AND U11183 ( .A(n10872), .B(n10875), .Z(n10894) );
  XNOR U11184 ( .A(n10872), .B(n10875), .Z(n10887) );
  XNOR U11185 ( .A(n10904), .B(n10905), .Z(n10875) );
  XNOR U11186 ( .A(n10906), .B(n10900), .Z(n10905) );
  XOR U11187 ( .A(n10907), .B(n10908), .Z(n10904) );
  XNOR U11188 ( .A(n10909), .B(n10902), .Z(n10908) );
  OR U11189 ( .A(n10801), .B(n10857), .Z(n10902) );
  XNOR U11190 ( .A(n10910), .B(n10941), .Z(n10857) );
  XNOR U11191 ( .A(n10803), .B(n10911), .Z(n10801) );
  ANDN U11192 ( .B(n10671), .A(n10808), .Z(n10909) );
  XNOR U11193 ( .A(n10912), .B(n10913), .Z(n10872) );
  XNOR U11194 ( .A(n10900), .B(n10914), .Z(n10913) );
  XNOR U11195 ( .A(n10817), .B(n10907), .Z(n10914) );
  XNOR U11196 ( .A(n10803), .B(n10910), .Z(n10900) );
  XNOR U11197 ( .A(n10915), .B(n10916), .Z(n10912) );
  XNOR U11198 ( .A(n10917), .B(n10918), .Z(n10916) );
  ANDN U11199 ( .B(n10919), .A(n10866), .Z(n10917) );
  XNOR U11200 ( .A(n10920), .B(n10921), .Z(n10884) );
  XNOR U11201 ( .A(n10906), .B(n10922), .Z(n10921) );
  XNOR U11202 ( .A(n10923), .B(n10899), .Z(n10922) );
  XOR U11203 ( .A(n10907), .B(n10924), .Z(n10899) );
  XNOR U11204 ( .A(n10925), .B(n10926), .Z(n10924) );
  NANDN U11205 ( .A(n10824), .B(n10862), .Z(n10926) );
  XNOR U11206 ( .A(n10927), .B(n10925), .Z(n10907) );
  OR U11207 ( .A(n10868), .B(n10827), .Z(n10925) );
  XOR U11208 ( .A(n10928), .B(n10824), .Z(n10827) );
  XNOR U11209 ( .A(n10671), .B(n10919), .Z(n10824) );
  IV U11210 ( .A(n10911), .Z(n10671) );
  XNOR U11211 ( .A(n10876), .B(n10862), .Z(n10868) );
  XNOR U11212 ( .A(n10866), .B(n10941), .Z(n10862) );
  IV U11213 ( .A(n10923), .Z(n10866) );
  ANDN U11214 ( .B(n10876), .A(n10829), .Z(n10927) );
  IV U11215 ( .A(n10928), .Z(n10829) );
  XOR U11216 ( .A(n10903), .B(n10817), .Z(n10928) );
  XOR U11217 ( .A(n10911), .B(n10808), .Z(n10906) );
  XOR U11218 ( .A(n10929), .B(n10930), .Z(n10808) );
  XOR U11219 ( .A(n10931), .B(n10932), .Z(n10911) );
  XOR U11220 ( .A(n10933), .B(n10930), .Z(n10932) );
  XNOR U11221 ( .A(n10813), .B(n10934), .Z(n10920) );
  XNOR U11222 ( .A(n10935), .B(n10918), .Z(n10934) );
  OR U11223 ( .A(n10819), .B(n10865), .Z(n10918) );
  XNOR U11224 ( .A(n10915), .B(n10923), .Z(n10865) );
  XOR U11225 ( .A(n10936), .B(n10937), .Z(n10923) );
  XNOR U11226 ( .A(n10938), .B(n10939), .Z(n10937) );
  XOR U11227 ( .A(n10915), .B(n10940), .Z(n10936) );
  XNOR U11228 ( .A(n10817), .B(n10919), .Z(n10819) );
  IV U11229 ( .A(n10813), .Z(n10919) );
  ANDN U11230 ( .B(n10817), .A(n10702), .Z(n10935) );
  XOR U11231 ( .A(n10938), .B(n10941), .Z(n10817) );
  XOR U11232 ( .A(n10942), .B(n10943), .Z(n10938) );
  XOR U11233 ( .A(n10356), .B(n10354), .Z(n10943) );
  XOR U11234 ( .A(n10944), .B(n9460), .Z(n10354) );
  IV U11235 ( .A(n10945), .Z(n9460) );
  XOR U11236 ( .A(n9478), .B(n10342), .Z(n10356) );
  XOR U11237 ( .A(n10946), .B(n10947), .Z(n10942) );
  XNOR U11238 ( .A(key[844]), .B(n9458), .Z(n10947) );
  XOR U11239 ( .A(n10948), .B(n10949), .Z(n9458) );
  XNOR U11240 ( .A(n10950), .B(n10951), .Z(n10813) );
  XOR U11241 ( .A(n10803), .B(n10931), .Z(n10951) );
  IV U11242 ( .A(n10903), .Z(n10803) );
  XOR U11243 ( .A(n10940), .B(n10941), .Z(n10903) );
  XNOR U11244 ( .A(n10929), .B(n10930), .Z(n10941) );
  IV U11245 ( .A(n10933), .Z(n10929) );
  XNOR U11246 ( .A(n10952), .B(n10953), .Z(n10933) );
  XNOR U11247 ( .A(n10954), .B(n10343), .Z(n10953) );
  XNOR U11248 ( .A(n10949), .B(n9446), .Z(n10343) );
  XNOR U11249 ( .A(n10955), .B(n10956), .Z(n10952) );
  XNOR U11250 ( .A(key[845]), .B(n10339), .Z(n10956) );
  XOR U11251 ( .A(n10957), .B(n10958), .Z(n10940) );
  XOR U11252 ( .A(n10372), .B(n10350), .Z(n10958) );
  XNOR U11253 ( .A(n10959), .B(n10960), .Z(n10350) );
  XNOR U11254 ( .A(key[847]), .B(n10961), .Z(n10957) );
  XOR U11255 ( .A(n10702), .B(n10858), .Z(n10876) );
  IV U11256 ( .A(n10910), .Z(n10858) );
  XNOR U11257 ( .A(n10939), .B(n10962), .Z(n10910) );
  XNOR U11258 ( .A(n10930), .B(n10950), .Z(n10962) );
  XOR U11259 ( .A(n10963), .B(n10964), .Z(n10950) );
  XOR U11260 ( .A(n10965), .B(n10966), .Z(n10964) );
  XOR U11261 ( .A(n9469), .B(n10967), .Z(n10963) );
  XNOR U11262 ( .A(n9431), .B(n10968), .Z(n9469) );
  XOR U11263 ( .A(n10969), .B(n10970), .Z(n10930) );
  XOR U11264 ( .A(n10336), .B(n10702), .Z(n10970) );
  XNOR U11265 ( .A(n9444), .B(n10349), .Z(n10336) );
  XOR U11266 ( .A(n9478), .B(n10971), .Z(n10349) );
  XOR U11267 ( .A(n10972), .B(n10955), .Z(n9444) );
  IV U11268 ( .A(n10973), .Z(n10955) );
  XNOR U11269 ( .A(n10974), .B(n10975), .Z(n10969) );
  XOR U11270 ( .A(key[846]), .B(n9440), .Z(n10975) );
  XOR U11271 ( .A(n9453), .B(n10959), .Z(n9440) );
  IV U11272 ( .A(n10976), .Z(n10959) );
  XOR U11273 ( .A(n10977), .B(n10978), .Z(n10939) );
  XOR U11274 ( .A(n10931), .B(n10979), .Z(n10978) );
  XNOR U11275 ( .A(n9429), .B(n10363), .Z(n10979) );
  XOR U11276 ( .A(n9473), .B(n10965), .Z(n9429) );
  IV U11277 ( .A(n10980), .Z(n10965) );
  IV U11278 ( .A(n10981), .Z(n9473) );
  XNOR U11279 ( .A(n10982), .B(n10983), .Z(n10931) );
  XNOR U11280 ( .A(n10984), .B(n10985), .Z(n10982) );
  XNOR U11281 ( .A(key[841]), .B(n9476), .Z(n10985) );
  XNOR U11282 ( .A(n10986), .B(n10987), .Z(n9476) );
  XNOR U11283 ( .A(n9465), .B(n10988), .Z(n10977) );
  XNOR U11284 ( .A(key[843]), .B(n10989), .Z(n10988) );
  XOR U11285 ( .A(n10948), .B(n10944), .Z(n9465) );
  IV U11286 ( .A(n10915), .Z(n10702) );
  XOR U11287 ( .A(n10990), .B(n10991), .Z(n10915) );
  XOR U11288 ( .A(n9477), .B(n10992), .Z(n10990) );
  XOR U11289 ( .A(n7496), .B(n6457), .Z(n7475) );
  XOR U11290 ( .A(n10680), .B(n10993), .Z(n6457) );
  XOR U11291 ( .A(n10709), .B(n10710), .Z(n10993) );
  IV U11292 ( .A(n10852), .Z(n10710) );
  XOR U11293 ( .A(n10845), .B(n10994), .Z(n10852) );
  XNOR U11294 ( .A(n10995), .B(n10996), .Z(n10994) );
  NANDN U11295 ( .A(n10724), .B(n10997), .Z(n10996) );
  XNOR U11296 ( .A(n10719), .B(n10998), .Z(n10845) );
  XNOR U11297 ( .A(n10999), .B(n11000), .Z(n10998) );
  NANDN U11298 ( .A(n11001), .B(n11002), .Z(n11000) );
  XOR U11299 ( .A(n11003), .B(n11004), .Z(n10709) );
  XNOR U11300 ( .A(n11005), .B(n11006), .Z(n11004) );
  NAND U11301 ( .A(n11007), .B(n10730), .Z(n11006) );
  XOR U11302 ( .A(n11008), .B(n10844), .Z(n10680) );
  XNOR U11303 ( .A(n10719), .B(n11009), .Z(n10844) );
  XNOR U11304 ( .A(n10995), .B(n11010), .Z(n11009) );
  NANDN U11305 ( .A(n11011), .B(n11012), .Z(n11010) );
  OR U11306 ( .A(n11013), .B(n11014), .Z(n10995) );
  XOR U11307 ( .A(n11015), .B(n10999), .Z(n10719) );
  NANDN U11308 ( .A(n11016), .B(n11017), .Z(n10999) );
  ANDN U11309 ( .B(n11018), .A(n11019), .Z(n11015) );
  IV U11310 ( .A(n6449), .Z(n7496) );
  XOR U11311 ( .A(n10648), .B(n11020), .Z(n6449) );
  XOR U11312 ( .A(n10632), .B(n10633), .Z(n11020) );
  XNOR U11313 ( .A(n11022), .B(n11023), .Z(n11021) );
  NANDN U11314 ( .A(n10740), .B(n11024), .Z(n11023) );
  XOR U11315 ( .A(n10742), .B(n11025), .Z(n10673) );
  XNOR U11316 ( .A(n11026), .B(n11027), .Z(n11025) );
  NAND U11317 ( .A(n11028), .B(n10840), .Z(n11027) );
  IV U11318 ( .A(n10650), .Z(n10632) );
  XOR U11319 ( .A(n10836), .B(n11029), .Z(n10650) );
  XOR U11320 ( .A(n10834), .B(n11030), .Z(n11029) );
  NAND U11321 ( .A(n11031), .B(n10745), .Z(n11030) );
  XOR U11322 ( .A(n10677), .B(n10745), .Z(n10747) );
  XOR U11323 ( .A(n10831), .B(n10630), .Z(n10648) );
  XNOR U11324 ( .A(n10742), .B(n11033), .Z(n10630) );
  XNOR U11325 ( .A(n11022), .B(n11034), .Z(n11033) );
  NANDN U11326 ( .A(n11035), .B(n11036), .Z(n11034) );
  OR U11327 ( .A(n11037), .B(n11038), .Z(n11022) );
  XNOR U11328 ( .A(n11039), .B(n11026), .Z(n10742) );
  NANDN U11329 ( .A(n11040), .B(n11041), .Z(n11026) );
  ANDN U11330 ( .B(n11042), .A(n11043), .Z(n11039) );
  XOR U11331 ( .A(n10836), .B(n11044), .Z(n10831) );
  XOR U11332 ( .A(n11045), .B(n10738), .Z(n11044) );
  OR U11333 ( .A(n11046), .B(n11037), .Z(n10738) );
  XNOR U11334 ( .A(n10740), .B(n11035), .Z(n11037) );
  NOR U11335 ( .A(n11047), .B(n11035), .Z(n11045) );
  XOR U11336 ( .A(n11048), .B(n10838), .Z(n10836) );
  OR U11337 ( .A(n11040), .B(n11049), .Z(n10838) );
  XNOR U11338 ( .A(n11050), .B(n10840), .Z(n11040) );
  XNOR U11339 ( .A(n11035), .B(n10745), .Z(n10840) );
  XOR U11340 ( .A(n11051), .B(n11052), .Z(n10745) );
  NANDN U11341 ( .A(n11053), .B(n11054), .Z(n11052) );
  XNOR U11342 ( .A(n11055), .B(n11056), .Z(n11035) );
  OR U11343 ( .A(n11053), .B(n11057), .Z(n11056) );
  ANDN U11344 ( .B(n11050), .A(n11058), .Z(n11048) );
  IV U11345 ( .A(n11043), .Z(n11050) );
  XOR U11346 ( .A(n10740), .B(n10677), .Z(n11043) );
  XNOR U11347 ( .A(n11059), .B(n11051), .Z(n10677) );
  NANDN U11348 ( .A(n11060), .B(n11061), .Z(n11051) );
  ANDN U11349 ( .B(n11062), .A(n11063), .Z(n11059) );
  NANDN U11350 ( .A(n11060), .B(n11065), .Z(n11055) );
  XOR U11351 ( .A(n11066), .B(n11053), .Z(n11060) );
  XNOR U11352 ( .A(n11067), .B(n11068), .Z(n11053) );
  XOR U11353 ( .A(n11069), .B(n11062), .Z(n11068) );
  XNOR U11354 ( .A(n11070), .B(n11071), .Z(n11067) );
  XNOR U11355 ( .A(n11072), .B(n11073), .Z(n11071) );
  ANDN U11356 ( .B(n11062), .A(n11074), .Z(n11072) );
  IV U11357 ( .A(n11075), .Z(n11062) );
  ANDN U11358 ( .B(n11066), .A(n11074), .Z(n11064) );
  IV U11359 ( .A(n11070), .Z(n11074) );
  IV U11360 ( .A(n11063), .Z(n11066) );
  XNOR U11361 ( .A(n11069), .B(n11076), .Z(n11063) );
  XOR U11362 ( .A(n11077), .B(n11073), .Z(n11076) );
  NAND U11363 ( .A(n11065), .B(n11061), .Z(n11073) );
  XNOR U11364 ( .A(n11054), .B(n11075), .Z(n11061) );
  XOR U11365 ( .A(n11078), .B(n11079), .Z(n11075) );
  XOR U11366 ( .A(n11080), .B(n11081), .Z(n11079) );
  XNOR U11367 ( .A(n11036), .B(n11082), .Z(n11081) );
  XNOR U11368 ( .A(n11083), .B(n11084), .Z(n11078) );
  XNOR U11369 ( .A(n11085), .B(n11086), .Z(n11084) );
  ANDN U11370 ( .B(n11024), .A(n10741), .Z(n11085) );
  XNOR U11371 ( .A(n11070), .B(n11057), .Z(n11065) );
  XOR U11372 ( .A(n11087), .B(n11088), .Z(n11070) );
  XNOR U11373 ( .A(n11089), .B(n11082), .Z(n11088) );
  XOR U11374 ( .A(n11090), .B(n11091), .Z(n11082) );
  XNOR U11375 ( .A(n11092), .B(n11093), .Z(n11091) );
  NAND U11376 ( .A(n10841), .B(n11028), .Z(n11093) );
  XNOR U11377 ( .A(n11094), .B(n11095), .Z(n11087) );
  ANDN U11378 ( .B(n11096), .A(n10835), .Z(n11094) );
  ANDN U11379 ( .B(n11054), .A(n11057), .Z(n11077) );
  XOR U11380 ( .A(n11057), .B(n11054), .Z(n11069) );
  XNOR U11381 ( .A(n11097), .B(n11098), .Z(n11054) );
  XNOR U11382 ( .A(n11090), .B(n11099), .Z(n11098) );
  XNOR U11383 ( .A(n11089), .B(n11024), .Z(n11099) );
  XNOR U11384 ( .A(n11100), .B(n11101), .Z(n11097) );
  XNOR U11385 ( .A(n11102), .B(n11086), .Z(n11101) );
  OR U11386 ( .A(n11038), .B(n11046), .Z(n11086) );
  XNOR U11387 ( .A(n11100), .B(n11083), .Z(n11046) );
  XNOR U11388 ( .A(n11024), .B(n11036), .Z(n11038) );
  ANDN U11389 ( .B(n11036), .A(n11047), .Z(n11102) );
  XOR U11390 ( .A(n11103), .B(n11104), .Z(n11057) );
  XOR U11391 ( .A(n11090), .B(n11080), .Z(n11104) );
  XOR U11392 ( .A(n11031), .B(n10746), .Z(n11080) );
  XOR U11393 ( .A(n11105), .B(n11092), .Z(n11090) );
  NANDN U11394 ( .A(n11049), .B(n11041), .Z(n11092) );
  XOR U11395 ( .A(n11042), .B(n11028), .Z(n11041) );
  XNOR U11396 ( .A(n11096), .B(n11106), .Z(n11036) );
  XNOR U11397 ( .A(n11107), .B(n11108), .Z(n11106) );
  XOR U11398 ( .A(n11058), .B(n10841), .Z(n11049) );
  XNOR U11399 ( .A(n11047), .B(n11031), .Z(n10841) );
  IV U11400 ( .A(n11083), .Z(n11047) );
  XOR U11401 ( .A(n11109), .B(n11110), .Z(n11083) );
  XOR U11402 ( .A(n11111), .B(n11112), .Z(n11110) );
  XOR U11403 ( .A(n11100), .B(n11113), .Z(n11109) );
  ANDN U11404 ( .B(n11042), .A(n11058), .Z(n11105) );
  XNOR U11405 ( .A(n11100), .B(n11114), .Z(n11058) );
  XOR U11406 ( .A(n11096), .B(n11024), .Z(n11042) );
  XNOR U11407 ( .A(n11115), .B(n11116), .Z(n11024) );
  XOR U11408 ( .A(n11117), .B(n11112), .Z(n11116) );
  XNOR U11409 ( .A(n11118), .B(n11119), .Z(n11112) );
  XOR U11410 ( .A(n9290), .B(n10194), .Z(n11119) );
  XOR U11411 ( .A(n10216), .B(n9276), .Z(n10194) );
  XNOR U11412 ( .A(n9294), .B(n11121), .Z(n11118) );
  XNOR U11413 ( .A(key[804]), .B(n11122), .Z(n11121) );
  XNOR U11414 ( .A(n11123), .B(n11124), .Z(n9294) );
  IV U11415 ( .A(n10678), .Z(n11096) );
  XOR U11416 ( .A(n11089), .B(n11125), .Z(n11103) );
  XNOR U11417 ( .A(n11126), .B(n11095), .Z(n11125) );
  OR U11418 ( .A(n10748), .B(n11032), .Z(n11095) );
  XNOR U11419 ( .A(n11114), .B(n11031), .Z(n11032) );
  XNOR U11420 ( .A(n10678), .B(n10746), .Z(n10748) );
  ANDN U11421 ( .B(n11031), .A(n10746), .Z(n11126) );
  XOR U11422 ( .A(n11115), .B(n11127), .Z(n10746) );
  XOR U11423 ( .A(n11107), .B(n11128), .Z(n11127) );
  XOR U11424 ( .A(n11117), .B(n11115), .Z(n11031) );
  XNOR U11425 ( .A(n10835), .B(n10678), .Z(n11089) );
  XOR U11426 ( .A(n11115), .B(n11129), .Z(n10678) );
  XNOR U11427 ( .A(n11117), .B(n11111), .Z(n11129) );
  XOR U11428 ( .A(n11130), .B(n11131), .Z(n11111) );
  XNOR U11429 ( .A(n11132), .B(n9286), .Z(n11131) );
  XNOR U11430 ( .A(key[807]), .B(n11134), .Z(n11130) );
  XNOR U11431 ( .A(n11135), .B(n11136), .Z(n11115) );
  XOR U11432 ( .A(n9277), .B(n11137), .Z(n11136) );
  XNOR U11433 ( .A(n10180), .B(n11138), .Z(n9277) );
  XNOR U11434 ( .A(key[805]), .B(n11124), .Z(n11135) );
  IV U11435 ( .A(n11114), .Z(n10835) );
  XNOR U11436 ( .A(n11108), .B(n11139), .Z(n11114) );
  XOR U11437 ( .A(n11113), .B(n11128), .Z(n11139) );
  IV U11438 ( .A(n11117), .Z(n11128) );
  XOR U11439 ( .A(n11140), .B(n11141), .Z(n11117) );
  XOR U11440 ( .A(n10174), .B(n10741), .Z(n11141) );
  IV U11441 ( .A(n11100), .Z(n10741) );
  XOR U11442 ( .A(n11142), .B(n11143), .Z(n11100) );
  XOR U11443 ( .A(n9287), .B(n10207), .Z(n11143) );
  XNOR U11444 ( .A(n9314), .B(n11123), .Z(n9287) );
  XNOR U11445 ( .A(n11134), .B(n9285), .Z(n10174) );
  XOR U11446 ( .A(n11145), .B(n11146), .Z(n11140) );
  XNOR U11447 ( .A(key[806]), .B(n9272), .Z(n11146) );
  XNOR U11448 ( .A(n11147), .B(n11132), .Z(n9272) );
  XNOR U11449 ( .A(n11123), .B(n11148), .Z(n11132) );
  XOR U11450 ( .A(n11149), .B(n11150), .Z(n11113) );
  XNOR U11451 ( .A(n11107), .B(n11151), .Z(n11150) );
  XNOR U11452 ( .A(n9261), .B(n10203), .Z(n11151) );
  XNOR U11453 ( .A(n10216), .B(n9292), .Z(n10203) );
  XOR U11454 ( .A(n11152), .B(n11153), .Z(n11107) );
  XNOR U11455 ( .A(n9303), .B(n10165), .Z(n11153) );
  XOR U11456 ( .A(key[801]), .B(n9316), .Z(n11152) );
  XNOR U11457 ( .A(n9299), .B(n11154), .Z(n11149) );
  XNOR U11458 ( .A(key[803]), .B(n9309), .Z(n11154) );
  XNOR U11459 ( .A(n11123), .B(n11122), .Z(n9309) );
  IV U11460 ( .A(n11155), .Z(n9299) );
  XOR U11461 ( .A(n11156), .B(n11157), .Z(n11108) );
  XNOR U11462 ( .A(key[802]), .B(n9306), .Z(n11156) );
  XOR U11463 ( .A(key[896]), .B(n6430), .Z(n10853) );
  XNOR U11464 ( .A(n8105), .B(n8119), .Z(n6430) );
  XOR U11465 ( .A(n11008), .B(n10726), .Z(n8119) );
  XNOR U11466 ( .A(n10720), .B(n11158), .Z(n10726) );
  XOR U11467 ( .A(n11159), .B(n11005), .Z(n11158) );
  NANDN U11468 ( .A(n11160), .B(n10849), .Z(n11005) );
  XOR U11469 ( .A(n10850), .B(n10730), .Z(n10849) );
  ANDN U11470 ( .B(n10850), .A(n11161), .Z(n11159) );
  XNOR U11471 ( .A(n11003), .B(n11162), .Z(n10720) );
  XNOR U11472 ( .A(n11163), .B(n11164), .Z(n11162) );
  NANDN U11473 ( .A(n11001), .B(n11165), .Z(n11164) );
  IV U11474 ( .A(n10760), .Z(n11008) );
  XNOR U11475 ( .A(n11003), .B(n11166), .Z(n10760) );
  XOR U11476 ( .A(n11167), .B(n10722), .Z(n11166) );
  OR U11477 ( .A(n11168), .B(n11013), .Z(n10722) );
  XNOR U11478 ( .A(n10724), .B(n11011), .Z(n11013) );
  NOR U11479 ( .A(n11169), .B(n11011), .Z(n11167) );
  XOR U11480 ( .A(n11170), .B(n11163), .Z(n11003) );
  OR U11481 ( .A(n11016), .B(n11171), .Z(n11163) );
  XOR U11482 ( .A(n11172), .B(n11001), .Z(n11016) );
  XOR U11483 ( .A(n11011), .B(n10730), .Z(n11001) );
  XOR U11484 ( .A(n11173), .B(n11174), .Z(n10730) );
  NANDN U11485 ( .A(n11175), .B(n11176), .Z(n11174) );
  XNOR U11486 ( .A(n11177), .B(n11178), .Z(n11011) );
  OR U11487 ( .A(n11175), .B(n11179), .Z(n11178) );
  ANDN U11488 ( .B(n11172), .A(n11180), .Z(n11170) );
  IV U11489 ( .A(n11019), .Z(n11172) );
  XOR U11490 ( .A(n10724), .B(n10850), .Z(n11019) );
  XNOR U11491 ( .A(n11181), .B(n11173), .Z(n10850) );
  NANDN U11492 ( .A(n11182), .B(n11183), .Z(n11173) );
  ANDN U11493 ( .B(n11184), .A(n11185), .Z(n11181) );
  NANDN U11494 ( .A(n11182), .B(n11187), .Z(n11177) );
  XOR U11495 ( .A(n11188), .B(n11175), .Z(n11182) );
  XNOR U11496 ( .A(n11189), .B(n11190), .Z(n11175) );
  XOR U11497 ( .A(n11191), .B(n11184), .Z(n11190) );
  XNOR U11498 ( .A(n11192), .B(n11193), .Z(n11189) );
  XNOR U11499 ( .A(n11194), .B(n11195), .Z(n11193) );
  ANDN U11500 ( .B(n11184), .A(n11196), .Z(n11194) );
  IV U11501 ( .A(n11197), .Z(n11184) );
  ANDN U11502 ( .B(n11188), .A(n11196), .Z(n11186) );
  IV U11503 ( .A(n11192), .Z(n11196) );
  IV U11504 ( .A(n11185), .Z(n11188) );
  XNOR U11505 ( .A(n11191), .B(n11198), .Z(n11185) );
  XOR U11506 ( .A(n11199), .B(n11195), .Z(n11198) );
  NAND U11507 ( .A(n11187), .B(n11183), .Z(n11195) );
  XNOR U11508 ( .A(n11176), .B(n11197), .Z(n11183) );
  XOR U11509 ( .A(n11200), .B(n11201), .Z(n11197) );
  XOR U11510 ( .A(n11202), .B(n11203), .Z(n11201) );
  XNOR U11511 ( .A(n11012), .B(n11204), .Z(n11203) );
  XNOR U11512 ( .A(n11205), .B(n11206), .Z(n11200) );
  XNOR U11513 ( .A(n11207), .B(n11208), .Z(n11206) );
  ANDN U11514 ( .B(n10997), .A(n10725), .Z(n11207) );
  XNOR U11515 ( .A(n11192), .B(n11179), .Z(n11187) );
  XOR U11516 ( .A(n11209), .B(n11210), .Z(n11192) );
  XNOR U11517 ( .A(n11211), .B(n11204), .Z(n11210) );
  XOR U11518 ( .A(n11212), .B(n11213), .Z(n11204) );
  XNOR U11519 ( .A(n11214), .B(n11215), .Z(n11213) );
  NAND U11520 ( .A(n11165), .B(n11002), .Z(n11215) );
  XNOR U11521 ( .A(n11216), .B(n11217), .Z(n11209) );
  ANDN U11522 ( .B(n11218), .A(n11161), .Z(n11216) );
  ANDN U11523 ( .B(n11176), .A(n11179), .Z(n11199) );
  XOR U11524 ( .A(n11179), .B(n11176), .Z(n11191) );
  XNOR U11525 ( .A(n11219), .B(n11220), .Z(n11176) );
  XNOR U11526 ( .A(n11212), .B(n11221), .Z(n11220) );
  XNOR U11527 ( .A(n11211), .B(n10997), .Z(n11221) );
  XNOR U11528 ( .A(n11222), .B(n11223), .Z(n11219) );
  XNOR U11529 ( .A(n11224), .B(n11208), .Z(n11223) );
  OR U11530 ( .A(n11014), .B(n11168), .Z(n11208) );
  XNOR U11531 ( .A(n11222), .B(n11205), .Z(n11168) );
  XNOR U11532 ( .A(n10997), .B(n11012), .Z(n11014) );
  ANDN U11533 ( .B(n11012), .A(n11169), .Z(n11224) );
  XOR U11534 ( .A(n11225), .B(n11226), .Z(n11179) );
  XOR U11535 ( .A(n11212), .B(n11202), .Z(n11226) );
  XOR U11536 ( .A(n11007), .B(n10731), .Z(n11202) );
  XOR U11537 ( .A(n11227), .B(n11214), .Z(n11212) );
  NANDN U11538 ( .A(n11171), .B(n11017), .Z(n11214) );
  XOR U11539 ( .A(n11018), .B(n11002), .Z(n11017) );
  XNOR U11540 ( .A(n11218), .B(n11228), .Z(n11012) );
  XNOR U11541 ( .A(n11229), .B(n11230), .Z(n11228) );
  XOR U11542 ( .A(n11180), .B(n11165), .Z(n11171) );
  XNOR U11543 ( .A(n11169), .B(n11007), .Z(n11165) );
  IV U11544 ( .A(n11205), .Z(n11169) );
  XOR U11545 ( .A(n11231), .B(n11232), .Z(n11205) );
  XOR U11546 ( .A(n11233), .B(n11234), .Z(n11232) );
  XOR U11547 ( .A(n11222), .B(n11235), .Z(n11231) );
  ANDN U11548 ( .B(n11018), .A(n11180), .Z(n11227) );
  XNOR U11549 ( .A(n11222), .B(n11236), .Z(n11180) );
  XOR U11550 ( .A(n11218), .B(n10997), .Z(n11018) );
  XNOR U11551 ( .A(n11237), .B(n11238), .Z(n10997) );
  XOR U11552 ( .A(n11239), .B(n11234), .Z(n11238) );
  XNOR U11553 ( .A(n11240), .B(n10036), .Z(n11234) );
  XOR U11554 ( .A(n11241), .B(n11242), .Z(n10036) );
  XNOR U11555 ( .A(n9130), .B(n11243), .Z(n11242) );
  XNOR U11556 ( .A(n11244), .B(n9172), .Z(n11241) );
  XOR U11557 ( .A(n11245), .B(n11246), .Z(n11240) );
  XNOR U11558 ( .A(key[796]), .B(n9128), .Z(n11246) );
  XNOR U11559 ( .A(n9142), .B(n11247), .Z(n9128) );
  IV U11560 ( .A(n10851), .Z(n11218) );
  XOR U11561 ( .A(n11211), .B(n11248), .Z(n11225) );
  XNOR U11562 ( .A(n11249), .B(n11217), .Z(n11248) );
  OR U11563 ( .A(n10848), .B(n11160), .Z(n11217) );
  XNOR U11564 ( .A(n11236), .B(n11007), .Z(n11160) );
  XNOR U11565 ( .A(n10851), .B(n10731), .Z(n10848) );
  ANDN U11566 ( .B(n11007), .A(n10731), .Z(n11249) );
  XOR U11567 ( .A(n11237), .B(n11250), .Z(n10731) );
  XOR U11568 ( .A(n11229), .B(n11251), .Z(n11250) );
  XOR U11569 ( .A(n11239), .B(n11237), .Z(n11007) );
  XNOR U11570 ( .A(n11161), .B(n10851), .Z(n11211) );
  XOR U11571 ( .A(n11237), .B(n11252), .Z(n10851) );
  XNOR U11572 ( .A(n11239), .B(n11233), .Z(n11252) );
  XOR U11573 ( .A(n11253), .B(n11254), .Z(n11233) );
  XOR U11574 ( .A(n10074), .B(n10050), .Z(n11254) );
  XNOR U11575 ( .A(n11255), .B(n11256), .Z(n10050) );
  XNOR U11576 ( .A(key[799]), .B(n11257), .Z(n11253) );
  XNOR U11577 ( .A(n11258), .B(n11259), .Z(n11237) );
  XNOR U11578 ( .A(n9135), .B(n11247), .Z(n10045) );
  XOR U11579 ( .A(n11260), .B(n11261), .Z(n11258) );
  XNOR U11580 ( .A(key[797]), .B(n11262), .Z(n11261) );
  IV U11581 ( .A(n11236), .Z(n11161) );
  XNOR U11582 ( .A(n11230), .B(n11263), .Z(n11236) );
  XOR U11583 ( .A(n11235), .B(n11251), .Z(n11263) );
  IV U11584 ( .A(n11239), .Z(n11251) );
  XOR U11585 ( .A(n11264), .B(n11265), .Z(n11239) );
  XOR U11586 ( .A(n10059), .B(n10725), .Z(n11265) );
  IV U11587 ( .A(n11222), .Z(n10725) );
  XOR U11588 ( .A(n11266), .B(n11267), .Z(n11222) );
  XNOR U11589 ( .A(n9171), .B(n10069), .Z(n11267) );
  XNOR U11590 ( .A(n11268), .B(n11269), .Z(n11266) );
  XOR U11591 ( .A(key[792]), .B(n9142), .Z(n11269) );
  XOR U11592 ( .A(n9137), .B(n10049), .Z(n10059) );
  XOR U11593 ( .A(n11270), .B(n11271), .Z(n10049) );
  XNOR U11594 ( .A(n11262), .B(n9154), .Z(n9137) );
  XNOR U11595 ( .A(n11272), .B(n11273), .Z(n11264) );
  XNOR U11596 ( .A(key[798]), .B(n9152), .Z(n11273) );
  XOR U11597 ( .A(n9142), .B(n11255), .Z(n9152) );
  XOR U11598 ( .A(n11274), .B(n11275), .Z(n11235) );
  XNOR U11599 ( .A(n11229), .B(n11276), .Z(n11275) );
  XOR U11600 ( .A(n9160), .B(n10064), .Z(n11276) );
  XOR U11601 ( .A(n11270), .B(n10039), .Z(n10064) );
  IV U11602 ( .A(n11277), .Z(n10039) );
  IV U11603 ( .A(n9172), .Z(n11270) );
  XOR U11604 ( .A(n9142), .B(n11243), .Z(n9160) );
  XOR U11605 ( .A(n11278), .B(n11279), .Z(n11229) );
  XOR U11606 ( .A(n11280), .B(n11281), .Z(n11279) );
  XNOR U11607 ( .A(n10055), .B(n11282), .Z(n11278) );
  XNOR U11608 ( .A(key[793]), .B(n9170), .Z(n11282) );
  XOR U11609 ( .A(n11283), .B(n11268), .Z(n9170) );
  XNOR U11610 ( .A(n11284), .B(n11285), .Z(n11274) );
  XOR U11611 ( .A(key[795]), .B(n9146), .Z(n11285) );
  XOR U11612 ( .A(n9161), .B(n11286), .Z(n9146) );
  IV U11613 ( .A(n11287), .Z(n9161) );
  XOR U11614 ( .A(n11288), .B(n11289), .Z(n11230) );
  XOR U11615 ( .A(n11286), .B(n10070), .Z(n11289) );
  IV U11616 ( .A(n11290), .Z(n11286) );
  XOR U11617 ( .A(n9166), .B(n11291), .Z(n11288) );
  XNOR U11618 ( .A(key[794]), .B(n11292), .Z(n11291) );
  XNOR U11619 ( .A(n9148), .B(n11281), .Z(n9166) );
  IV U11620 ( .A(n6459), .Z(n8105) );
  XOR U11621 ( .A(n10657), .B(n10714), .Z(n6459) );
  XNOR U11622 ( .A(n10790), .B(n11293), .Z(n10714) );
  XOR U11623 ( .A(n11294), .B(n10689), .Z(n11293) );
  OR U11624 ( .A(n11295), .B(n10778), .Z(n10689) );
  XNOR U11625 ( .A(n10692), .B(n10774), .Z(n10778) );
  ANDN U11626 ( .B(n11296), .A(n11297), .Z(n11294) );
  IV U11627 ( .A(n10713), .Z(n10657) );
  XNOR U11628 ( .A(n11299), .B(n10792), .Z(n11298) );
  XOR U11629 ( .A(n11301), .B(n10661), .Z(n10766) );
  ANDN U11630 ( .B(n11302), .A(n10769), .Z(n11299) );
  IV U11631 ( .A(n11301), .Z(n10769) );
  XNOR U11632 ( .A(n10790), .B(n11303), .Z(n10687) );
  XNOR U11633 ( .A(n11304), .B(n11305), .Z(n11303) );
  NANDN U11634 ( .A(n10783), .B(n11306), .Z(n11305) );
  XOR U11635 ( .A(n11307), .B(n11304), .Z(n10790) );
  OR U11636 ( .A(n10786), .B(n11308), .Z(n11304) );
  XNOR U11637 ( .A(n10789), .B(n10783), .Z(n10786) );
  XNOR U11638 ( .A(n10774), .B(n10661), .Z(n10783) );
  XOR U11639 ( .A(n11309), .B(n11310), .Z(n10661) );
  NANDN U11640 ( .A(n11311), .B(n11312), .Z(n11310) );
  IV U11641 ( .A(n11297), .Z(n10774) );
  XNOR U11642 ( .A(n11313), .B(n11314), .Z(n11297) );
  NANDN U11643 ( .A(n11311), .B(n11315), .Z(n11314) );
  NOR U11644 ( .A(n10789), .B(n11316), .Z(n11307) );
  XNOR U11645 ( .A(n11301), .B(n10692), .Z(n10789) );
  XNOR U11646 ( .A(n11317), .B(n11313), .Z(n10692) );
  NANDN U11647 ( .A(n11318), .B(n11319), .Z(n11313) );
  XOR U11648 ( .A(n11315), .B(n11320), .Z(n11319) );
  ANDN U11649 ( .B(n11320), .A(n11321), .Z(n11317) );
  XNOR U11650 ( .A(n11322), .B(n11309), .Z(n11301) );
  NANDN U11651 ( .A(n11318), .B(n11323), .Z(n11309) );
  XOR U11652 ( .A(n11324), .B(n11312), .Z(n11323) );
  XNOR U11653 ( .A(n11325), .B(n11326), .Z(n11311) );
  XOR U11654 ( .A(n11327), .B(n11328), .Z(n11326) );
  XNOR U11655 ( .A(n11329), .B(n11330), .Z(n11325) );
  XNOR U11656 ( .A(n11331), .B(n11332), .Z(n11330) );
  ANDN U11657 ( .B(n11324), .A(n11328), .Z(n11331) );
  ANDN U11658 ( .B(n11324), .A(n11321), .Z(n11322) );
  XNOR U11659 ( .A(n11327), .B(n11333), .Z(n11321) );
  XOR U11660 ( .A(n11334), .B(n11332), .Z(n11333) );
  NAND U11661 ( .A(n11335), .B(n11336), .Z(n11332) );
  XNOR U11662 ( .A(n11329), .B(n11312), .Z(n11336) );
  IV U11663 ( .A(n11324), .Z(n11329) );
  XNOR U11664 ( .A(n11315), .B(n11328), .Z(n11335) );
  IV U11665 ( .A(n11320), .Z(n11328) );
  XOR U11666 ( .A(n11337), .B(n11338), .Z(n11320) );
  XNOR U11667 ( .A(n11339), .B(n11340), .Z(n11338) );
  XNOR U11668 ( .A(n11341), .B(n11342), .Z(n11337) );
  ANDN U11669 ( .B(n11302), .A(n11343), .Z(n11341) );
  AND U11670 ( .A(n11312), .B(n11315), .Z(n11334) );
  XNOR U11671 ( .A(n11312), .B(n11315), .Z(n11327) );
  XNOR U11672 ( .A(n11344), .B(n11345), .Z(n11315) );
  XNOR U11673 ( .A(n11346), .B(n11340), .Z(n11345) );
  XOR U11674 ( .A(n11347), .B(n11348), .Z(n11344) );
  XNOR U11675 ( .A(n11349), .B(n11342), .Z(n11348) );
  OR U11676 ( .A(n10767), .B(n11300), .Z(n11342) );
  XNOR U11677 ( .A(n11302), .B(n11350), .Z(n11300) );
  XNOR U11678 ( .A(n11343), .B(n10662), .Z(n10767) );
  ANDN U11679 ( .B(n11351), .A(n10794), .Z(n11349) );
  XNOR U11680 ( .A(n11352), .B(n11353), .Z(n11312) );
  XNOR U11681 ( .A(n11340), .B(n11354), .Z(n11353) );
  XOR U11682 ( .A(n10777), .B(n11347), .Z(n11354) );
  XNOR U11683 ( .A(n11302), .B(n11343), .Z(n11340) );
  XNOR U11684 ( .A(n11355), .B(n11356), .Z(n11352) );
  XNOR U11685 ( .A(n11357), .B(n11358), .Z(n11356) );
  ANDN U11686 ( .B(n11296), .A(n10773), .Z(n11357) );
  XNOR U11687 ( .A(n11359), .B(n11360), .Z(n11324) );
  XNOR U11688 ( .A(n11346), .B(n11361), .Z(n11360) );
  XNOR U11689 ( .A(n10773), .B(n11339), .Z(n11361) );
  XOR U11690 ( .A(n11347), .B(n11362), .Z(n11339) );
  XNOR U11691 ( .A(n11363), .B(n11364), .Z(n11362) );
  NAND U11692 ( .A(n11306), .B(n10784), .Z(n11364) );
  XNOR U11693 ( .A(n11365), .B(n11363), .Z(n11347) );
  NANDN U11694 ( .A(n11308), .B(n10787), .Z(n11363) );
  XOR U11695 ( .A(n10788), .B(n10784), .Z(n10787) );
  XNOR U11696 ( .A(n11366), .B(n10662), .Z(n10784) );
  XOR U11697 ( .A(n11316), .B(n11306), .Z(n11308) );
  XOR U11698 ( .A(n11296), .B(n11350), .Z(n11306) );
  ANDN U11699 ( .B(n10788), .A(n11316), .Z(n11365) );
  XNOR U11700 ( .A(n11355), .B(n11302), .Z(n11316) );
  XNOR U11701 ( .A(n11367), .B(n11368), .Z(n11302) );
  XNOR U11702 ( .A(n11369), .B(n11370), .Z(n11368) );
  XOR U11703 ( .A(n11371), .B(n10768), .Z(n10788) );
  XOR U11704 ( .A(n11350), .B(n11351), .Z(n11346) );
  IV U11705 ( .A(n10662), .Z(n11351) );
  XOR U11706 ( .A(n11372), .B(n11373), .Z(n10662) );
  XNOR U11707 ( .A(n11374), .B(n11370), .Z(n11373) );
  IV U11708 ( .A(n10794), .Z(n11350) );
  XOR U11709 ( .A(n11370), .B(n11375), .Z(n10794) );
  XNOR U11710 ( .A(n11296), .B(n11376), .Z(n11359) );
  XNOR U11711 ( .A(n11377), .B(n11358), .Z(n11376) );
  OR U11712 ( .A(n10779), .B(n11295), .Z(n11358) );
  XNOR U11713 ( .A(n11355), .B(n11296), .Z(n11295) );
  XOR U11714 ( .A(n10777), .B(n11366), .Z(n10779) );
  IV U11715 ( .A(n10773), .Z(n11366) );
  XOR U11716 ( .A(n10768), .B(n11378), .Z(n10773) );
  XNOR U11717 ( .A(n11374), .B(n11367), .Z(n11378) );
  XOR U11718 ( .A(n11379), .B(n11380), .Z(n11367) );
  XNOR U11719 ( .A(n9633), .B(n10507), .Z(n11380) );
  IV U11720 ( .A(n11381), .Z(n9633) );
  XNOR U11721 ( .A(key[882]), .B(n9626), .Z(n11379) );
  IV U11722 ( .A(n11343), .Z(n10768) );
  XOR U11723 ( .A(n11372), .B(n11382), .Z(n11343) );
  XOR U11724 ( .A(n11370), .B(n11383), .Z(n11382) );
  ANDN U11725 ( .B(n11371), .A(n10691), .Z(n11377) );
  IV U11726 ( .A(n10777), .Z(n11371) );
  XOR U11727 ( .A(n11372), .B(n11384), .Z(n10777) );
  XOR U11728 ( .A(n11370), .B(n11385), .Z(n11384) );
  XOR U11729 ( .A(n11386), .B(n11387), .Z(n11370) );
  XOR U11730 ( .A(n10497), .B(n10691), .Z(n11387) );
  IV U11731 ( .A(n11355), .Z(n10691) );
  XOR U11732 ( .A(n10504), .B(n9591), .Z(n10497) );
  XOR U11733 ( .A(n9598), .B(n11388), .Z(n11386) );
  XNOR U11734 ( .A(key[886]), .B(n9606), .Z(n11388) );
  XNOR U11735 ( .A(n11389), .B(n11390), .Z(n9606) );
  IV U11736 ( .A(n11375), .Z(n11372) );
  XOR U11737 ( .A(n11391), .B(n11392), .Z(n11375) );
  XOR U11738 ( .A(n9597), .B(n11393), .Z(n11392) );
  XNOR U11739 ( .A(key[885]), .B(n11395), .Z(n11391) );
  XOR U11740 ( .A(n11396), .B(n11397), .Z(n11296) );
  XNOR U11741 ( .A(n11385), .B(n11383), .Z(n11397) );
  XNOR U11742 ( .A(n11398), .B(n11399), .Z(n11383) );
  XNOR U11743 ( .A(n11390), .B(n9592), .Z(n11399) );
  XOR U11744 ( .A(n10484), .B(n11400), .Z(n9592) );
  XOR U11745 ( .A(n11401), .B(n11402), .Z(n11390) );
  XNOR U11746 ( .A(n11403), .B(n11404), .Z(n11385) );
  XOR U11747 ( .A(n9578), .B(n10473), .Z(n11404) );
  XOR U11748 ( .A(n10504), .B(n9596), .Z(n10473) );
  XOR U11749 ( .A(n11405), .B(n11406), .Z(n9578) );
  XNOR U11750 ( .A(n9582), .B(n11407), .Z(n11403) );
  XNOR U11751 ( .A(key[884]), .B(n11408), .Z(n11407) );
  XOR U11752 ( .A(n11401), .B(n11395), .Z(n9582) );
  XOR U11753 ( .A(n11355), .B(n11369), .Z(n11396) );
  XOR U11754 ( .A(n11409), .B(n11410), .Z(n11369) );
  XNOR U11755 ( .A(n11374), .B(n11411), .Z(n11410) );
  XNOR U11756 ( .A(n9632), .B(n10509), .Z(n11411) );
  XOR U11757 ( .A(n10504), .B(n9580), .Z(n10509) );
  XOR U11758 ( .A(n11412), .B(n11413), .Z(n11374) );
  XOR U11759 ( .A(n9623), .B(n11414), .Z(n11413) );
  XOR U11760 ( .A(n9619), .B(n11415), .Z(n11409) );
  XNOR U11761 ( .A(key[883]), .B(n9629), .Z(n11415) );
  XOR U11762 ( .A(n11401), .B(n11408), .Z(n9629) );
  XOR U11763 ( .A(n11416), .B(n11417), .Z(n11355) );
  XOR U11764 ( .A(n9593), .B(n10513), .Z(n11417) );
  XNOR U11765 ( .A(n9612), .B(n11418), .Z(n9593) );
  XNOR U11766 ( .A(key[880]), .B(n11419), .Z(n11416) );
  XOR U11767 ( .A(n8640), .B(n8630), .Z(n3010) );
  IV U11768 ( .A(n8500), .Z(n8630) );
  XOR U11769 ( .A(n8562), .B(n11420), .Z(n8500) );
  XOR U11770 ( .A(n8559), .B(n11421), .Z(n11420) );
  NANDN U11771 ( .A(n11422), .B(n8544), .Z(n11421) );
  XOR U11772 ( .A(n8629), .B(n8544), .Z(n8626) );
  XNOR U11773 ( .A(n8562), .B(n11424), .Z(n8640) );
  XOR U11774 ( .A(n11425), .B(n8537), .Z(n11424) );
  OR U11775 ( .A(n11426), .B(n8644), .Z(n8537) );
  XNOR U11776 ( .A(n8540), .B(n8639), .Z(n8644) );
  ANDN U11777 ( .B(n8639), .A(n11427), .Z(n11425) );
  XOR U11778 ( .A(n11428), .B(n8564), .Z(n8562) );
  OR U11779 ( .A(n8651), .B(n11429), .Z(n8564) );
  XNOR U11780 ( .A(n8654), .B(n8566), .Z(n8651) );
  XNOR U11781 ( .A(n8639), .B(n8544), .Z(n8566) );
  XOR U11782 ( .A(n11430), .B(n11431), .Z(n8544) );
  NANDN U11783 ( .A(n11432), .B(n11433), .Z(n11431) );
  XOR U11784 ( .A(n11434), .B(n11435), .Z(n8639) );
  NANDN U11785 ( .A(n11432), .B(n11436), .Z(n11435) );
  NOR U11786 ( .A(n8654), .B(n11437), .Z(n11428) );
  XNOR U11787 ( .A(n8629), .B(n8540), .Z(n8654) );
  XNOR U11788 ( .A(n11438), .B(n11434), .Z(n8540) );
  NANDN U11789 ( .A(n11439), .B(n11440), .Z(n11434) );
  XOR U11790 ( .A(n11436), .B(n11441), .Z(n11440) );
  ANDN U11791 ( .B(n11441), .A(n11442), .Z(n11438) );
  XNOR U11792 ( .A(n11443), .B(n11430), .Z(n8629) );
  NANDN U11793 ( .A(n11439), .B(n11444), .Z(n11430) );
  XOR U11794 ( .A(n11445), .B(n11433), .Z(n11444) );
  XNOR U11795 ( .A(n11446), .B(n11447), .Z(n11432) );
  XOR U11796 ( .A(n11448), .B(n11449), .Z(n11447) );
  XNOR U11797 ( .A(n11450), .B(n11451), .Z(n11446) );
  XNOR U11798 ( .A(n11452), .B(n11453), .Z(n11451) );
  ANDN U11799 ( .B(n11445), .A(n11449), .Z(n11452) );
  ANDN U11800 ( .B(n11445), .A(n11442), .Z(n11443) );
  XNOR U11801 ( .A(n11448), .B(n11454), .Z(n11442) );
  XOR U11802 ( .A(n11455), .B(n11453), .Z(n11454) );
  NAND U11803 ( .A(n11456), .B(n11457), .Z(n11453) );
  XNOR U11804 ( .A(n11450), .B(n11433), .Z(n11457) );
  IV U11805 ( .A(n11445), .Z(n11450) );
  XNOR U11806 ( .A(n11436), .B(n11449), .Z(n11456) );
  IV U11807 ( .A(n11441), .Z(n11449) );
  XOR U11808 ( .A(n11458), .B(n11459), .Z(n11441) );
  XNOR U11809 ( .A(n11460), .B(n11461), .Z(n11459) );
  XNOR U11810 ( .A(n11462), .B(n11463), .Z(n11458) );
  ANDN U11811 ( .B(n8560), .A(n11464), .Z(n11462) );
  AND U11812 ( .A(n11433), .B(n11436), .Z(n11455) );
  XNOR U11813 ( .A(n11433), .B(n11436), .Z(n11448) );
  XNOR U11814 ( .A(n11465), .B(n11466), .Z(n11436) );
  XNOR U11815 ( .A(n11467), .B(n11461), .Z(n11466) );
  XOR U11816 ( .A(n11468), .B(n11469), .Z(n11465) );
  XNOR U11817 ( .A(n11470), .B(n11463), .Z(n11469) );
  OR U11818 ( .A(n8627), .B(n11423), .Z(n11463) );
  XNOR U11819 ( .A(n8560), .B(n11471), .Z(n11423) );
  XNOR U11820 ( .A(n11464), .B(n8545), .Z(n8627) );
  ANDN U11821 ( .B(n11472), .A(n11422), .Z(n11470) );
  XNOR U11822 ( .A(n11473), .B(n11474), .Z(n11433) );
  XNOR U11823 ( .A(n11461), .B(n11475), .Z(n11474) );
  XOR U11824 ( .A(n8643), .B(n11468), .Z(n11475) );
  XNOR U11825 ( .A(n8560), .B(n11464), .Z(n11461) );
  XOR U11826 ( .A(n8539), .B(n11476), .Z(n11473) );
  XNOR U11827 ( .A(n11477), .B(n11478), .Z(n11476) );
  ANDN U11828 ( .B(n11479), .A(n11427), .Z(n11477) );
  XNOR U11829 ( .A(n11480), .B(n11481), .Z(n11445) );
  XNOR U11830 ( .A(n11467), .B(n11482), .Z(n11481) );
  XNOR U11831 ( .A(n8638), .B(n11460), .Z(n11482) );
  XOR U11832 ( .A(n11468), .B(n11483), .Z(n11460) );
  XNOR U11833 ( .A(n11484), .B(n11485), .Z(n11483) );
  NAND U11834 ( .A(n8567), .B(n8649), .Z(n11485) );
  XNOR U11835 ( .A(n11486), .B(n11484), .Z(n11468) );
  NANDN U11836 ( .A(n11429), .B(n8652), .Z(n11484) );
  XOR U11837 ( .A(n8653), .B(n8649), .Z(n8652) );
  XNOR U11838 ( .A(n11479), .B(n8545), .Z(n8649) );
  XOR U11839 ( .A(n11437), .B(n8567), .Z(n11429) );
  XNOR U11840 ( .A(n11427), .B(n11471), .Z(n8567) );
  ANDN U11841 ( .B(n8653), .A(n11437), .Z(n11486) );
  XOR U11842 ( .A(n8539), .B(n8560), .Z(n11437) );
  XNOR U11843 ( .A(n11487), .B(n11488), .Z(n8560) );
  XNOR U11844 ( .A(n11489), .B(n11490), .Z(n11488) );
  XOR U11845 ( .A(n11471), .B(n11472), .Z(n11467) );
  IV U11846 ( .A(n8545), .Z(n11472) );
  XOR U11847 ( .A(n11491), .B(n11492), .Z(n8545) );
  XOR U11848 ( .A(n11493), .B(n11490), .Z(n11492) );
  IV U11849 ( .A(n11422), .Z(n11471) );
  XOR U11850 ( .A(n11490), .B(n11494), .Z(n11422) );
  XNOR U11851 ( .A(n11495), .B(n11496), .Z(n11480) );
  XNOR U11852 ( .A(n11497), .B(n11478), .Z(n11496) );
  OR U11853 ( .A(n8645), .B(n11426), .Z(n11478) );
  XNOR U11854 ( .A(n8539), .B(n11427), .Z(n11426) );
  IV U11855 ( .A(n11495), .Z(n11427) );
  XOR U11856 ( .A(n8643), .B(n11479), .Z(n8645) );
  IV U11857 ( .A(n8638), .Z(n11479) );
  XOR U11858 ( .A(n8628), .B(n11498), .Z(n8638) );
  XOR U11859 ( .A(n11499), .B(n11500), .Z(n11487) );
  XNOR U11860 ( .A(n6305), .B(n6263), .Z(n11500) );
  XNOR U11861 ( .A(n7220), .B(n6307), .Z(n6263) );
  XNOR U11862 ( .A(key[978]), .B(n7221), .Z(n11499) );
  XOR U11863 ( .A(n6312), .B(n6264), .Z(n7221) );
  IV U11864 ( .A(n7228), .Z(n6312) );
  XNOR U11865 ( .A(n11501), .B(n11502), .Z(n7228) );
  XOR U11866 ( .A(n11503), .B(n11504), .Z(n11502) );
  XNOR U11867 ( .A(n11505), .B(n11506), .Z(n11501) );
  IV U11868 ( .A(n11464), .Z(n8628) );
  XOR U11869 ( .A(n11491), .B(n11507), .Z(n11464) );
  XOR U11870 ( .A(n11490), .B(n11508), .Z(n11507) );
  NOR U11871 ( .A(n8643), .B(n8539), .Z(n11497) );
  XOR U11872 ( .A(n11491), .B(n11509), .Z(n8643) );
  XOR U11873 ( .A(n11490), .B(n11510), .Z(n11509) );
  XOR U11874 ( .A(n11511), .B(n11512), .Z(n11490) );
  XOR U11875 ( .A(n8539), .B(n6274), .Z(n11512) );
  XNOR U11876 ( .A(n8361), .B(n11513), .Z(n6274) );
  XOR U11877 ( .A(n6283), .B(n7201), .Z(n8361) );
  XOR U11878 ( .A(n11514), .B(n11515), .Z(n7201) );
  XOR U11879 ( .A(n11516), .B(n11517), .Z(n6283) );
  XNOR U11880 ( .A(n11518), .B(n11519), .Z(n11517) );
  XNOR U11881 ( .A(n6281), .B(n11520), .Z(n11511) );
  XNOR U11882 ( .A(key[982]), .B(n7209), .Z(n11520) );
  XOR U11883 ( .A(n7231), .B(n6288), .Z(n7209) );
  XNOR U11884 ( .A(n11521), .B(n11522), .Z(n6288) );
  XOR U11885 ( .A(n11523), .B(n11524), .Z(n11522) );
  XOR U11886 ( .A(n11525), .B(n11506), .Z(n11521) );
  IV U11887 ( .A(n11494), .Z(n11491) );
  XOR U11888 ( .A(n11526), .B(n11527), .Z(n11494) );
  XOR U11889 ( .A(n8362), .B(n6280), .Z(n11527) );
  XOR U11890 ( .A(n8363), .B(n7203), .Z(n6280) );
  XNOR U11891 ( .A(n11528), .B(n11529), .Z(n7203) );
  XNOR U11892 ( .A(n11530), .B(n11531), .Z(n11529) );
  XNOR U11893 ( .A(n11532), .B(n11533), .Z(n11528) );
  XNOR U11894 ( .A(n11534), .B(n11535), .Z(n11533) );
  ANDN U11895 ( .B(n11536), .A(n11537), .Z(n11534) );
  XNOR U11896 ( .A(n11538), .B(n11539), .Z(n8363) );
  XOR U11897 ( .A(n11540), .B(n11541), .Z(n11539) );
  XNOR U11898 ( .A(n11542), .B(n11543), .Z(n11538) );
  XOR U11899 ( .A(n11544), .B(n11545), .Z(n11543) );
  ANDN U11900 ( .B(n11546), .A(n11547), .Z(n11545) );
  XNOR U11901 ( .A(key[981]), .B(n8357), .Z(n11526) );
  XOR U11902 ( .A(n6281), .B(n6276), .Z(n8357) );
  XNOR U11903 ( .A(n11548), .B(n11549), .Z(n11504) );
  XNOR U11904 ( .A(n11550), .B(n11551), .Z(n11549) );
  ANDN U11905 ( .B(n11552), .A(n11553), .Z(n11550) );
  XNOR U11906 ( .A(n11554), .B(n11555), .Z(n6281) );
  XNOR U11907 ( .A(n11556), .B(n11557), .Z(n11555) );
  XOR U11908 ( .A(n11558), .B(n11559), .Z(n11495) );
  XNOR U11909 ( .A(n11510), .B(n11508), .Z(n11559) );
  XNOR U11910 ( .A(n11560), .B(n11561), .Z(n11508) );
  XNOR U11911 ( .A(n11513), .B(n6289), .Z(n11561) );
  XNOR U11912 ( .A(n8370), .B(n7198), .Z(n6289) );
  XNOR U11913 ( .A(n11562), .B(n11563), .Z(n7198) );
  XNOR U11914 ( .A(n11564), .B(n11531), .Z(n11563) );
  XNOR U11915 ( .A(n11565), .B(n11566), .Z(n11531) );
  XNOR U11916 ( .A(n11567), .B(n11568), .Z(n11566) );
  OR U11917 ( .A(n11569), .B(n11570), .Z(n11568) );
  XOR U11918 ( .A(n11571), .B(n11572), .Z(n11562) );
  XNOR U11919 ( .A(n11573), .B(n11574), .Z(n8370) );
  XNOR U11920 ( .A(n11575), .B(n11541), .Z(n11574) );
  XNOR U11921 ( .A(n11576), .B(n11577), .Z(n11541) );
  XNOR U11922 ( .A(n11578), .B(n11579), .Z(n11577) );
  NANDN U11923 ( .A(n11580), .B(n11581), .Z(n11579) );
  XOR U11924 ( .A(n11582), .B(n11514), .Z(n11573) );
  XNOR U11925 ( .A(n11583), .B(n11584), .Z(n8368) );
  XNOR U11926 ( .A(n11585), .B(n11586), .Z(n11584) );
  XNOR U11927 ( .A(n11587), .B(n11588), .Z(n11583) );
  XNOR U11928 ( .A(key[983]), .B(n7231), .Z(n11560) );
  XNOR U11929 ( .A(n11589), .B(n11590), .Z(n11510) );
  XNOR U11930 ( .A(n6295), .B(n6293), .Z(n11590) );
  XOR U11931 ( .A(n11532), .B(n6307), .Z(n7186) );
  XNOR U11932 ( .A(n11518), .B(n11571), .Z(n6307) );
  XOR U11933 ( .A(n7220), .B(n11540), .Z(n8375) );
  XOR U11934 ( .A(n11591), .B(n11592), .Z(n7220) );
  XNOR U11935 ( .A(n8385), .B(n8362), .Z(n6295) );
  XOR U11936 ( .A(n11593), .B(n11594), .Z(n8362) );
  XNOR U11937 ( .A(n11595), .B(n11586), .Z(n11594) );
  XNOR U11938 ( .A(n11596), .B(n11597), .Z(n11586) );
  XNOR U11939 ( .A(n11598), .B(n11599), .Z(n11597) );
  OR U11940 ( .A(n11600), .B(n11601), .Z(n11599) );
  XNOR U11941 ( .A(n11602), .B(n11603), .Z(n11593) );
  XNOR U11942 ( .A(n11604), .B(n11605), .Z(n11603) );
  ANDN U11943 ( .B(n11606), .A(n11607), .Z(n11605) );
  XNOR U11944 ( .A(n8373), .B(n11608), .Z(n11589) );
  XNOR U11945 ( .A(key[980]), .B(n7188), .Z(n11608) );
  XOR U11946 ( .A(n7231), .B(n6279), .Z(n7188) );
  XNOR U11947 ( .A(n11609), .B(n11610), .Z(n6279) );
  XNOR U11948 ( .A(n11611), .B(n11524), .Z(n11610) );
  XNOR U11949 ( .A(n11612), .B(n11613), .Z(n11524) );
  XNOR U11950 ( .A(n11614), .B(n11615), .Z(n11613) );
  OR U11951 ( .A(n11616), .B(n11617), .Z(n11615) );
  XOR U11952 ( .A(n11618), .B(n11619), .Z(n11609) );
  XOR U11953 ( .A(n11551), .B(n11620), .Z(n11619) );
  ANDN U11954 ( .B(n11621), .A(n11622), .Z(n11620) );
  ANDN U11955 ( .B(n11623), .A(n11624), .Z(n11551) );
  XNOR U11956 ( .A(n8539), .B(n11489), .Z(n11558) );
  XOR U11957 ( .A(n11625), .B(n11626), .Z(n11489) );
  XNOR U11958 ( .A(n6302), .B(n11627), .Z(n11626) );
  XOR U11959 ( .A(n6310), .B(n11493), .Z(n11627) );
  XNOR U11960 ( .A(n11628), .B(n11629), .Z(n11493) );
  XNOR U11961 ( .A(n7226), .B(n6306), .Z(n11629) );
  XOR U11962 ( .A(n7232), .B(n6315), .Z(n6306) );
  XOR U11963 ( .A(n11564), .B(n11630), .Z(n6315) );
  IV U11964 ( .A(n8381), .Z(n7232) );
  XOR U11965 ( .A(n11592), .B(n11631), .Z(n8381) );
  XNOR U11966 ( .A(n11582), .B(n11514), .Z(n11631) );
  XOR U11967 ( .A(n11632), .B(n11633), .Z(n11514) );
  XNOR U11968 ( .A(n6262), .B(n6305), .Z(n7226) );
  XOR U11969 ( .A(key[977]), .B(n6317), .Z(n11628) );
  IV U11970 ( .A(n8348), .Z(n6310) );
  XOR U11971 ( .A(n6266), .B(n7225), .Z(n8348) );
  XOR U11972 ( .A(n11634), .B(n11635), .Z(n7225) );
  XNOR U11973 ( .A(n11575), .B(n11515), .Z(n11635) );
  XNOR U11974 ( .A(n11636), .B(n11637), .Z(n11515) );
  XNOR U11975 ( .A(n11638), .B(n11544), .Z(n11637) );
  NOR U11976 ( .A(n11639), .B(n11640), .Z(n11544) );
  ANDN U11977 ( .B(n11641), .A(n11642), .Z(n11638) );
  IV U11978 ( .A(n11592), .Z(n11575) );
  XOR U11979 ( .A(n11643), .B(n11644), .Z(n11592) );
  XOR U11980 ( .A(n11645), .B(n11646), .Z(n11644) );
  NANDN U11981 ( .A(n11647), .B(n11648), .Z(n11646) );
  XOR U11982 ( .A(n11582), .B(n11633), .Z(n11634) );
  XOR U11983 ( .A(n11542), .B(n11649), .Z(n11633) );
  XNOR U11984 ( .A(n11650), .B(n11651), .Z(n11649) );
  NANDN U11985 ( .A(n11652), .B(n11653), .Z(n11651) );
  XNOR U11986 ( .A(n11650), .B(n11655), .Z(n11654) );
  NAND U11987 ( .A(n11656), .B(n11581), .Z(n11655) );
  OR U11988 ( .A(n11657), .B(n11658), .Z(n11650) );
  XNOR U11989 ( .A(n11542), .B(n11659), .Z(n11636) );
  XNOR U11990 ( .A(n11660), .B(n11661), .Z(n11659) );
  OR U11991 ( .A(n11662), .B(n11663), .Z(n11661) );
  XOR U11992 ( .A(n11664), .B(n11660), .Z(n11542) );
  OR U11993 ( .A(n11665), .B(n11666), .Z(n11660) );
  ANDN U11994 ( .B(n11667), .A(n11668), .Z(n11664) );
  XOR U11995 ( .A(n11669), .B(n11630), .Z(n6266) );
  XNOR U11996 ( .A(n11571), .B(n11572), .Z(n11630) );
  XOR U11997 ( .A(n11670), .B(n11671), .Z(n11572) );
  XNOR U11998 ( .A(n11672), .B(n11673), .Z(n11671) );
  NANDN U11999 ( .A(n11569), .B(n11674), .Z(n11673) );
  XOR U12000 ( .A(n11675), .B(n11676), .Z(n11571) );
  XOR U12001 ( .A(n11677), .B(n11678), .Z(n11676) );
  NAND U12002 ( .A(n11679), .B(n11536), .Z(n11678) );
  XOR U12003 ( .A(n11519), .B(n11516), .Z(n11669) );
  XNOR U12004 ( .A(n11530), .B(n11680), .Z(n11516) );
  XOR U12005 ( .A(n11681), .B(n11672), .Z(n11680) );
  OR U12006 ( .A(n11682), .B(n11683), .Z(n11672) );
  AND U12007 ( .A(n11684), .B(n11685), .Z(n11681) );
  XNOR U12008 ( .A(n11670), .B(n11686), .Z(n11519) );
  XNOR U12009 ( .A(n11535), .B(n11687), .Z(n11686) );
  NANDN U12010 ( .A(n11688), .B(n11689), .Z(n11687) );
  NANDN U12011 ( .A(n11690), .B(n11691), .Z(n11535) );
  XNOR U12012 ( .A(n11530), .B(n11692), .Z(n11670) );
  XNOR U12013 ( .A(n11693), .B(n11694), .Z(n11692) );
  NANDN U12014 ( .A(n11695), .B(n11696), .Z(n11694) );
  XOR U12015 ( .A(n11697), .B(n11693), .Z(n11530) );
  NANDN U12016 ( .A(n11698), .B(n11699), .Z(n11693) );
  ANDN U12017 ( .B(n11700), .A(n11701), .Z(n11697) );
  XNOR U12018 ( .A(n8385), .B(n8373), .Z(n6302) );
  XOR U12019 ( .A(n11602), .B(n6305), .Z(n8373) );
  XNOR U12020 ( .A(n11702), .B(n11588), .Z(n6305) );
  XNOR U12021 ( .A(n7215), .B(n11703), .Z(n11625) );
  XOR U12022 ( .A(key[979]), .B(n6264), .Z(n11703) );
  XNOR U12023 ( .A(n11704), .B(n11705), .Z(n6264) );
  XOR U12024 ( .A(n11588), .B(n11554), .Z(n11705) );
  XNOR U12025 ( .A(n11706), .B(n11707), .Z(n11554) );
  XOR U12026 ( .A(n11708), .B(n11604), .Z(n11707) );
  NANDN U12027 ( .A(n11709), .B(n11710), .Z(n11604) );
  NOR U12028 ( .A(n11711), .B(n11712), .Z(n11708) );
  XNOR U12029 ( .A(n11587), .B(n11557), .Z(n11704) );
  XNOR U12030 ( .A(n7231), .B(n6297), .Z(n7215) );
  XNOR U12031 ( .A(n11611), .B(n6262), .Z(n6297) );
  XOR U12032 ( .A(n11505), .B(n11713), .Z(n6262) );
  XOR U12033 ( .A(n11713), .B(n11611), .Z(n7231) );
  XNOR U12034 ( .A(n11612), .B(n11714), .Z(n11611) );
  XNOR U12035 ( .A(n11715), .B(n11716), .Z(n11714) );
  ANDN U12036 ( .B(n11552), .A(n11717), .Z(n11715) );
  XNOR U12037 ( .A(n11718), .B(n11719), .Z(n11612) );
  XNOR U12038 ( .A(n11720), .B(n11721), .Z(n11719) );
  NAND U12039 ( .A(n11722), .B(n11723), .Z(n11721) );
  XNOR U12040 ( .A(n11724), .B(n11725), .Z(n8539) );
  XNOR U12041 ( .A(n7218), .B(n8369), .Z(n11725) );
  XNOR U12042 ( .A(n11632), .B(n11540), .Z(n8369) );
  XOR U12043 ( .A(n11576), .B(n11726), .Z(n11540) );
  XNOR U12044 ( .A(n11727), .B(n11645), .Z(n11726) );
  NOR U12045 ( .A(n11639), .B(n11728), .Z(n11645) );
  XNOR U12046 ( .A(n11641), .B(n11648), .Z(n11639) );
  ANDN U12047 ( .B(n11641), .A(n11729), .Z(n11727) );
  XNOR U12048 ( .A(n11643), .B(n11730), .Z(n11576) );
  XNOR U12049 ( .A(n11731), .B(n11732), .Z(n11730) );
  NANDN U12050 ( .A(n11662), .B(n11733), .Z(n11732) );
  IV U12051 ( .A(n11591), .Z(n11632) );
  XNOR U12052 ( .A(n11643), .B(n11734), .Z(n11591) );
  XOR U12053 ( .A(n11735), .B(n11578), .Z(n11734) );
  OR U12054 ( .A(n11736), .B(n11657), .Z(n11578) );
  XNOR U12055 ( .A(n11581), .B(n11653), .Z(n11657) );
  ANDN U12056 ( .B(n11653), .A(n11737), .Z(n11735) );
  XOR U12057 ( .A(n11738), .B(n11731), .Z(n11643) );
  OR U12058 ( .A(n11665), .B(n11739), .Z(n11731) );
  XOR U12059 ( .A(n11667), .B(n11662), .Z(n11665) );
  XOR U12060 ( .A(n11653), .B(n11547), .Z(n11662) );
  IV U12061 ( .A(n11648), .Z(n11547) );
  XOR U12062 ( .A(n11740), .B(n11741), .Z(n11648) );
  NANDN U12063 ( .A(n11742), .B(n11743), .Z(n11741) );
  XOR U12064 ( .A(n11744), .B(n11745), .Z(n11653) );
  NANDN U12065 ( .A(n11742), .B(n11746), .Z(n11745) );
  AND U12066 ( .A(n11747), .B(n11667), .Z(n11738) );
  XOR U12067 ( .A(n11641), .B(n11581), .Z(n11667) );
  XNOR U12068 ( .A(n11748), .B(n11744), .Z(n11581) );
  NANDN U12069 ( .A(n11749), .B(n11750), .Z(n11744) );
  XOR U12070 ( .A(n11746), .B(n11751), .Z(n11750) );
  ANDN U12071 ( .B(n11751), .A(n11752), .Z(n11748) );
  NANDN U12072 ( .A(n11749), .B(n11754), .Z(n11740) );
  XOR U12073 ( .A(n11755), .B(n11743), .Z(n11754) );
  XNOR U12074 ( .A(n11756), .B(n11757), .Z(n11742) );
  XOR U12075 ( .A(n11758), .B(n11759), .Z(n11757) );
  XNOR U12076 ( .A(n11760), .B(n11761), .Z(n11756) );
  XNOR U12077 ( .A(n11762), .B(n11763), .Z(n11761) );
  ANDN U12078 ( .B(n11755), .A(n11759), .Z(n11762) );
  ANDN U12079 ( .B(n11755), .A(n11752), .Z(n11753) );
  XNOR U12080 ( .A(n11758), .B(n11764), .Z(n11752) );
  XOR U12081 ( .A(n11765), .B(n11763), .Z(n11764) );
  NAND U12082 ( .A(n11766), .B(n11767), .Z(n11763) );
  XNOR U12083 ( .A(n11760), .B(n11743), .Z(n11767) );
  IV U12084 ( .A(n11755), .Z(n11760) );
  XNOR U12085 ( .A(n11746), .B(n11759), .Z(n11766) );
  IV U12086 ( .A(n11751), .Z(n11759) );
  XOR U12087 ( .A(n11768), .B(n11769), .Z(n11751) );
  XNOR U12088 ( .A(n11770), .B(n11771), .Z(n11769) );
  XNOR U12089 ( .A(n11772), .B(n11773), .Z(n11768) );
  ANDN U12090 ( .B(n11774), .A(n11729), .Z(n11772) );
  AND U12091 ( .A(n11743), .B(n11746), .Z(n11765) );
  XNOR U12092 ( .A(n11743), .B(n11746), .Z(n11758) );
  XNOR U12093 ( .A(n11775), .B(n11776), .Z(n11746) );
  XNOR U12094 ( .A(n11777), .B(n11771), .Z(n11776) );
  XOR U12095 ( .A(n11778), .B(n11779), .Z(n11775) );
  XNOR U12096 ( .A(n11780), .B(n11773), .Z(n11779) );
  OR U12097 ( .A(n11640), .B(n11728), .Z(n11773) );
  XNOR U12098 ( .A(n11781), .B(n11812), .Z(n11728) );
  XNOR U12099 ( .A(n11642), .B(n11782), .Z(n11640) );
  ANDN U12100 ( .B(n11546), .A(n11647), .Z(n11780) );
  XNOR U12101 ( .A(n11783), .B(n11784), .Z(n11743) );
  XNOR U12102 ( .A(n11771), .B(n11785), .Z(n11784) );
  XNOR U12103 ( .A(n11656), .B(n11778), .Z(n11785) );
  XNOR U12104 ( .A(n11642), .B(n11781), .Z(n11771) );
  XNOR U12105 ( .A(n11786), .B(n11787), .Z(n11783) );
  XNOR U12106 ( .A(n11788), .B(n11789), .Z(n11787) );
  ANDN U12107 ( .B(n11790), .A(n11737), .Z(n11788) );
  XNOR U12108 ( .A(n11791), .B(n11792), .Z(n11755) );
  XNOR U12109 ( .A(n11777), .B(n11793), .Z(n11792) );
  XNOR U12110 ( .A(n11794), .B(n11770), .Z(n11793) );
  XOR U12111 ( .A(n11778), .B(n11795), .Z(n11770) );
  XNOR U12112 ( .A(n11796), .B(n11797), .Z(n11795) );
  NANDN U12113 ( .A(n11663), .B(n11733), .Z(n11797) );
  XNOR U12114 ( .A(n11798), .B(n11796), .Z(n11778) );
  OR U12115 ( .A(n11739), .B(n11666), .Z(n11796) );
  XOR U12116 ( .A(n11799), .B(n11663), .Z(n11666) );
  XNOR U12117 ( .A(n11546), .B(n11790), .Z(n11663) );
  IV U12118 ( .A(n11782), .Z(n11546) );
  XNOR U12119 ( .A(n11747), .B(n11733), .Z(n11739) );
  XNOR U12120 ( .A(n11737), .B(n11812), .Z(n11733) );
  IV U12121 ( .A(n11794), .Z(n11737) );
  ANDN U12122 ( .B(n11747), .A(n11668), .Z(n11798) );
  IV U12123 ( .A(n11799), .Z(n11668) );
  XOR U12124 ( .A(n11774), .B(n11656), .Z(n11799) );
  XOR U12125 ( .A(n11782), .B(n11647), .Z(n11777) );
  XOR U12126 ( .A(n11800), .B(n11801), .Z(n11647) );
  XOR U12127 ( .A(n11802), .B(n11803), .Z(n11782) );
  XOR U12128 ( .A(n11804), .B(n11801), .Z(n11803) );
  XNOR U12129 ( .A(n11652), .B(n11805), .Z(n11791) );
  XNOR U12130 ( .A(n11806), .B(n11789), .Z(n11805) );
  OR U12131 ( .A(n11658), .B(n11736), .Z(n11789) );
  XNOR U12132 ( .A(n11786), .B(n11794), .Z(n11736) );
  XOR U12133 ( .A(n11807), .B(n11808), .Z(n11794) );
  XNOR U12134 ( .A(n11809), .B(n11810), .Z(n11808) );
  XOR U12135 ( .A(n11786), .B(n11811), .Z(n11807) );
  XNOR U12136 ( .A(n11656), .B(n11790), .Z(n11658) );
  IV U12137 ( .A(n11652), .Z(n11790) );
  ANDN U12138 ( .B(n11656), .A(n11580), .Z(n11806) );
  XOR U12139 ( .A(n11809), .B(n11812), .Z(n11656) );
  XOR U12140 ( .A(n11813), .B(n11814), .Z(n11809) );
  XNOR U12141 ( .A(n9457), .B(n10355), .Z(n11814) );
  XOR U12142 ( .A(n10351), .B(n10954), .Z(n10355) );
  XOR U12143 ( .A(n10358), .B(n10946), .Z(n9457) );
  XOR U12144 ( .A(n11815), .B(n10329), .Z(n10358) );
  IV U12145 ( .A(n11816), .Z(n10329) );
  XNOR U12146 ( .A(n9456), .B(n11817), .Z(n11813) );
  XNOR U12147 ( .A(key[860]), .B(n10944), .Z(n11817) );
  XNOR U12148 ( .A(n10968), .B(n11818), .Z(n10944) );
  XNOR U12149 ( .A(n10373), .B(n9446), .Z(n9456) );
  XNOR U12150 ( .A(n11819), .B(n11820), .Z(n9446) );
  XNOR U12151 ( .A(n11821), .B(n11822), .Z(n11820) );
  XNOR U12152 ( .A(n11823), .B(n11824), .Z(n11819) );
  XOR U12153 ( .A(n11825), .B(n11826), .Z(n11824) );
  ANDN U12154 ( .B(n11827), .A(n11828), .Z(n11826) );
  XNOR U12155 ( .A(n11829), .B(n11830), .Z(n11652) );
  XOR U12156 ( .A(n11642), .B(n11802), .Z(n11830) );
  IV U12157 ( .A(n11774), .Z(n11642) );
  XOR U12158 ( .A(n11811), .B(n11812), .Z(n11774) );
  XNOR U12159 ( .A(n11800), .B(n11801), .Z(n11812) );
  IV U12160 ( .A(n11804), .Z(n11800) );
  XNOR U12161 ( .A(n11831), .B(n11832), .Z(n11804) );
  XOR U12162 ( .A(n10949), .B(n9445), .Z(n11832) );
  XOR U12163 ( .A(n10342), .B(n10954), .Z(n9445) );
  XNOR U12164 ( .A(n11833), .B(n11834), .Z(n10954) );
  XNOR U12165 ( .A(n11835), .B(n11836), .Z(n11834) );
  XNOR U12166 ( .A(n11837), .B(n11838), .Z(n11833) );
  XOR U12167 ( .A(n11839), .B(n11840), .Z(n11838) );
  ANDN U12168 ( .B(n11841), .A(n11842), .Z(n11840) );
  XNOR U12169 ( .A(n11843), .B(n11844), .Z(n10342) );
  XNOR U12170 ( .A(n11845), .B(n11846), .Z(n11844) );
  XNOR U12171 ( .A(n11815), .B(n11847), .Z(n11843) );
  XOR U12172 ( .A(n11848), .B(n11849), .Z(n11847) );
  ANDN U12173 ( .B(n11850), .A(n11851), .Z(n11849) );
  XOR U12174 ( .A(n11852), .B(n11853), .Z(n10949) );
  XOR U12175 ( .A(n11818), .B(n11854), .Z(n11853) );
  XNOR U12176 ( .A(n11855), .B(n11856), .Z(n11852) );
  XNOR U12177 ( .A(n11857), .B(n11858), .Z(n11856) );
  ANDN U12178 ( .B(n11859), .A(n11860), .Z(n11857) );
  XNOR U12179 ( .A(n10974), .B(n11861), .Z(n11831) );
  XOR U12180 ( .A(key[861]), .B(n10972), .Z(n11861) );
  IV U12181 ( .A(n9438), .Z(n10972) );
  XOR U12182 ( .A(n11862), .B(n11863), .Z(n9438) );
  XOR U12183 ( .A(n11864), .B(n11865), .Z(n11811) );
  XNOR U12184 ( .A(n10976), .B(n9452), .Z(n11865) );
  XNOR U12185 ( .A(n10971), .B(n10961), .Z(n9452) );
  XNOR U12186 ( .A(n11866), .B(n11867), .Z(n10971) );
  XNOR U12187 ( .A(n11868), .B(n11846), .Z(n11867) );
  XNOR U12188 ( .A(n11869), .B(n11870), .Z(n11846) );
  XNOR U12189 ( .A(n11871), .B(n11872), .Z(n11870) );
  NANDN U12190 ( .A(n11873), .B(n11874), .Z(n11872) );
  XNOR U12191 ( .A(n11875), .B(n11876), .Z(n11866) );
  XNOR U12192 ( .A(n11877), .B(n11878), .Z(n10976) );
  XOR U12193 ( .A(n11879), .B(n11854), .Z(n11878) );
  XNOR U12194 ( .A(n11880), .B(n11881), .Z(n11854) );
  XNOR U12195 ( .A(n11882), .B(n11883), .Z(n11881) );
  OR U12196 ( .A(n11884), .B(n11885), .Z(n11883) );
  XNOR U12197 ( .A(n11886), .B(n11887), .Z(n11877) );
  XOR U12198 ( .A(key[863]), .B(n9477), .Z(n11864) );
  XOR U12199 ( .A(n10373), .B(n10351), .Z(n9477) );
  XOR U12200 ( .A(n11580), .B(n11729), .Z(n11747) );
  IV U12201 ( .A(n11781), .Z(n11729) );
  XNOR U12202 ( .A(n11810), .B(n11888), .Z(n11781) );
  XNOR U12203 ( .A(n11801), .B(n11829), .Z(n11888) );
  XOR U12204 ( .A(n11889), .B(n11890), .Z(n11829) );
  XOR U12205 ( .A(n11816), .B(n10966), .Z(n9430) );
  XNOR U12206 ( .A(n11891), .B(n11876), .Z(n11816) );
  XOR U12207 ( .A(n11892), .B(n11887), .Z(n10968) );
  XNOR U12208 ( .A(n10989), .B(n11893), .Z(n11889) );
  XOR U12209 ( .A(key[858]), .B(n10981), .Z(n11893) );
  XNOR U12210 ( .A(n11894), .B(n11895), .Z(n10981) );
  XOR U12211 ( .A(n11896), .B(n11863), .Z(n11895) );
  XNOR U12212 ( .A(n11897), .B(n11898), .Z(n11863) );
  XNOR U12213 ( .A(n11899), .B(n11825), .Z(n11898) );
  NOR U12214 ( .A(n11900), .B(n11901), .Z(n11825) );
  NOR U12215 ( .A(n11902), .B(n11903), .Z(n11899) );
  XNOR U12216 ( .A(n11904), .B(n11905), .Z(n11894) );
  XOR U12217 ( .A(n11906), .B(n11907), .Z(n11801) );
  XOR U12218 ( .A(n10337), .B(n11580), .Z(n11907) );
  XOR U12219 ( .A(n11908), .B(n11909), .Z(n10961) );
  XOR U12220 ( .A(n11910), .B(n11836), .Z(n11909) );
  XNOR U12221 ( .A(n11911), .B(n11912), .Z(n11836) );
  XNOR U12222 ( .A(n11913), .B(n11914), .Z(n11912) );
  OR U12223 ( .A(n11915), .B(n11916), .Z(n11914) );
  XNOR U12224 ( .A(n11917), .B(n11918), .Z(n11908) );
  XOR U12225 ( .A(n10973), .B(n11919), .Z(n11906) );
  XOR U12226 ( .A(key[862]), .B(n9439), .Z(n11919) );
  XOR U12227 ( .A(n10344), .B(n9451), .Z(n9439) );
  XNOR U12228 ( .A(n10373), .B(n10960), .Z(n9451) );
  XNOR U12229 ( .A(n11920), .B(n11921), .Z(n10960) );
  XOR U12230 ( .A(n11896), .B(n11822), .Z(n11921) );
  XNOR U12231 ( .A(n11922), .B(n11923), .Z(n11822) );
  XNOR U12232 ( .A(n11924), .B(n11925), .Z(n11923) );
  NANDN U12233 ( .A(n11926), .B(n11927), .Z(n11925) );
  XOR U12234 ( .A(n11904), .B(n11862), .Z(n11920) );
  XNOR U12235 ( .A(n10339), .B(n10974), .Z(n10344) );
  XOR U12236 ( .A(n11928), .B(n11929), .Z(n10974) );
  XNOR U12237 ( .A(n11930), .B(n11931), .Z(n10339) );
  XOR U12238 ( .A(n11891), .B(n11932), .Z(n11931) );
  XOR U12239 ( .A(n11933), .B(n11934), .Z(n10973) );
  XNOR U12240 ( .A(n11892), .B(n11935), .Z(n11934) );
  XOR U12241 ( .A(n11936), .B(n11937), .Z(n11810) );
  XOR U12242 ( .A(n11802), .B(n11938), .Z(n11937) );
  XNOR U12243 ( .A(n10980), .B(n10361), .Z(n11938) );
  XOR U12244 ( .A(n10351), .B(n10946), .Z(n10361) );
  XNOR U12245 ( .A(n11837), .B(n10966), .Z(n10946) );
  XNOR U12246 ( .A(n11939), .B(n11940), .Z(n10980) );
  XOR U12247 ( .A(n11879), .B(n11933), .Z(n11940) );
  XNOR U12248 ( .A(n11941), .B(n11942), .Z(n11933) );
  XNOR U12249 ( .A(n11858), .B(n11943), .Z(n11942) );
  OR U12250 ( .A(n11944), .B(n11945), .Z(n11943) );
  NANDN U12251 ( .A(n11946), .B(n11947), .Z(n11858) );
  XOR U12252 ( .A(n11935), .B(n11887), .Z(n11939) );
  XNOR U12253 ( .A(n11948), .B(n11949), .Z(n11802) );
  XOR U12254 ( .A(n9431), .B(n10966), .Z(n11949) );
  XOR U12255 ( .A(n11950), .B(n11951), .Z(n10966) );
  XNOR U12256 ( .A(n9468), .B(n11952), .Z(n11948) );
  XOR U12257 ( .A(key[857]), .B(n10987), .Z(n11952) );
  XNOR U12258 ( .A(n11879), .B(n11953), .Z(n10987) );
  XOR U12259 ( .A(n11886), .B(n11887), .Z(n11953) );
  XOR U12260 ( .A(n11954), .B(n11955), .Z(n11887) );
  XNOR U12261 ( .A(n11956), .B(n11957), .Z(n11955) );
  NAND U12262 ( .A(n11958), .B(n11859), .Z(n11957) );
  XOR U12263 ( .A(n11959), .B(n11935), .Z(n11886) );
  XOR U12264 ( .A(n11855), .B(n11960), .Z(n11935) );
  XOR U12265 ( .A(n11961), .B(n11962), .Z(n11960) );
  AND U12266 ( .A(n11963), .B(n11964), .Z(n11961) );
  XOR U12267 ( .A(n11941), .B(n11965), .Z(n11879) );
  XNOR U12268 ( .A(n11962), .B(n11966), .Z(n11965) );
  OR U12269 ( .A(n11884), .B(n11967), .Z(n11966) );
  OR U12270 ( .A(n11968), .B(n11969), .Z(n11962) );
  XNOR U12271 ( .A(n11855), .B(n11970), .Z(n11941) );
  XNOR U12272 ( .A(n11971), .B(n11972), .Z(n11970) );
  NAND U12273 ( .A(n11973), .B(n11974), .Z(n11972) );
  XOR U12274 ( .A(n11975), .B(n11971), .Z(n11855) );
  NANDN U12275 ( .A(n11976), .B(n11977), .Z(n11971) );
  AND U12276 ( .A(n11978), .B(n11979), .Z(n11975) );
  XOR U12277 ( .A(n10984), .B(n10366), .Z(n9468) );
  XOR U12278 ( .A(n11868), .B(n11980), .Z(n10366) );
  XNOR U12279 ( .A(n11875), .B(n11981), .Z(n11980) );
  XNOR U12280 ( .A(n11982), .B(n11932), .Z(n11868) );
  XNOR U12281 ( .A(n9463), .B(n11983), .Z(n11936) );
  XNOR U12282 ( .A(key[859]), .B(n9471), .Z(n11983) );
  XOR U12283 ( .A(n10989), .B(n10369), .Z(n9471) );
  XNOR U12284 ( .A(n11984), .B(n11985), .Z(n10369) );
  XNOR U12285 ( .A(n11876), .B(n11930), .Z(n11985) );
  XNOR U12286 ( .A(n11986), .B(n11987), .Z(n11930) );
  XNOR U12287 ( .A(n11988), .B(n11848), .Z(n11987) );
  NOR U12288 ( .A(n11989), .B(n11990), .Z(n11848) );
  ANDN U12289 ( .B(n11991), .A(n11992), .Z(n11988) );
  IV U12290 ( .A(n11981), .Z(n11876) );
  XNOR U12291 ( .A(n11994), .B(n11995), .Z(n11993) );
  NANDN U12292 ( .A(n11851), .B(n11996), .Z(n11995) );
  XNOR U12293 ( .A(n11875), .B(n11932), .Z(n11984) );
  XNOR U12294 ( .A(n11845), .B(n11998), .Z(n11932) );
  XNOR U12295 ( .A(n11999), .B(n12000), .Z(n11998) );
  NANDN U12296 ( .A(n12001), .B(n12002), .Z(n12000) );
  XOR U12297 ( .A(n12004), .B(n11999), .Z(n12003) );
  OR U12298 ( .A(n12005), .B(n12006), .Z(n11999) );
  AND U12299 ( .A(n11874), .B(n12007), .Z(n12004) );
  XNOR U12300 ( .A(n11845), .B(n12008), .Z(n11986) );
  XNOR U12301 ( .A(n12009), .B(n12010), .Z(n12008) );
  NAND U12302 ( .A(n12011), .B(n12012), .Z(n12010) );
  XOR U12303 ( .A(n12013), .B(n12009), .Z(n11845) );
  NANDN U12304 ( .A(n12014), .B(n12015), .Z(n12009) );
  ANDN U12305 ( .B(n12016), .A(n12017), .Z(n12013) );
  XOR U12306 ( .A(n12018), .B(n12019), .Z(n10989) );
  XOR U12307 ( .A(n11918), .B(n11928), .Z(n12019) );
  XNOR U12308 ( .A(n12020), .B(n12021), .Z(n11928) );
  XNOR U12309 ( .A(n12022), .B(n11839), .Z(n12021) );
  ANDN U12310 ( .B(n12023), .A(n12024), .Z(n11839) );
  ANDN U12311 ( .B(n12025), .A(n12026), .Z(n12022) );
  IV U12312 ( .A(n11951), .Z(n11918) );
  XOR U12313 ( .A(n11917), .B(n12027), .Z(n12018) );
  XNOR U12314 ( .A(n10373), .B(n10945), .Z(n9463) );
  XOR U12315 ( .A(n11821), .B(n9431), .Z(n10945) );
  XOR U12316 ( .A(n12028), .B(n11896), .Z(n9431) );
  XOR U12317 ( .A(n12028), .B(n11821), .Z(n10373) );
  XNOR U12318 ( .A(n11922), .B(n12029), .Z(n11821) );
  XOR U12319 ( .A(n12030), .B(n12031), .Z(n12029) );
  ANDN U12320 ( .B(n12032), .A(n11903), .Z(n12030) );
  XNOR U12321 ( .A(n12033), .B(n12034), .Z(n11922) );
  XNOR U12322 ( .A(n12035), .B(n12036), .Z(n12034) );
  NANDN U12323 ( .A(n12037), .B(n12038), .Z(n12036) );
  IV U12324 ( .A(n11786), .Z(n11580) );
  XOR U12325 ( .A(n12039), .B(n12040), .Z(n11786) );
  XNOR U12326 ( .A(n10984), .B(n10372), .Z(n12040) );
  XNOR U12327 ( .A(n9478), .B(n9453), .Z(n10372) );
  IV U12328 ( .A(n10948), .Z(n9453) );
  XOR U12329 ( .A(n11892), .B(n11818), .Z(n10948) );
  XOR U12330 ( .A(n11880), .B(n12041), .Z(n11818) );
  XOR U12331 ( .A(n12042), .B(n11956), .Z(n12041) );
  NANDN U12332 ( .A(n12043), .B(n11947), .Z(n11956) );
  XNOR U12333 ( .A(n11944), .B(n11859), .Z(n11947) );
  NOR U12334 ( .A(n12044), .B(n11944), .Z(n12042) );
  XNOR U12335 ( .A(n11954), .B(n12045), .Z(n11880) );
  XNOR U12336 ( .A(n12046), .B(n12047), .Z(n12045) );
  NAND U12337 ( .A(n11974), .B(n12048), .Z(n12047) );
  IV U12338 ( .A(n11959), .Z(n11892) );
  XNOR U12339 ( .A(n11954), .B(n12049), .Z(n11959) );
  XOR U12340 ( .A(n12050), .B(n11882), .Z(n12049) );
  OR U12341 ( .A(n11969), .B(n12051), .Z(n11882) );
  XOR U12342 ( .A(n11884), .B(n11964), .Z(n11969) );
  ANDN U12343 ( .B(n11964), .A(n12052), .Z(n12050) );
  XOR U12344 ( .A(n12053), .B(n12046), .Z(n11954) );
  OR U12345 ( .A(n11976), .B(n12054), .Z(n12046) );
  XNOR U12346 ( .A(n11978), .B(n11974), .Z(n11976) );
  XOR U12347 ( .A(n11964), .B(n11859), .Z(n11974) );
  XOR U12348 ( .A(n12055), .B(n12056), .Z(n11859) );
  NANDN U12349 ( .A(n12057), .B(n12058), .Z(n12056) );
  XOR U12350 ( .A(n12059), .B(n12060), .Z(n11964) );
  OR U12351 ( .A(n12057), .B(n12061), .Z(n12060) );
  ANDN U12352 ( .B(n11978), .A(n12062), .Z(n12053) );
  XOR U12353 ( .A(n11884), .B(n11944), .Z(n11978) );
  XOR U12354 ( .A(n12063), .B(n12055), .Z(n11944) );
  NANDN U12355 ( .A(n12064), .B(n12065), .Z(n12055) );
  ANDN U12356 ( .B(n12066), .A(n12067), .Z(n12063) );
  NANDN U12357 ( .A(n12064), .B(n12069), .Z(n12059) );
  XOR U12358 ( .A(n12070), .B(n12057), .Z(n12064) );
  XNOR U12359 ( .A(n12071), .B(n12072), .Z(n12057) );
  XOR U12360 ( .A(n12073), .B(n12066), .Z(n12072) );
  XNOR U12361 ( .A(n12074), .B(n12075), .Z(n12071) );
  XNOR U12362 ( .A(n12076), .B(n12077), .Z(n12075) );
  ANDN U12363 ( .B(n12066), .A(n12078), .Z(n12076) );
  IV U12364 ( .A(n12079), .Z(n12066) );
  ANDN U12365 ( .B(n12070), .A(n12078), .Z(n12068) );
  IV U12366 ( .A(n12074), .Z(n12078) );
  IV U12367 ( .A(n12067), .Z(n12070) );
  XNOR U12368 ( .A(n12073), .B(n12080), .Z(n12067) );
  XOR U12369 ( .A(n12081), .B(n12077), .Z(n12080) );
  NAND U12370 ( .A(n12069), .B(n12065), .Z(n12077) );
  XNOR U12371 ( .A(n12058), .B(n12079), .Z(n12065) );
  XOR U12372 ( .A(n12082), .B(n12083), .Z(n12079) );
  XOR U12373 ( .A(n12084), .B(n12085), .Z(n12083) );
  XNOR U12374 ( .A(n11963), .B(n12086), .Z(n12085) );
  XNOR U12375 ( .A(n12087), .B(n12088), .Z(n12082) );
  XNOR U12376 ( .A(n12089), .B(n12090), .Z(n12088) );
  ANDN U12377 ( .B(n12091), .A(n11885), .Z(n12089) );
  XNOR U12378 ( .A(n12074), .B(n12061), .Z(n12069) );
  XOR U12379 ( .A(n12092), .B(n12093), .Z(n12074) );
  XNOR U12380 ( .A(n12094), .B(n12086), .Z(n12093) );
  XOR U12381 ( .A(n12095), .B(n12096), .Z(n12086) );
  XNOR U12382 ( .A(n12097), .B(n12098), .Z(n12096) );
  NAND U12383 ( .A(n12048), .B(n11973), .Z(n12098) );
  XNOR U12384 ( .A(n12099), .B(n12100), .Z(n12092) );
  ANDN U12385 ( .B(n12101), .A(n12044), .Z(n12099) );
  ANDN U12386 ( .B(n12058), .A(n12061), .Z(n12081) );
  XOR U12387 ( .A(n12061), .B(n12058), .Z(n12073) );
  XNOR U12388 ( .A(n12102), .B(n12103), .Z(n12058) );
  XNOR U12389 ( .A(n12095), .B(n12104), .Z(n12103) );
  XOR U12390 ( .A(n12094), .B(n11967), .Z(n12104) );
  XOR U12391 ( .A(n11885), .B(n12105), .Z(n12102) );
  XNOR U12392 ( .A(n12106), .B(n12090), .Z(n12105) );
  OR U12393 ( .A(n11968), .B(n12051), .Z(n12090) );
  XNOR U12394 ( .A(n11885), .B(n12052), .Z(n12051) );
  XOR U12395 ( .A(n11967), .B(n11963), .Z(n11968) );
  ANDN U12396 ( .B(n11963), .A(n12052), .Z(n12106) );
  XOR U12397 ( .A(n12107), .B(n12108), .Z(n12061) );
  XOR U12398 ( .A(n12095), .B(n12084), .Z(n12108) );
  XOR U12399 ( .A(n11958), .B(n11860), .Z(n12084) );
  XOR U12400 ( .A(n12109), .B(n12097), .Z(n12095) );
  NANDN U12401 ( .A(n12054), .B(n11977), .Z(n12097) );
  XOR U12402 ( .A(n11979), .B(n11973), .Z(n11977) );
  XNOR U12403 ( .A(n12101), .B(n12110), .Z(n11963) );
  XOR U12404 ( .A(n12111), .B(n12112), .Z(n12110) );
  XOR U12405 ( .A(n12062), .B(n12048), .Z(n12054) );
  XNOR U12406 ( .A(n12052), .B(n11958), .Z(n12048) );
  IV U12407 ( .A(n12087), .Z(n12052) );
  XOR U12408 ( .A(n12113), .B(n12114), .Z(n12087) );
  XOR U12409 ( .A(n12115), .B(n12116), .Z(n12114) );
  XNOR U12410 ( .A(n11885), .B(n12117), .Z(n12113) );
  ANDN U12411 ( .B(n11979), .A(n12062), .Z(n12109) );
  XNOR U12412 ( .A(n11885), .B(n12044), .Z(n12062) );
  XOR U12413 ( .A(n12101), .B(n12091), .Z(n11979) );
  IV U12414 ( .A(n11967), .Z(n12091) );
  XOR U12415 ( .A(n12118), .B(n12119), .Z(n11967) );
  XOR U12416 ( .A(n12120), .B(n12116), .Z(n12119) );
  XNOR U12417 ( .A(n12121), .B(n12122), .Z(n12116) );
  XNOR U12418 ( .A(n12123), .B(n12124), .Z(n12122) );
  XOR U12419 ( .A(n12125), .B(n12126), .Z(n12121) );
  XNOR U12420 ( .A(key[740]), .B(n12127), .Z(n12126) );
  IV U12421 ( .A(n11945), .Z(n12101) );
  XOR U12422 ( .A(n12094), .B(n12128), .Z(n12107) );
  XNOR U12423 ( .A(n12129), .B(n12100), .Z(n12128) );
  OR U12424 ( .A(n11946), .B(n12043), .Z(n12100) );
  XNOR U12425 ( .A(n12130), .B(n11958), .Z(n12043) );
  XNOR U12426 ( .A(n11945), .B(n11860), .Z(n11946) );
  ANDN U12427 ( .B(n11958), .A(n11860), .Z(n12129) );
  XOR U12428 ( .A(n12118), .B(n12131), .Z(n11860) );
  XNOR U12429 ( .A(n12112), .B(n12132), .Z(n12131) );
  XOR U12430 ( .A(n12120), .B(n12118), .Z(n11958) );
  XNOR U12431 ( .A(n12044), .B(n11945), .Z(n12094) );
  XOR U12432 ( .A(n12118), .B(n12133), .Z(n11945) );
  XNOR U12433 ( .A(n12120), .B(n12115), .Z(n12133) );
  XOR U12434 ( .A(n12134), .B(n12135), .Z(n12115) );
  XNOR U12435 ( .A(n12136), .B(n12137), .Z(n12135) );
  XNOR U12436 ( .A(key[743]), .B(n12138), .Z(n12134) );
  XNOR U12437 ( .A(n12139), .B(n12140), .Z(n12118) );
  XOR U12438 ( .A(n12141), .B(n12142), .Z(n12140) );
  XNOR U12439 ( .A(key[741]), .B(n12143), .Z(n12139) );
  IV U12440 ( .A(n12130), .Z(n12044) );
  XOR U12441 ( .A(n12132), .B(n12144), .Z(n12130) );
  XNOR U12442 ( .A(n12111), .B(n12117), .Z(n12144) );
  XOR U12443 ( .A(n12145), .B(n12146), .Z(n12117) );
  XNOR U12444 ( .A(n12147), .B(n12148), .Z(n12146) );
  XOR U12445 ( .A(n12112), .B(n12149), .Z(n12148) );
  XNOR U12446 ( .A(n12150), .B(n12151), .Z(n12112) );
  XNOR U12447 ( .A(n12152), .B(n12153), .Z(n12151) );
  XOR U12448 ( .A(key[737]), .B(n12154), .Z(n12150) );
  XNOR U12449 ( .A(n12155), .B(n12156), .Z(n12145) );
  XOR U12450 ( .A(key[739]), .B(n12157), .Z(n12156) );
  XOR U12451 ( .A(n12158), .B(n12159), .Z(n12111) );
  XNOR U12452 ( .A(n12160), .B(n12161), .Z(n12159) );
  XNOR U12453 ( .A(key[738]), .B(n12162), .Z(n12158) );
  IV U12454 ( .A(n12120), .Z(n12132) );
  XOR U12455 ( .A(n12163), .B(n12164), .Z(n12120) );
  XOR U12456 ( .A(n11885), .B(n12165), .Z(n12164) );
  XNOR U12457 ( .A(n12166), .B(n12167), .Z(n11885) );
  XOR U12458 ( .A(n12168), .B(n12169), .Z(n12167) );
  XOR U12459 ( .A(key[736]), .B(n12170), .Z(n12166) );
  XNOR U12460 ( .A(n12171), .B(n12172), .Z(n12163) );
  XNOR U12461 ( .A(key[742]), .B(n12173), .Z(n12172) );
  XOR U12462 ( .A(n11891), .B(n11815), .Z(n9478) );
  XNOR U12463 ( .A(n11869), .B(n12174), .Z(n11815) );
  XNOR U12464 ( .A(n11994), .B(n12175), .Z(n12174) );
  NANDN U12465 ( .A(n12176), .B(n11991), .Z(n12175) );
  OR U12466 ( .A(n12177), .B(n11989), .Z(n11994) );
  XNOR U12467 ( .A(n11991), .B(n12178), .Z(n11989) );
  XOR U12468 ( .A(n11997), .B(n12179), .Z(n11869) );
  XNOR U12469 ( .A(n12180), .B(n12181), .Z(n12179) );
  NAND U12470 ( .A(n12012), .B(n12182), .Z(n12181) );
  IV U12471 ( .A(n11982), .Z(n11891) );
  XOR U12472 ( .A(n11997), .B(n12183), .Z(n11982) );
  XOR U12473 ( .A(n12184), .B(n11871), .Z(n12183) );
  OR U12474 ( .A(n12185), .B(n12005), .Z(n11871) );
  XOR U12475 ( .A(n11874), .B(n12001), .Z(n12005) );
  NOR U12476 ( .A(n12186), .B(n12001), .Z(n12184) );
  XNOR U12477 ( .A(n12187), .B(n12180), .Z(n11997) );
  OR U12478 ( .A(n12188), .B(n12014), .Z(n12180) );
  XOR U12479 ( .A(n12017), .B(n12012), .Z(n12014) );
  XOR U12480 ( .A(n12001), .B(n11851), .Z(n12012) );
  IV U12481 ( .A(n12178), .Z(n11851) );
  XOR U12482 ( .A(n12189), .B(n12190), .Z(n12178) );
  NANDN U12483 ( .A(n12191), .B(n12192), .Z(n12190) );
  XNOR U12484 ( .A(n12193), .B(n12194), .Z(n12001) );
  OR U12485 ( .A(n12191), .B(n12195), .Z(n12194) );
  ANDN U12486 ( .B(n12196), .A(n12017), .Z(n12187) );
  XNOR U12487 ( .A(n11874), .B(n11991), .Z(n12017) );
  XOR U12488 ( .A(n12189), .B(n12197), .Z(n11991) );
  NANDN U12489 ( .A(n12198), .B(n12199), .Z(n12197) );
  NANDN U12490 ( .A(n12200), .B(n12201), .Z(n12189) );
  OR U12491 ( .A(n12203), .B(n12200), .Z(n12193) );
  XOR U12492 ( .A(n12204), .B(n12191), .Z(n12200) );
  XNOR U12493 ( .A(n12205), .B(n12206), .Z(n12191) );
  XOR U12494 ( .A(n12207), .B(n12199), .Z(n12206) );
  XNOR U12495 ( .A(n12208), .B(n12209), .Z(n12205) );
  XNOR U12496 ( .A(n12210), .B(n12211), .Z(n12209) );
  ANDN U12497 ( .B(n12199), .A(n12212), .Z(n12210) );
  IV U12498 ( .A(n12213), .Z(n12199) );
  ANDN U12499 ( .B(n12204), .A(n12212), .Z(n12202) );
  IV U12500 ( .A(n12198), .Z(n12204) );
  XNOR U12501 ( .A(n12207), .B(n12214), .Z(n12198) );
  XNOR U12502 ( .A(n12211), .B(n12215), .Z(n12214) );
  NANDN U12503 ( .A(n12195), .B(n12192), .Z(n12215) );
  NANDN U12504 ( .A(n12203), .B(n12201), .Z(n12211) );
  XNOR U12505 ( .A(n12192), .B(n12213), .Z(n12201) );
  XOR U12506 ( .A(n12216), .B(n12217), .Z(n12213) );
  XOR U12507 ( .A(n12218), .B(n12219), .Z(n12217) );
  XNOR U12508 ( .A(n12002), .B(n12220), .Z(n12219) );
  XNOR U12509 ( .A(n12221), .B(n12222), .Z(n12216) );
  XNOR U12510 ( .A(n12223), .B(n12224), .Z(n12222) );
  ANDN U12511 ( .B(n12007), .A(n11873), .Z(n12223) );
  XNOR U12512 ( .A(n12212), .B(n12195), .Z(n12203) );
  IV U12513 ( .A(n12208), .Z(n12212) );
  XOR U12514 ( .A(n12225), .B(n12226), .Z(n12208) );
  XNOR U12515 ( .A(n12227), .B(n12220), .Z(n12226) );
  XOR U12516 ( .A(n12228), .B(n12229), .Z(n12220) );
  XNOR U12517 ( .A(n12230), .B(n12231), .Z(n12229) );
  NAND U12518 ( .A(n12182), .B(n12011), .Z(n12231) );
  XNOR U12519 ( .A(n12232), .B(n12233), .Z(n12225) );
  ANDN U12520 ( .B(n12234), .A(n12176), .Z(n12232) );
  XOR U12521 ( .A(n12195), .B(n12192), .Z(n12207) );
  XNOR U12522 ( .A(n12235), .B(n12236), .Z(n12192) );
  XNOR U12523 ( .A(n12228), .B(n12237), .Z(n12236) );
  XNOR U12524 ( .A(n12227), .B(n12007), .Z(n12237) );
  XNOR U12525 ( .A(n12238), .B(n12239), .Z(n12235) );
  XNOR U12526 ( .A(n12240), .B(n12224), .Z(n12239) );
  OR U12527 ( .A(n12006), .B(n12185), .Z(n12224) );
  XNOR U12528 ( .A(n12238), .B(n12221), .Z(n12185) );
  XNOR U12529 ( .A(n12007), .B(n12002), .Z(n12006) );
  ANDN U12530 ( .B(n12002), .A(n12186), .Z(n12240) );
  XOR U12531 ( .A(n12241), .B(n12242), .Z(n12195) );
  XOR U12532 ( .A(n12228), .B(n12218), .Z(n12242) );
  XNOR U12533 ( .A(n11996), .B(n11850), .Z(n12218) );
  XOR U12534 ( .A(n12243), .B(n12230), .Z(n12228) );
  NANDN U12535 ( .A(n12188), .B(n12015), .Z(n12230) );
  XOR U12536 ( .A(n12016), .B(n12011), .Z(n12015) );
  XOR U12537 ( .A(n11850), .B(n12002), .Z(n12011) );
  XNOR U12538 ( .A(n12234), .B(n12244), .Z(n12002) );
  XOR U12539 ( .A(n12245), .B(n12246), .Z(n12244) );
  XNOR U12540 ( .A(n12196), .B(n12182), .Z(n12188) );
  XNOR U12541 ( .A(n12186), .B(n11996), .Z(n12182) );
  IV U12542 ( .A(n12221), .Z(n12186) );
  XOR U12543 ( .A(n12247), .B(n12248), .Z(n12221) );
  XOR U12544 ( .A(n12249), .B(n12250), .Z(n12248) );
  XOR U12545 ( .A(n12238), .B(n12251), .Z(n12247) );
  AND U12546 ( .A(n12016), .B(n12196), .Z(n12243) );
  XOR U12547 ( .A(n12234), .B(n12007), .Z(n12016) );
  XNOR U12548 ( .A(n12252), .B(n12253), .Z(n12007) );
  XOR U12549 ( .A(n12254), .B(n12250), .Z(n12253) );
  XNOR U12550 ( .A(n12255), .B(n12256), .Z(n12250) );
  XNOR U12551 ( .A(n12257), .B(n12258), .Z(n12256) );
  XOR U12552 ( .A(key[652]), .B(n12259), .Z(n12255) );
  XOR U12553 ( .A(n12227), .B(n12260), .Z(n12241) );
  XNOR U12554 ( .A(n12261), .B(n12233), .Z(n12260) );
  OR U12555 ( .A(n11990), .B(n12177), .Z(n12233) );
  XNOR U12556 ( .A(n12262), .B(n11996), .Z(n12177) );
  XNOR U12557 ( .A(n12234), .B(n11850), .Z(n11990) );
  IV U12558 ( .A(n11992), .Z(n12234) );
  AND U12559 ( .A(n11850), .B(n11996), .Z(n12261) );
  XOR U12560 ( .A(n12254), .B(n12252), .Z(n11996) );
  XNOR U12561 ( .A(n12252), .B(n12263), .Z(n11850) );
  XNOR U12562 ( .A(n12264), .B(n12254), .Z(n12263) );
  XNOR U12563 ( .A(n12176), .B(n11992), .Z(n12227) );
  XOR U12564 ( .A(n12252), .B(n12265), .Z(n11992) );
  XNOR U12565 ( .A(n12254), .B(n12249), .Z(n12265) );
  XOR U12566 ( .A(n12266), .B(n12267), .Z(n12249) );
  XOR U12567 ( .A(n12268), .B(n12269), .Z(n12267) );
  XOR U12568 ( .A(key[655]), .B(n12270), .Z(n12266) );
  XNOR U12569 ( .A(n12271), .B(n12272), .Z(n12252) );
  XNOR U12570 ( .A(n12273), .B(n12274), .Z(n12272) );
  XNOR U12571 ( .A(n12275), .B(n12276), .Z(n12271) );
  XNOR U12572 ( .A(key[653]), .B(n12277), .Z(n12276) );
  XOR U12573 ( .A(n11873), .B(n12176), .Z(n12196) );
  IV U12574 ( .A(n12262), .Z(n12176) );
  XNOR U12575 ( .A(n12245), .B(n12251), .Z(n12278) );
  XOR U12576 ( .A(n12279), .B(n12280), .Z(n12251) );
  XNOR U12577 ( .A(n12281), .B(n12282), .Z(n12280) );
  XNOR U12578 ( .A(n12283), .B(n12246), .Z(n12282) );
  IV U12579 ( .A(n12264), .Z(n12246) );
  XOR U12580 ( .A(n12284), .B(n12285), .Z(n12264) );
  XNOR U12581 ( .A(n12286), .B(n12287), .Z(n12285) );
  XNOR U12582 ( .A(n12288), .B(n12289), .Z(n12284) );
  XNOR U12583 ( .A(key[649]), .B(n12290), .Z(n12289) );
  XNOR U12584 ( .A(n12291), .B(n12292), .Z(n12279) );
  XNOR U12585 ( .A(key[651]), .B(n12293), .Z(n12292) );
  XOR U12586 ( .A(n12294), .B(n12295), .Z(n12245) );
  XOR U12587 ( .A(n12296), .B(n12297), .Z(n12295) );
  XNOR U12588 ( .A(n12298), .B(n12299), .Z(n12294) );
  XNOR U12589 ( .A(key[650]), .B(n12300), .Z(n12299) );
  XOR U12590 ( .A(n12301), .B(n12302), .Z(n12254) );
  XNOR U12591 ( .A(n12238), .B(n12303), .Z(n12302) );
  XNOR U12592 ( .A(n12304), .B(n12305), .Z(n12301) );
  XNOR U12593 ( .A(key[654]), .B(n12306), .Z(n12305) );
  IV U12594 ( .A(n12238), .Z(n11873) );
  XOR U12595 ( .A(n12307), .B(n12308), .Z(n12238) );
  XOR U12596 ( .A(n12309), .B(n12310), .Z(n12308) );
  XOR U12597 ( .A(n12311), .B(n12312), .Z(n12307) );
  XNOR U12598 ( .A(key[648]), .B(n12313), .Z(n12312) );
  XOR U12599 ( .A(n11910), .B(n12314), .Z(n10984) );
  XNOR U12600 ( .A(n11917), .B(n11951), .Z(n12314) );
  XOR U12601 ( .A(n12315), .B(n12316), .Z(n11951) );
  XOR U12602 ( .A(n12317), .B(n12318), .Z(n12316) );
  NAND U12603 ( .A(n12319), .B(n11841), .Z(n12318) );
  XNOR U12604 ( .A(n12020), .B(n12320), .Z(n11917) );
  XNOR U12605 ( .A(n12321), .B(n12322), .Z(n12320) );
  OR U12606 ( .A(n11915), .B(n12323), .Z(n12322) );
  XOR U12607 ( .A(n11835), .B(n12324), .Z(n12020) );
  XNOR U12608 ( .A(n12325), .B(n12326), .Z(n12324) );
  NAND U12609 ( .A(n12327), .B(n12328), .Z(n12326) );
  IV U12610 ( .A(n11929), .Z(n11910) );
  XNOR U12611 ( .A(n11950), .B(n12027), .Z(n11929) );
  XOR U12612 ( .A(n11835), .B(n12329), .Z(n12027) );
  XNOR U12613 ( .A(n12321), .B(n12330), .Z(n12329) );
  NANDN U12614 ( .A(n12331), .B(n12332), .Z(n12330) );
  OR U12615 ( .A(n12333), .B(n12334), .Z(n12321) );
  XOR U12616 ( .A(n12335), .B(n12325), .Z(n11835) );
  NANDN U12617 ( .A(n12336), .B(n12337), .Z(n12325) );
  ANDN U12618 ( .B(n12338), .A(n12339), .Z(n12335) );
  XOR U12619 ( .A(n10351), .B(n12340), .Z(n12039) );
  XOR U12620 ( .A(key[856]), .B(n10986), .Z(n12340) );
  IV U12621 ( .A(n9470), .Z(n10986) );
  XOR U12622 ( .A(n11896), .B(n12341), .Z(n9470) );
  XNOR U12623 ( .A(n11904), .B(n11862), .Z(n12341) );
  XOR U12624 ( .A(n12028), .B(n11905), .Z(n11862) );
  XNOR U12625 ( .A(n11823), .B(n12342), .Z(n11905) );
  XNOR U12626 ( .A(n12343), .B(n12344), .Z(n12342) );
  NANDN U12627 ( .A(n12345), .B(n12346), .Z(n12344) );
  XNOR U12628 ( .A(n12033), .B(n12347), .Z(n12028) );
  XOR U12629 ( .A(n12348), .B(n11924), .Z(n12347) );
  OR U12630 ( .A(n12349), .B(n12350), .Z(n11924) );
  ANDN U12631 ( .B(n12346), .A(n12351), .Z(n12348) );
  XNOR U12632 ( .A(n12343), .B(n12353), .Z(n12352) );
  NAND U12633 ( .A(n12354), .B(n11927), .Z(n12353) );
  OR U12634 ( .A(n12349), .B(n12355), .Z(n12343) );
  XNOR U12635 ( .A(n11927), .B(n12346), .Z(n12349) );
  XNOR U12636 ( .A(n11823), .B(n12356), .Z(n11897) );
  XNOR U12637 ( .A(n12357), .B(n12358), .Z(n12356) );
  NANDN U12638 ( .A(n12359), .B(n12360), .Z(n12358) );
  XOR U12639 ( .A(n12361), .B(n12357), .Z(n11823) );
  OR U12640 ( .A(n12362), .B(n12363), .Z(n12357) );
  ANDN U12641 ( .B(n12364), .A(n12365), .Z(n12361) );
  XOR U12642 ( .A(n12033), .B(n12366), .Z(n11896) );
  XNOR U12643 ( .A(n12031), .B(n12367), .Z(n12366) );
  NANDN U12644 ( .A(n12368), .B(n11827), .Z(n12367) );
  OR U12645 ( .A(n12369), .B(n11900), .Z(n12031) );
  XOR U12646 ( .A(n11903), .B(n11827), .Z(n11900) );
  XOR U12647 ( .A(n12370), .B(n12035), .Z(n12033) );
  OR U12648 ( .A(n12362), .B(n12371), .Z(n12035) );
  XNOR U12649 ( .A(n12364), .B(n12360), .Z(n12362) );
  IV U12650 ( .A(n12037), .Z(n12360) );
  XNOR U12651 ( .A(n12346), .B(n11827), .Z(n12037) );
  XOR U12652 ( .A(n12372), .B(n12373), .Z(n11827) );
  NANDN U12653 ( .A(n12374), .B(n12375), .Z(n12373) );
  XOR U12654 ( .A(n12376), .B(n12377), .Z(n12346) );
  NANDN U12655 ( .A(n12374), .B(n12378), .Z(n12377) );
  AND U12656 ( .A(n12379), .B(n12364), .Z(n12370) );
  XNOR U12657 ( .A(n11903), .B(n11927), .Z(n12364) );
  XNOR U12658 ( .A(n12380), .B(n12376), .Z(n11927) );
  NANDN U12659 ( .A(n12381), .B(n12382), .Z(n12376) );
  XOR U12660 ( .A(n12378), .B(n12383), .Z(n12382) );
  ANDN U12661 ( .B(n12383), .A(n12384), .Z(n12380) );
  NANDN U12662 ( .A(n12381), .B(n12386), .Z(n12372) );
  XOR U12663 ( .A(n12387), .B(n12375), .Z(n12386) );
  XNOR U12664 ( .A(n12388), .B(n12389), .Z(n12374) );
  XOR U12665 ( .A(n12390), .B(n12391), .Z(n12389) );
  XNOR U12666 ( .A(n12392), .B(n12393), .Z(n12388) );
  XNOR U12667 ( .A(n12394), .B(n12395), .Z(n12393) );
  ANDN U12668 ( .B(n12387), .A(n12391), .Z(n12394) );
  ANDN U12669 ( .B(n12387), .A(n12384), .Z(n12385) );
  XNOR U12670 ( .A(n12390), .B(n12396), .Z(n12384) );
  XOR U12671 ( .A(n12397), .B(n12395), .Z(n12396) );
  NAND U12672 ( .A(n12398), .B(n12399), .Z(n12395) );
  XNOR U12673 ( .A(n12392), .B(n12375), .Z(n12399) );
  IV U12674 ( .A(n12387), .Z(n12392) );
  XNOR U12675 ( .A(n12378), .B(n12391), .Z(n12398) );
  IV U12676 ( .A(n12383), .Z(n12391) );
  XOR U12677 ( .A(n12400), .B(n12401), .Z(n12383) );
  XNOR U12678 ( .A(n12402), .B(n12403), .Z(n12401) );
  XNOR U12679 ( .A(n12404), .B(n12405), .Z(n12400) );
  ANDN U12680 ( .B(n12032), .A(n11902), .Z(n12404) );
  AND U12681 ( .A(n12375), .B(n12378), .Z(n12397) );
  XNOR U12682 ( .A(n12375), .B(n12378), .Z(n12390) );
  XNOR U12683 ( .A(n12406), .B(n12407), .Z(n12378) );
  XNOR U12684 ( .A(n12408), .B(n12403), .Z(n12407) );
  XOR U12685 ( .A(n12409), .B(n12410), .Z(n12406) );
  XNOR U12686 ( .A(n12411), .B(n12405), .Z(n12410) );
  OR U12687 ( .A(n11901), .B(n12369), .Z(n12405) );
  XNOR U12688 ( .A(n12032), .B(n12442), .Z(n12369) );
  XNOR U12689 ( .A(n11902), .B(n11828), .Z(n11901) );
  ANDN U12690 ( .B(n12412), .A(n12368), .Z(n12411) );
  XNOR U12691 ( .A(n12413), .B(n12414), .Z(n12375) );
  XNOR U12692 ( .A(n12403), .B(n12415), .Z(n12414) );
  XNOR U12693 ( .A(n12354), .B(n12409), .Z(n12415) );
  XNOR U12694 ( .A(n11902), .B(n12032), .Z(n12403) );
  XOR U12695 ( .A(n11926), .B(n12416), .Z(n12413) );
  XNOR U12696 ( .A(n12417), .B(n12418), .Z(n12416) );
  ANDN U12697 ( .B(n12419), .A(n12351), .Z(n12417) );
  XNOR U12698 ( .A(n12420), .B(n12421), .Z(n12387) );
  XNOR U12699 ( .A(n12408), .B(n12422), .Z(n12421) );
  XNOR U12700 ( .A(n12423), .B(n12402), .Z(n12422) );
  XOR U12701 ( .A(n12409), .B(n12424), .Z(n12402) );
  XNOR U12702 ( .A(n12425), .B(n12426), .Z(n12424) );
  NANDN U12703 ( .A(n12359), .B(n12038), .Z(n12426) );
  XNOR U12704 ( .A(n12427), .B(n12425), .Z(n12409) );
  OR U12705 ( .A(n12371), .B(n12363), .Z(n12425) );
  XOR U12706 ( .A(n12428), .B(n12359), .Z(n12363) );
  XNOR U12707 ( .A(n12412), .B(n12419), .Z(n12359) );
  IV U12708 ( .A(n11828), .Z(n12412) );
  XNOR U12709 ( .A(n12379), .B(n12038), .Z(n12371) );
  XNOR U12710 ( .A(n12351), .B(n12442), .Z(n12038) );
  ANDN U12711 ( .B(n12379), .A(n12365), .Z(n12427) );
  IV U12712 ( .A(n12428), .Z(n12365) );
  XOR U12713 ( .A(n12429), .B(n12354), .Z(n12428) );
  XOR U12714 ( .A(n11828), .B(n12368), .Z(n12408) );
  XOR U12715 ( .A(n12430), .B(n12431), .Z(n12368) );
  XOR U12716 ( .A(n12432), .B(n12433), .Z(n11828) );
  XOR U12717 ( .A(n12434), .B(n12431), .Z(n12433) );
  XNOR U12718 ( .A(n12345), .B(n12435), .Z(n12420) );
  XNOR U12719 ( .A(n12436), .B(n12418), .Z(n12435) );
  OR U12720 ( .A(n12355), .B(n12350), .Z(n12418) );
  XNOR U12721 ( .A(n11926), .B(n12351), .Z(n12350) );
  IV U12722 ( .A(n12423), .Z(n12351) );
  XOR U12723 ( .A(n12437), .B(n12438), .Z(n12423) );
  XNOR U12724 ( .A(n12439), .B(n12440), .Z(n12438) );
  XNOR U12725 ( .A(n11926), .B(n12441), .Z(n12437) );
  XNOR U12726 ( .A(n12354), .B(n12419), .Z(n12355) );
  IV U12727 ( .A(n12345), .Z(n12419) );
  ANDN U12728 ( .B(n12354), .A(n11926), .Z(n12436) );
  XOR U12729 ( .A(n12439), .B(n12442), .Z(n12354) );
  XOR U12730 ( .A(n12443), .B(n12444), .Z(n12439) );
  XNOR U12731 ( .A(n12445), .B(n12446), .Z(n12444) );
  XNOR U12732 ( .A(n12447), .B(n12448), .Z(n12443) );
  XNOR U12733 ( .A(key[732]), .B(n12449), .Z(n12448) );
  XNOR U12734 ( .A(n12450), .B(n12451), .Z(n12345) );
  XOR U12735 ( .A(n11902), .B(n12432), .Z(n12451) );
  IV U12736 ( .A(n12429), .Z(n11902) );
  XOR U12737 ( .A(n12441), .B(n12442), .Z(n12429) );
  XNOR U12738 ( .A(n12430), .B(n12431), .Z(n12442) );
  IV U12739 ( .A(n12434), .Z(n12430) );
  XNOR U12740 ( .A(n12452), .B(n12453), .Z(n12434) );
  XOR U12741 ( .A(n12454), .B(n12455), .Z(n12453) );
  XNOR U12742 ( .A(n12456), .B(n12457), .Z(n12452) );
  XNOR U12743 ( .A(key[733]), .B(n12458), .Z(n12457) );
  XOR U12744 ( .A(n12459), .B(n12460), .Z(n12441) );
  XOR U12745 ( .A(n12461), .B(n12462), .Z(n12460) );
  XOR U12746 ( .A(key[735]), .B(n12463), .Z(n12459) );
  XNOR U12747 ( .A(n11926), .B(n12032), .Z(n12379) );
  XNOR U12748 ( .A(n12440), .B(n12464), .Z(n12032) );
  XNOR U12749 ( .A(n12431), .B(n12450), .Z(n12464) );
  XOR U12750 ( .A(n12465), .B(n12466), .Z(n12450) );
  XOR U12751 ( .A(n12467), .B(n12468), .Z(n12466) );
  XNOR U12752 ( .A(n12469), .B(n12470), .Z(n12465) );
  XOR U12753 ( .A(key[730]), .B(n12471), .Z(n12470) );
  XOR U12754 ( .A(n12472), .B(n12473), .Z(n12431) );
  XOR U12755 ( .A(n11926), .B(n12474), .Z(n12473) );
  XNOR U12756 ( .A(n12475), .B(n12476), .Z(n12472) );
  XNOR U12757 ( .A(key[734]), .B(n12477), .Z(n12476) );
  XOR U12758 ( .A(n12478), .B(n12479), .Z(n12440) );
  XNOR U12759 ( .A(n12480), .B(n12481), .Z(n12479) );
  XOR U12760 ( .A(n12482), .B(n12432), .Z(n12481) );
  XNOR U12761 ( .A(n12483), .B(n12484), .Z(n12432) );
  XOR U12762 ( .A(n12485), .B(n12486), .Z(n12484) );
  XNOR U12763 ( .A(n12487), .B(n12488), .Z(n12483) );
  XNOR U12764 ( .A(key[729]), .B(n12489), .Z(n12488) );
  XNOR U12765 ( .A(n12490), .B(n12491), .Z(n12478) );
  XNOR U12766 ( .A(key[731]), .B(n12492), .Z(n12491) );
  XNOR U12767 ( .A(n12493), .B(n12494), .Z(n11926) );
  XOR U12768 ( .A(n12495), .B(n12496), .Z(n12494) );
  XOR U12769 ( .A(n12497), .B(n12498), .Z(n12493) );
  XNOR U12770 ( .A(key[728]), .B(n12499), .Z(n12498) );
  XNOR U12771 ( .A(n11950), .B(n11837), .Z(n10351) );
  XNOR U12772 ( .A(n11911), .B(n12500), .Z(n11837) );
  XNOR U12773 ( .A(n12501), .B(n12317), .Z(n12500) );
  XOR U12774 ( .A(n12025), .B(n11841), .Z(n12023) );
  ANDN U12775 ( .B(n12025), .A(n12503), .Z(n12501) );
  XNOR U12776 ( .A(n12315), .B(n12504), .Z(n11911) );
  XNOR U12777 ( .A(n12505), .B(n12506), .Z(n12504) );
  NAND U12778 ( .A(n12328), .B(n12507), .Z(n12506) );
  XOR U12779 ( .A(n12315), .B(n12508), .Z(n11950) );
  XOR U12780 ( .A(n12509), .B(n11913), .Z(n12508) );
  OR U12781 ( .A(n12510), .B(n12333), .Z(n11913) );
  XNOR U12782 ( .A(n11915), .B(n12331), .Z(n12333) );
  NOR U12783 ( .A(n12511), .B(n12331), .Z(n12509) );
  XOR U12784 ( .A(n12512), .B(n12505), .Z(n12315) );
  OR U12785 ( .A(n12336), .B(n12513), .Z(n12505) );
  XNOR U12786 ( .A(n12514), .B(n12328), .Z(n12336) );
  XNOR U12787 ( .A(n12331), .B(n11841), .Z(n12328) );
  XOR U12788 ( .A(n12515), .B(n12516), .Z(n11841) );
  NANDN U12789 ( .A(n12517), .B(n12518), .Z(n12516) );
  XNOR U12790 ( .A(n12519), .B(n12520), .Z(n12331) );
  OR U12791 ( .A(n12517), .B(n12521), .Z(n12520) );
  ANDN U12792 ( .B(n12514), .A(n12522), .Z(n12512) );
  IV U12793 ( .A(n12339), .Z(n12514) );
  XOR U12794 ( .A(n11915), .B(n12025), .Z(n12339) );
  XNOR U12795 ( .A(n12523), .B(n12515), .Z(n12025) );
  NANDN U12796 ( .A(n12524), .B(n12525), .Z(n12515) );
  ANDN U12797 ( .B(n12526), .A(n12527), .Z(n12523) );
  NANDN U12798 ( .A(n12524), .B(n12529), .Z(n12519) );
  XOR U12799 ( .A(n12530), .B(n12517), .Z(n12524) );
  XNOR U12800 ( .A(n12531), .B(n12532), .Z(n12517) );
  XOR U12801 ( .A(n12533), .B(n12526), .Z(n12532) );
  XNOR U12802 ( .A(n12534), .B(n12535), .Z(n12531) );
  XNOR U12803 ( .A(n12536), .B(n12537), .Z(n12535) );
  ANDN U12804 ( .B(n12526), .A(n12538), .Z(n12536) );
  IV U12805 ( .A(n12539), .Z(n12526) );
  ANDN U12806 ( .B(n12530), .A(n12538), .Z(n12528) );
  IV U12807 ( .A(n12534), .Z(n12538) );
  IV U12808 ( .A(n12527), .Z(n12530) );
  XNOR U12809 ( .A(n12533), .B(n12540), .Z(n12527) );
  XOR U12810 ( .A(n12541), .B(n12537), .Z(n12540) );
  NAND U12811 ( .A(n12529), .B(n12525), .Z(n12537) );
  XNOR U12812 ( .A(n12518), .B(n12539), .Z(n12525) );
  XOR U12813 ( .A(n12542), .B(n12543), .Z(n12539) );
  XOR U12814 ( .A(n12544), .B(n12545), .Z(n12543) );
  XNOR U12815 ( .A(n12332), .B(n12546), .Z(n12545) );
  XNOR U12816 ( .A(n12547), .B(n12548), .Z(n12542) );
  XNOR U12817 ( .A(n12549), .B(n12550), .Z(n12548) );
  ANDN U12818 ( .B(n12551), .A(n11916), .Z(n12549) );
  XNOR U12819 ( .A(n12534), .B(n12521), .Z(n12529) );
  XOR U12820 ( .A(n12552), .B(n12553), .Z(n12534) );
  XNOR U12821 ( .A(n12554), .B(n12546), .Z(n12553) );
  XOR U12822 ( .A(n12555), .B(n12556), .Z(n12546) );
  XNOR U12823 ( .A(n12557), .B(n12558), .Z(n12556) );
  NAND U12824 ( .A(n12507), .B(n12327), .Z(n12558) );
  XNOR U12825 ( .A(n12559), .B(n12560), .Z(n12552) );
  ANDN U12826 ( .B(n12561), .A(n12503), .Z(n12559) );
  ANDN U12827 ( .B(n12518), .A(n12521), .Z(n12541) );
  XOR U12828 ( .A(n12521), .B(n12518), .Z(n12533) );
  XNOR U12829 ( .A(n12562), .B(n12563), .Z(n12518) );
  XNOR U12830 ( .A(n12555), .B(n12564), .Z(n12563) );
  XOR U12831 ( .A(n12554), .B(n12323), .Z(n12564) );
  XOR U12832 ( .A(n11916), .B(n12565), .Z(n12562) );
  XNOR U12833 ( .A(n12566), .B(n12550), .Z(n12565) );
  OR U12834 ( .A(n12334), .B(n12510), .Z(n12550) );
  XNOR U12835 ( .A(n11916), .B(n12511), .Z(n12510) );
  XOR U12836 ( .A(n12323), .B(n12332), .Z(n12334) );
  ANDN U12837 ( .B(n12332), .A(n12511), .Z(n12566) );
  XOR U12838 ( .A(n12567), .B(n12568), .Z(n12521) );
  XOR U12839 ( .A(n12555), .B(n12544), .Z(n12568) );
  XOR U12840 ( .A(n12319), .B(n11842), .Z(n12544) );
  XOR U12841 ( .A(n12569), .B(n12557), .Z(n12555) );
  NANDN U12842 ( .A(n12513), .B(n12337), .Z(n12557) );
  XOR U12843 ( .A(n12338), .B(n12327), .Z(n12337) );
  XNOR U12844 ( .A(n12561), .B(n12570), .Z(n12332) );
  XNOR U12845 ( .A(n12571), .B(n12572), .Z(n12570) );
  XOR U12846 ( .A(n12522), .B(n12507), .Z(n12513) );
  XNOR U12847 ( .A(n12511), .B(n12319), .Z(n12507) );
  IV U12848 ( .A(n12547), .Z(n12511) );
  XOR U12849 ( .A(n12573), .B(n12574), .Z(n12547) );
  XOR U12850 ( .A(n12575), .B(n12576), .Z(n12574) );
  XNOR U12851 ( .A(n11916), .B(n12577), .Z(n12573) );
  ANDN U12852 ( .B(n12338), .A(n12522), .Z(n12569) );
  XNOR U12853 ( .A(n11916), .B(n12503), .Z(n12522) );
  XOR U12854 ( .A(n12561), .B(n12551), .Z(n12338) );
  IV U12855 ( .A(n12323), .Z(n12551) );
  XOR U12856 ( .A(n12578), .B(n12579), .Z(n12323) );
  XOR U12857 ( .A(n12580), .B(n12576), .Z(n12579) );
  XNOR U12858 ( .A(n12581), .B(n12582), .Z(n12576) );
  XNOR U12859 ( .A(n12583), .B(n12584), .Z(n12582) );
  XOR U12860 ( .A(n12585), .B(n12586), .Z(n12581) );
  XNOR U12861 ( .A(key[692]), .B(n12587), .Z(n12586) );
  IV U12862 ( .A(n12026), .Z(n12561) );
  XOR U12863 ( .A(n12554), .B(n12588), .Z(n12567) );
  XNOR U12864 ( .A(n12589), .B(n12560), .Z(n12588) );
  OR U12865 ( .A(n12024), .B(n12502), .Z(n12560) );
  XNOR U12866 ( .A(n12590), .B(n12319), .Z(n12502) );
  XNOR U12867 ( .A(n12026), .B(n11842), .Z(n12024) );
  ANDN U12868 ( .B(n12319), .A(n11842), .Z(n12589) );
  XOR U12869 ( .A(n12578), .B(n12591), .Z(n11842) );
  XOR U12870 ( .A(n12571), .B(n12592), .Z(n12591) );
  XOR U12871 ( .A(n12580), .B(n12578), .Z(n12319) );
  XNOR U12872 ( .A(n12503), .B(n12026), .Z(n12554) );
  XOR U12873 ( .A(n12578), .B(n12593), .Z(n12026) );
  XNOR U12874 ( .A(n12580), .B(n12575), .Z(n12593) );
  XOR U12875 ( .A(n12594), .B(n12595), .Z(n12575) );
  XNOR U12876 ( .A(n12596), .B(n12597), .Z(n12595) );
  XNOR U12877 ( .A(key[695]), .B(n12598), .Z(n12594) );
  XNOR U12878 ( .A(n12599), .B(n12600), .Z(n12578) );
  XOR U12879 ( .A(n12601), .B(n12602), .Z(n12600) );
  XNOR U12880 ( .A(key[693]), .B(n12603), .Z(n12599) );
  IV U12881 ( .A(n12590), .Z(n12503) );
  XNOR U12882 ( .A(n12572), .B(n12604), .Z(n12590) );
  XOR U12883 ( .A(n12577), .B(n12592), .Z(n12604) );
  IV U12884 ( .A(n12580), .Z(n12592) );
  XOR U12885 ( .A(n12605), .B(n12606), .Z(n12580) );
  XNOR U12886 ( .A(n11916), .B(n12607), .Z(n12606) );
  XNOR U12887 ( .A(n12608), .B(n12609), .Z(n11916) );
  XOR U12888 ( .A(n12610), .B(n12611), .Z(n12609) );
  XOR U12889 ( .A(key[688]), .B(n12612), .Z(n12608) );
  XNOR U12890 ( .A(n12613), .B(n12614), .Z(n12605) );
  XNOR U12891 ( .A(key[694]), .B(n12615), .Z(n12614) );
  XOR U12892 ( .A(n12616), .B(n12617), .Z(n12577) );
  XNOR U12893 ( .A(n12618), .B(n12619), .Z(n12617) );
  XNOR U12894 ( .A(n12571), .B(n12620), .Z(n12619) );
  XOR U12895 ( .A(n12621), .B(n12622), .Z(n12571) );
  XNOR U12896 ( .A(n12623), .B(n12624), .Z(n12622) );
  XNOR U12897 ( .A(key[689]), .B(n12625), .Z(n12621) );
  XOR U12898 ( .A(n12626), .B(n12627), .Z(n12616) );
  XNOR U12899 ( .A(key[691]), .B(n12628), .Z(n12627) );
  XOR U12900 ( .A(n12629), .B(n12630), .Z(n12572) );
  XNOR U12901 ( .A(n12631), .B(n12632), .Z(n12630) );
  XOR U12902 ( .A(key[690]), .B(n12633), .Z(n12629) );
  XNOR U12903 ( .A(n7233), .B(n6317), .Z(n7218) );
  XOR U12904 ( .A(n11585), .B(n12634), .Z(n6317) );
  XOR U12905 ( .A(n11587), .B(n11588), .Z(n12634) );
  XOR U12906 ( .A(n12635), .B(n12636), .Z(n11588) );
  XNOR U12907 ( .A(n12637), .B(n12638), .Z(n12636) );
  NANDN U12908 ( .A(n11607), .B(n12639), .Z(n12638) );
  XNOR U12909 ( .A(n11706), .B(n12640), .Z(n11587) );
  XOR U12910 ( .A(n12641), .B(n12642), .Z(n12640) );
  ANDN U12911 ( .B(n12643), .A(n11600), .Z(n12641) );
  XNOR U12912 ( .A(n11595), .B(n12644), .Z(n11706) );
  XNOR U12913 ( .A(n12645), .B(n12646), .Z(n12644) );
  NAND U12914 ( .A(n12647), .B(n12648), .Z(n12646) );
  XOR U12915 ( .A(n11702), .B(n11557), .Z(n11585) );
  XOR U12916 ( .A(n11595), .B(n12649), .Z(n11557) );
  XNOR U12917 ( .A(n12642), .B(n12650), .Z(n12649) );
  NANDN U12918 ( .A(n12651), .B(n12652), .Z(n12650) );
  OR U12919 ( .A(n12653), .B(n12654), .Z(n12642) );
  XOR U12920 ( .A(n12655), .B(n12645), .Z(n11595) );
  NANDN U12921 ( .A(n12656), .B(n12657), .Z(n12645) );
  AND U12922 ( .A(n12658), .B(n12659), .Z(n12655) );
  IV U12923 ( .A(n6309), .Z(n7233) );
  XOR U12924 ( .A(n11523), .B(n12660), .Z(n6309) );
  XOR U12925 ( .A(n11505), .B(n11506), .Z(n12660) );
  XNOR U12926 ( .A(n12662), .B(n12663), .Z(n12661) );
  NANDN U12927 ( .A(n11616), .B(n12664), .Z(n12663) );
  XOR U12928 ( .A(n11618), .B(n12665), .Z(n11548) );
  XNOR U12929 ( .A(n12666), .B(n12667), .Z(n12665) );
  NAND U12930 ( .A(n12668), .B(n11722), .Z(n12667) );
  IV U12931 ( .A(n11525), .Z(n11505) );
  XOR U12932 ( .A(n11718), .B(n12669), .Z(n11525) );
  XOR U12933 ( .A(n11716), .B(n12670), .Z(n12669) );
  NAND U12934 ( .A(n12671), .B(n11621), .Z(n12670) );
  XOR U12935 ( .A(n11552), .B(n11621), .Z(n11623) );
  XOR U12936 ( .A(n11713), .B(n11503), .Z(n11523) );
  XNOR U12937 ( .A(n11618), .B(n12673), .Z(n11503) );
  XNOR U12938 ( .A(n12662), .B(n12674), .Z(n12673) );
  NANDN U12939 ( .A(n12675), .B(n12676), .Z(n12674) );
  OR U12940 ( .A(n12677), .B(n12678), .Z(n12662) );
  XNOR U12941 ( .A(n12679), .B(n12666), .Z(n11618) );
  NANDN U12942 ( .A(n12680), .B(n12681), .Z(n12666) );
  ANDN U12943 ( .B(n12682), .A(n12683), .Z(n12679) );
  XOR U12944 ( .A(n11718), .B(n12684), .Z(n11713) );
  XOR U12945 ( .A(n12685), .B(n11614), .Z(n12684) );
  OR U12946 ( .A(n12686), .B(n12677), .Z(n11614) );
  XNOR U12947 ( .A(n11616), .B(n12675), .Z(n12677) );
  NOR U12948 ( .A(n12687), .B(n12675), .Z(n12685) );
  XOR U12949 ( .A(n12688), .B(n11720), .Z(n11718) );
  OR U12950 ( .A(n12680), .B(n12689), .Z(n11720) );
  XNOR U12951 ( .A(n12690), .B(n11722), .Z(n12680) );
  XNOR U12952 ( .A(n12675), .B(n11621), .Z(n11722) );
  XOR U12953 ( .A(n12691), .B(n12692), .Z(n11621) );
  NANDN U12954 ( .A(n12693), .B(n12694), .Z(n12692) );
  XNOR U12955 ( .A(n12695), .B(n12696), .Z(n12675) );
  OR U12956 ( .A(n12693), .B(n12697), .Z(n12696) );
  ANDN U12957 ( .B(n12690), .A(n12698), .Z(n12688) );
  IV U12958 ( .A(n12683), .Z(n12690) );
  XOR U12959 ( .A(n11616), .B(n11552), .Z(n12683) );
  XNOR U12960 ( .A(n12699), .B(n12691), .Z(n11552) );
  NANDN U12961 ( .A(n12700), .B(n12701), .Z(n12691) );
  ANDN U12962 ( .B(n12702), .A(n12703), .Z(n12699) );
  NANDN U12963 ( .A(n12700), .B(n12705), .Z(n12695) );
  XOR U12964 ( .A(n12706), .B(n12693), .Z(n12700) );
  XNOR U12965 ( .A(n12707), .B(n12708), .Z(n12693) );
  XOR U12966 ( .A(n12709), .B(n12702), .Z(n12708) );
  XNOR U12967 ( .A(n12710), .B(n12711), .Z(n12707) );
  XNOR U12968 ( .A(n12712), .B(n12713), .Z(n12711) );
  ANDN U12969 ( .B(n12702), .A(n12714), .Z(n12712) );
  IV U12970 ( .A(n12715), .Z(n12702) );
  ANDN U12971 ( .B(n12706), .A(n12714), .Z(n12704) );
  IV U12972 ( .A(n12710), .Z(n12714) );
  IV U12973 ( .A(n12703), .Z(n12706) );
  XNOR U12974 ( .A(n12709), .B(n12716), .Z(n12703) );
  XOR U12975 ( .A(n12717), .B(n12713), .Z(n12716) );
  NAND U12976 ( .A(n12705), .B(n12701), .Z(n12713) );
  XNOR U12977 ( .A(n12694), .B(n12715), .Z(n12701) );
  XOR U12978 ( .A(n12718), .B(n12719), .Z(n12715) );
  XOR U12979 ( .A(n12720), .B(n12721), .Z(n12719) );
  XNOR U12980 ( .A(n12676), .B(n12722), .Z(n12721) );
  XNOR U12981 ( .A(n12723), .B(n12724), .Z(n12718) );
  XNOR U12982 ( .A(n12725), .B(n12726), .Z(n12724) );
  ANDN U12983 ( .B(n12664), .A(n11617), .Z(n12725) );
  XNOR U12984 ( .A(n12710), .B(n12697), .Z(n12705) );
  XOR U12985 ( .A(n12727), .B(n12728), .Z(n12710) );
  XNOR U12986 ( .A(n12729), .B(n12722), .Z(n12728) );
  XOR U12987 ( .A(n12730), .B(n12731), .Z(n12722) );
  XNOR U12988 ( .A(n12732), .B(n12733), .Z(n12731) );
  NAND U12989 ( .A(n11723), .B(n12668), .Z(n12733) );
  XNOR U12990 ( .A(n12734), .B(n12735), .Z(n12727) );
  ANDN U12991 ( .B(n12736), .A(n11717), .Z(n12734) );
  ANDN U12992 ( .B(n12694), .A(n12697), .Z(n12717) );
  XOR U12993 ( .A(n12697), .B(n12694), .Z(n12709) );
  XNOR U12994 ( .A(n12737), .B(n12738), .Z(n12694) );
  XNOR U12995 ( .A(n12730), .B(n12739), .Z(n12738) );
  XNOR U12996 ( .A(n12729), .B(n12664), .Z(n12739) );
  XNOR U12997 ( .A(n12740), .B(n12741), .Z(n12737) );
  XNOR U12998 ( .A(n12742), .B(n12726), .Z(n12741) );
  OR U12999 ( .A(n12678), .B(n12686), .Z(n12726) );
  XNOR U13000 ( .A(n12740), .B(n12723), .Z(n12686) );
  XNOR U13001 ( .A(n12664), .B(n12676), .Z(n12678) );
  ANDN U13002 ( .B(n12676), .A(n12687), .Z(n12742) );
  XOR U13003 ( .A(n12743), .B(n12744), .Z(n12697) );
  XOR U13004 ( .A(n12730), .B(n12720), .Z(n12744) );
  XOR U13005 ( .A(n12671), .B(n11622), .Z(n12720) );
  XOR U13006 ( .A(n12745), .B(n12732), .Z(n12730) );
  NANDN U13007 ( .A(n12689), .B(n12681), .Z(n12732) );
  XOR U13008 ( .A(n12682), .B(n12668), .Z(n12681) );
  XNOR U13009 ( .A(n12736), .B(n12746), .Z(n12676) );
  XNOR U13010 ( .A(n12747), .B(n12748), .Z(n12746) );
  XOR U13011 ( .A(n12698), .B(n11723), .Z(n12689) );
  XNOR U13012 ( .A(n12687), .B(n12671), .Z(n11723) );
  IV U13013 ( .A(n12723), .Z(n12687) );
  XOR U13014 ( .A(n12749), .B(n12750), .Z(n12723) );
  XOR U13015 ( .A(n12751), .B(n12752), .Z(n12750) );
  XOR U13016 ( .A(n12740), .B(n12753), .Z(n12749) );
  ANDN U13017 ( .B(n12682), .A(n12698), .Z(n12745) );
  XNOR U13018 ( .A(n12740), .B(n12754), .Z(n12698) );
  XOR U13019 ( .A(n12736), .B(n12664), .Z(n12682) );
  XNOR U13020 ( .A(n12755), .B(n12756), .Z(n12664) );
  XOR U13021 ( .A(n12757), .B(n12752), .Z(n12756) );
  XNOR U13022 ( .A(n12758), .B(n12759), .Z(n12752) );
  XNOR U13023 ( .A(n10196), .B(n10195), .Z(n12759) );
  XNOR U13024 ( .A(n11122), .B(n9292), .Z(n10195) );
  XNOR U13025 ( .A(n12760), .B(n9259), .Z(n9292) );
  XOR U13026 ( .A(n12761), .B(n12762), .Z(n11122) );
  XNOR U13027 ( .A(n11144), .B(n11138), .Z(n10196) );
  XNOR U13028 ( .A(n9291), .B(n12763), .Z(n12758) );
  XNOR U13029 ( .A(key[820]), .B(n11120), .Z(n12763) );
  XNOR U13030 ( .A(n9314), .B(n10180), .Z(n9291) );
  XOR U13031 ( .A(n12764), .B(n12765), .Z(n10180) );
  XNOR U13032 ( .A(n12766), .B(n12767), .Z(n12765) );
  XNOR U13033 ( .A(n12768), .B(n12769), .Z(n12764) );
  XOR U13034 ( .A(n12770), .B(n12771), .Z(n12769) );
  ANDN U13035 ( .B(n12772), .A(n12773), .Z(n12771) );
  IV U13036 ( .A(n11553), .Z(n12736) );
  XOR U13037 ( .A(n12729), .B(n12774), .Z(n12743) );
  XNOR U13038 ( .A(n12775), .B(n12735), .Z(n12774) );
  OR U13039 ( .A(n11624), .B(n12672), .Z(n12735) );
  XNOR U13040 ( .A(n12754), .B(n12671), .Z(n12672) );
  XNOR U13041 ( .A(n11553), .B(n11622), .Z(n11624) );
  ANDN U13042 ( .B(n12671), .A(n11622), .Z(n12775) );
  XOR U13043 ( .A(n12755), .B(n12776), .Z(n11622) );
  XOR U13044 ( .A(n12747), .B(n12777), .Z(n12776) );
  XOR U13045 ( .A(n12757), .B(n12755), .Z(n12671) );
  XNOR U13046 ( .A(n11717), .B(n11553), .Z(n12729) );
  XOR U13047 ( .A(n12755), .B(n12778), .Z(n11553) );
  XNOR U13048 ( .A(n12757), .B(n12751), .Z(n12778) );
  XOR U13049 ( .A(n12779), .B(n12780), .Z(n12751) );
  XNOR U13050 ( .A(n12781), .B(n10190), .Z(n12780) );
  XNOR U13051 ( .A(n11148), .B(n9285), .Z(n10190) );
  XOR U13052 ( .A(n12782), .B(n12783), .Z(n9285) );
  XOR U13053 ( .A(n12784), .B(n12785), .Z(n12783) );
  XNOR U13054 ( .A(n12786), .B(n12787), .Z(n12782) );
  XOR U13055 ( .A(n12788), .B(n12789), .Z(n11148) );
  XOR U13056 ( .A(n12790), .B(n12791), .Z(n12789) );
  XNOR U13057 ( .A(n12792), .B(n12793), .Z(n12788) );
  XNOR U13058 ( .A(key[823]), .B(n9314), .Z(n12779) );
  XNOR U13059 ( .A(n12794), .B(n12795), .Z(n12755) );
  XOR U13060 ( .A(n11138), .B(n10181), .Z(n12795) );
  XOR U13061 ( .A(n11124), .B(n9276), .Z(n10181) );
  XNOR U13062 ( .A(n12796), .B(n12797), .Z(n9276) );
  XNOR U13063 ( .A(n12798), .B(n12785), .Z(n12797) );
  XNOR U13064 ( .A(n12799), .B(n12800), .Z(n12785) );
  XNOR U13065 ( .A(n12801), .B(n12802), .Z(n12800) );
  NANDN U13066 ( .A(n12803), .B(n12804), .Z(n12802) );
  XOR U13067 ( .A(n12805), .B(n12806), .Z(n12796) );
  XOR U13068 ( .A(n12807), .B(n12808), .Z(n12806) );
  ANDN U13069 ( .B(n12809), .A(n12810), .Z(n12808) );
  XOR U13070 ( .A(n12811), .B(n12812), .Z(n11124) );
  XNOR U13071 ( .A(n12761), .B(n12791), .Z(n12812) );
  XNOR U13072 ( .A(n12813), .B(n12814), .Z(n12791) );
  XNOR U13073 ( .A(n12815), .B(n12816), .Z(n12814) );
  NANDN U13074 ( .A(n12817), .B(n12818), .Z(n12816) );
  XNOR U13075 ( .A(n12819), .B(n12820), .Z(n12811) );
  XNOR U13076 ( .A(n12821), .B(n12822), .Z(n12820) );
  ANDN U13077 ( .B(n12823), .A(n12824), .Z(n12822) );
  XNOR U13078 ( .A(n12825), .B(n12826), .Z(n11138) );
  XNOR U13079 ( .A(n12827), .B(n12828), .Z(n12826) );
  XNOR U13080 ( .A(n12829), .B(n12830), .Z(n12825) );
  XOR U13081 ( .A(n12831), .B(n12832), .Z(n12830) );
  ANDN U13082 ( .B(n12833), .A(n12834), .Z(n12832) );
  XNOR U13083 ( .A(key[821]), .B(n11147), .Z(n12794) );
  XOR U13084 ( .A(n10177), .B(n10184), .Z(n11147) );
  IV U13085 ( .A(n9280), .Z(n10177) );
  XOR U13086 ( .A(n12835), .B(n12836), .Z(n9280) );
  IV U13087 ( .A(n12754), .Z(n11717) );
  XNOR U13088 ( .A(n12748), .B(n12837), .Z(n12754) );
  XOR U13089 ( .A(n12753), .B(n12777), .Z(n12837) );
  IV U13090 ( .A(n12757), .Z(n12777) );
  XOR U13091 ( .A(n12838), .B(n12839), .Z(n12757) );
  XNOR U13092 ( .A(n10175), .B(n11617), .Z(n12839) );
  IV U13093 ( .A(n12740), .Z(n11617) );
  XOR U13094 ( .A(n12840), .B(n12841), .Z(n12740) );
  XNOR U13095 ( .A(n11123), .B(n9303), .Z(n12841) );
  XOR U13096 ( .A(n10209), .B(n10214), .Z(n9303) );
  IV U13097 ( .A(n9312), .Z(n10209) );
  XOR U13098 ( .A(n12842), .B(n12843), .Z(n9312) );
  XNOR U13099 ( .A(n12844), .B(n12835), .Z(n12843) );
  XNOR U13100 ( .A(n12845), .B(n12761), .Z(n11123) );
  XNOR U13101 ( .A(n12813), .B(n12846), .Z(n12761) );
  XOR U13102 ( .A(n12847), .B(n12848), .Z(n12846) );
  ANDN U13103 ( .B(n12849), .A(n12850), .Z(n12847) );
  XOR U13104 ( .A(n12851), .B(n12852), .Z(n12813) );
  XNOR U13105 ( .A(n12853), .B(n12854), .Z(n12852) );
  NANDN U13106 ( .A(n12855), .B(n12856), .Z(n12854) );
  XNOR U13107 ( .A(key[816]), .B(n10191), .Z(n12840) );
  XNOR U13108 ( .A(n10216), .B(n11144), .Z(n10191) );
  IV U13109 ( .A(n11134), .Z(n10216) );
  XNOR U13110 ( .A(n12805), .B(n12857), .Z(n11134) );
  IV U13111 ( .A(n12760), .Z(n12805) );
  XNOR U13112 ( .A(n12859), .B(n12860), .Z(n12858) );
  ANDN U13113 ( .B(n12861), .A(n12862), .Z(n12859) );
  XOR U13114 ( .A(n12863), .B(n12864), .Z(n12799) );
  XNOR U13115 ( .A(n12865), .B(n12866), .Z(n12864) );
  NAND U13116 ( .A(n12867), .B(n12868), .Z(n12866) );
  XOR U13117 ( .A(n11137), .B(n12781), .Z(n10175) );
  XNOR U13118 ( .A(n11144), .B(n11133), .Z(n12781) );
  XNOR U13119 ( .A(n12869), .B(n12870), .Z(n11133) );
  XNOR U13120 ( .A(n12871), .B(n12828), .Z(n12870) );
  XNOR U13121 ( .A(n12872), .B(n12873), .Z(n12828) );
  XNOR U13122 ( .A(n12874), .B(n12875), .Z(n12873) );
  OR U13123 ( .A(n12876), .B(n12877), .Z(n12875) );
  XOR U13124 ( .A(n12878), .B(n12879), .Z(n12869) );
  XOR U13125 ( .A(n9270), .B(n11145), .Z(n11137) );
  IV U13126 ( .A(n9278), .Z(n11145) );
  XNOR U13127 ( .A(n12793), .B(n12880), .Z(n9278) );
  IV U13128 ( .A(n10182), .Z(n9270) );
  XNOR U13129 ( .A(n12881), .B(n12784), .Z(n10182) );
  XOR U13130 ( .A(n9271), .B(n12882), .Z(n12838) );
  XNOR U13131 ( .A(key[822]), .B(n10184), .Z(n12882) );
  XNOR U13132 ( .A(n12871), .B(n12883), .Z(n10184) );
  XOR U13133 ( .A(n9314), .B(n10189), .Z(n9271) );
  XOR U13134 ( .A(n12884), .B(n12885), .Z(n10189) );
  XNOR U13135 ( .A(n12886), .B(n12767), .Z(n12885) );
  XNOR U13136 ( .A(n12887), .B(n12888), .Z(n12767) );
  XNOR U13137 ( .A(n12889), .B(n12890), .Z(n12888) );
  NANDN U13138 ( .A(n12891), .B(n12892), .Z(n12890) );
  XOR U13139 ( .A(n12844), .B(n12835), .Z(n12884) );
  XOR U13140 ( .A(n12893), .B(n12894), .Z(n12835) );
  XOR U13141 ( .A(n12895), .B(n12896), .Z(n12753) );
  XNOR U13142 ( .A(n12747), .B(n12897), .Z(n12896) );
  XNOR U13143 ( .A(n10210), .B(n10201), .Z(n12897) );
  XOR U13144 ( .A(n9307), .B(n9261), .Z(n10201) );
  XNOR U13145 ( .A(n12898), .B(n12899), .Z(n9261) );
  XOR U13146 ( .A(n12790), .B(n12880), .Z(n12899) );
  XNOR U13147 ( .A(n12900), .B(n12901), .Z(n12880) );
  XOR U13148 ( .A(n12902), .B(n12821), .Z(n12901) );
  NANDN U13149 ( .A(n12903), .B(n12904), .Z(n12821) );
  NOR U13150 ( .A(n12905), .B(n12850), .Z(n12902) );
  XNOR U13151 ( .A(n12792), .B(n12906), .Z(n12898) );
  IV U13152 ( .A(n10167), .Z(n9307) );
  XNOR U13153 ( .A(n12907), .B(n12908), .Z(n10167) );
  XNOR U13154 ( .A(n12787), .B(n12881), .Z(n12908) );
  XNOR U13155 ( .A(n12909), .B(n12910), .Z(n12881) );
  XNOR U13156 ( .A(n12911), .B(n12807), .Z(n12910) );
  ANDN U13157 ( .B(n12912), .A(n12913), .Z(n12807) );
  NOR U13158 ( .A(n12914), .B(n12862), .Z(n12911) );
  IV U13159 ( .A(n12915), .Z(n12787) );
  XOR U13160 ( .A(n12786), .B(n12916), .Z(n12907) );
  XOR U13161 ( .A(n11144), .B(n11120), .Z(n10210) );
  XOR U13162 ( .A(n12829), .B(n10206), .Z(n11120) );
  XNOR U13163 ( .A(n12917), .B(n12829), .Z(n11144) );
  XNOR U13164 ( .A(n12872), .B(n12918), .Z(n12829) );
  XNOR U13165 ( .A(n12919), .B(n12920), .Z(n12918) );
  NOR U13166 ( .A(n12921), .B(n12922), .Z(n12919) );
  XNOR U13167 ( .A(n12923), .B(n12924), .Z(n12872) );
  XNOR U13168 ( .A(n12925), .B(n12926), .Z(n12924) );
  NAND U13169 ( .A(n12927), .B(n12928), .Z(n12926) );
  XOR U13170 ( .A(n12929), .B(n12930), .Z(n12747) );
  XNOR U13171 ( .A(n9260), .B(n10207), .Z(n12930) );
  XOR U13172 ( .A(n9316), .B(n9304), .Z(n10207) );
  XNOR U13173 ( .A(n12784), .B(n12931), .Z(n9304) );
  XNOR U13174 ( .A(n12786), .B(n12915), .Z(n12931) );
  XNOR U13175 ( .A(n12933), .B(n12934), .Z(n12932) );
  NANDN U13176 ( .A(n12935), .B(n12804), .Z(n12934) );
  XNOR U13177 ( .A(n12798), .B(n12936), .Z(n12909) );
  XNOR U13178 ( .A(n12937), .B(n12938), .Z(n12936) );
  NAND U13179 ( .A(n12939), .B(n12867), .Z(n12938) );
  XOR U13180 ( .A(n12857), .B(n12916), .Z(n12784) );
  XOR U13181 ( .A(n12798), .B(n12940), .Z(n12916) );
  XNOR U13182 ( .A(n12933), .B(n12941), .Z(n12940) );
  NANDN U13183 ( .A(n12942), .B(n12943), .Z(n12941) );
  OR U13184 ( .A(n12944), .B(n12945), .Z(n12933) );
  XOR U13185 ( .A(n12946), .B(n12937), .Z(n12798) );
  NANDN U13186 ( .A(n12947), .B(n12948), .Z(n12937) );
  ANDN U13187 ( .B(n12949), .A(n12950), .Z(n12946) );
  XNOR U13188 ( .A(n12790), .B(n12951), .Z(n9316) );
  XOR U13189 ( .A(n12792), .B(n12793), .Z(n12951) );
  XOR U13190 ( .A(n12952), .B(n12906), .Z(n12793) );
  XNOR U13191 ( .A(n12819), .B(n12953), .Z(n12906) );
  XNOR U13192 ( .A(n12954), .B(n12955), .Z(n12953) );
  NANDN U13193 ( .A(n12956), .B(n12957), .Z(n12955) );
  XNOR U13194 ( .A(n12954), .B(n12959), .Z(n12958) );
  NAND U13195 ( .A(n12960), .B(n12818), .Z(n12959) );
  OR U13196 ( .A(n12961), .B(n12962), .Z(n12954) );
  XNOR U13197 ( .A(n12819), .B(n12963), .Z(n12900) );
  XNOR U13198 ( .A(n12964), .B(n12965), .Z(n12963) );
  NANDN U13199 ( .A(n12966), .B(n12967), .Z(n12965) );
  XOR U13200 ( .A(n12968), .B(n12964), .Z(n12819) );
  OR U13201 ( .A(n12969), .B(n12970), .Z(n12964) );
  ANDN U13202 ( .B(n12971), .A(n12972), .Z(n12968) );
  XNOR U13203 ( .A(n9302), .B(n10206), .Z(n9260) );
  XNOR U13204 ( .A(key[817]), .B(n10214), .Z(n12929) );
  XOR U13205 ( .A(n12878), .B(n12974), .Z(n12973) );
  XNOR U13206 ( .A(n12917), .B(n12975), .Z(n12871) );
  XNOR U13207 ( .A(n9297), .B(n12976), .Z(n12895) );
  XNOR U13208 ( .A(key[819]), .B(n10164), .Z(n12976) );
  XOR U13209 ( .A(n9314), .B(n10198), .Z(n9297) );
  XOR U13210 ( .A(n12768), .B(n9302), .Z(n10198) );
  XOR U13211 ( .A(n12893), .B(n12842), .Z(n9302) );
  IV U13212 ( .A(n12977), .Z(n12893) );
  XOR U13213 ( .A(n12768), .B(n12977), .Z(n9314) );
  XOR U13214 ( .A(n12978), .B(n12979), .Z(n12977) );
  XOR U13215 ( .A(n12980), .B(n12889), .Z(n12979) );
  OR U13216 ( .A(n12981), .B(n12982), .Z(n12889) );
  ANDN U13217 ( .B(n12983), .A(n12984), .Z(n12980) );
  XNOR U13218 ( .A(n12887), .B(n12985), .Z(n12768) );
  XNOR U13219 ( .A(n12986), .B(n12987), .Z(n12985) );
  ANDN U13220 ( .B(n12988), .A(n12989), .Z(n12986) );
  XOR U13221 ( .A(n12990), .B(n12991), .Z(n12887) );
  XNOR U13222 ( .A(n12992), .B(n12993), .Z(n12991) );
  NAND U13223 ( .A(n12994), .B(n12995), .Z(n12993) );
  XOR U13224 ( .A(n12996), .B(n12997), .Z(n12748) );
  XOR U13225 ( .A(n10206), .B(n10165), .Z(n12997) );
  XOR U13226 ( .A(n12762), .B(n9259), .Z(n10165) );
  XOR U13227 ( .A(n12998), .B(n12999), .Z(n12915) );
  XOR U13228 ( .A(n12860), .B(n13000), .Z(n12999) );
  NANDN U13229 ( .A(n13001), .B(n12809), .Z(n13000) );
  XNOR U13230 ( .A(n12862), .B(n12809), .Z(n12912) );
  XOR U13231 ( .A(n12998), .B(n13003), .Z(n12857) );
  XOR U13232 ( .A(n13004), .B(n12801), .Z(n13003) );
  OR U13233 ( .A(n13005), .B(n12944), .Z(n12801) );
  XNOR U13234 ( .A(n12804), .B(n12943), .Z(n12944) );
  ANDN U13235 ( .B(n12943), .A(n13006), .Z(n13004) );
  IV U13236 ( .A(n12863), .Z(n12998) );
  XNOR U13237 ( .A(n13007), .B(n12865), .Z(n12863) );
  OR U13238 ( .A(n13008), .B(n12947), .Z(n12865) );
  XOR U13239 ( .A(n12950), .B(n12867), .Z(n12947) );
  XOR U13240 ( .A(n12943), .B(n12809), .Z(n12867) );
  XOR U13241 ( .A(n13009), .B(n13010), .Z(n12809) );
  NANDN U13242 ( .A(n13011), .B(n13012), .Z(n13010) );
  XOR U13243 ( .A(n13013), .B(n13014), .Z(n12943) );
  NANDN U13244 ( .A(n13011), .B(n13015), .Z(n13014) );
  NOR U13245 ( .A(n12950), .B(n13016), .Z(n13007) );
  XOR U13246 ( .A(n12862), .B(n12804), .Z(n12950) );
  XNOR U13247 ( .A(n13017), .B(n13013), .Z(n12804) );
  NANDN U13248 ( .A(n13018), .B(n13019), .Z(n13013) );
  XOR U13249 ( .A(n13015), .B(n13020), .Z(n13019) );
  ANDN U13250 ( .B(n13020), .A(n13021), .Z(n13017) );
  XOR U13251 ( .A(n13022), .B(n13009), .Z(n12862) );
  NANDN U13252 ( .A(n13018), .B(n13023), .Z(n13009) );
  XOR U13253 ( .A(n13024), .B(n13012), .Z(n13023) );
  XNOR U13254 ( .A(n13025), .B(n13026), .Z(n13011) );
  XOR U13255 ( .A(n13027), .B(n13028), .Z(n13026) );
  XNOR U13256 ( .A(n13029), .B(n13030), .Z(n13025) );
  XNOR U13257 ( .A(n13031), .B(n13032), .Z(n13030) );
  ANDN U13258 ( .B(n13024), .A(n13028), .Z(n13031) );
  ANDN U13259 ( .B(n13024), .A(n13021), .Z(n13022) );
  XNOR U13260 ( .A(n13027), .B(n13033), .Z(n13021) );
  XOR U13261 ( .A(n13034), .B(n13032), .Z(n13033) );
  NAND U13262 ( .A(n13035), .B(n13036), .Z(n13032) );
  XNOR U13263 ( .A(n13029), .B(n13012), .Z(n13036) );
  IV U13264 ( .A(n13024), .Z(n13029) );
  XNOR U13265 ( .A(n13015), .B(n13028), .Z(n13035) );
  IV U13266 ( .A(n13020), .Z(n13028) );
  XOR U13267 ( .A(n13037), .B(n13038), .Z(n13020) );
  XNOR U13268 ( .A(n13039), .B(n13040), .Z(n13038) );
  XNOR U13269 ( .A(n13041), .B(n13042), .Z(n13037) );
  ANDN U13270 ( .B(n12861), .A(n12914), .Z(n13041) );
  AND U13271 ( .A(n13012), .B(n13015), .Z(n13034) );
  XNOR U13272 ( .A(n13012), .B(n13015), .Z(n13027) );
  XNOR U13273 ( .A(n13043), .B(n13044), .Z(n13015) );
  XNOR U13274 ( .A(n13045), .B(n13040), .Z(n13044) );
  XOR U13275 ( .A(n13046), .B(n13047), .Z(n13043) );
  XNOR U13276 ( .A(n13048), .B(n13042), .Z(n13047) );
  OR U13277 ( .A(n12913), .B(n13002), .Z(n13042) );
  XNOR U13278 ( .A(n12861), .B(n13049), .Z(n13002) );
  XNOR U13279 ( .A(n12914), .B(n12810), .Z(n12913) );
  ANDN U13280 ( .B(n13050), .A(n13001), .Z(n13048) );
  XNOR U13281 ( .A(n13051), .B(n13052), .Z(n13012) );
  XNOR U13282 ( .A(n13040), .B(n13053), .Z(n13052) );
  XOR U13283 ( .A(n12935), .B(n13046), .Z(n13053) );
  XNOR U13284 ( .A(n12861), .B(n12914), .Z(n13040) );
  XOR U13285 ( .A(n12803), .B(n13054), .Z(n13051) );
  XNOR U13286 ( .A(n13055), .B(n13056), .Z(n13054) );
  ANDN U13287 ( .B(n13057), .A(n13006), .Z(n13055) );
  XNOR U13288 ( .A(n13058), .B(n13059), .Z(n13024) );
  XNOR U13289 ( .A(n13045), .B(n13060), .Z(n13059) );
  XNOR U13290 ( .A(n12942), .B(n13039), .Z(n13060) );
  XOR U13291 ( .A(n13046), .B(n13061), .Z(n13039) );
  XNOR U13292 ( .A(n13062), .B(n13063), .Z(n13061) );
  NAND U13293 ( .A(n12868), .B(n12939), .Z(n13063) );
  XNOR U13294 ( .A(n13064), .B(n13062), .Z(n13046) );
  NANDN U13295 ( .A(n13008), .B(n12948), .Z(n13062) );
  XOR U13296 ( .A(n12949), .B(n12939), .Z(n12948) );
  XNOR U13297 ( .A(n13057), .B(n12810), .Z(n12939) );
  XOR U13298 ( .A(n13016), .B(n12868), .Z(n13008) );
  XNOR U13299 ( .A(n13006), .B(n13049), .Z(n12868) );
  ANDN U13300 ( .B(n12949), .A(n13016), .Z(n13064) );
  XOR U13301 ( .A(n12803), .B(n12861), .Z(n13016) );
  XNOR U13302 ( .A(n13065), .B(n13066), .Z(n12861) );
  XNOR U13303 ( .A(n13067), .B(n13068), .Z(n13066) );
  XOR U13304 ( .A(n13049), .B(n13050), .Z(n13045) );
  IV U13305 ( .A(n12810), .Z(n13050) );
  XOR U13306 ( .A(n13070), .B(n13071), .Z(n12810) );
  XNOR U13307 ( .A(n13072), .B(n13068), .Z(n13071) );
  IV U13308 ( .A(n13001), .Z(n13049) );
  XOR U13309 ( .A(n13068), .B(n13073), .Z(n13001) );
  XNOR U13310 ( .A(n13074), .B(n13075), .Z(n13058) );
  XNOR U13311 ( .A(n13076), .B(n13056), .Z(n13075) );
  OR U13312 ( .A(n12945), .B(n13005), .Z(n13056) );
  XNOR U13313 ( .A(n12803), .B(n13006), .Z(n13005) );
  IV U13314 ( .A(n13074), .Z(n13006) );
  XOR U13315 ( .A(n12935), .B(n13057), .Z(n12945) );
  IV U13316 ( .A(n12942), .Z(n13057) );
  XOR U13317 ( .A(n13069), .B(n13077), .Z(n12942) );
  XNOR U13318 ( .A(n13072), .B(n13065), .Z(n13077) );
  XOR U13319 ( .A(n13078), .B(n13079), .Z(n13065) );
  XOR U13320 ( .A(n13080), .B(n12468), .Z(n13079) );
  XNOR U13321 ( .A(key[706]), .B(n12487), .Z(n13078) );
  IV U13322 ( .A(n12914), .Z(n13069) );
  XOR U13323 ( .A(n13070), .B(n13081), .Z(n12914) );
  XOR U13324 ( .A(n13068), .B(n13082), .Z(n13081) );
  NOR U13325 ( .A(n12935), .B(n12803), .Z(n13076) );
  XOR U13326 ( .A(n13070), .B(n13083), .Z(n12935) );
  XOR U13327 ( .A(n13068), .B(n13084), .Z(n13083) );
  XOR U13328 ( .A(n13085), .B(n13086), .Z(n13068) );
  XNOR U13329 ( .A(n12477), .B(n12456), .Z(n13086) );
  XOR U13330 ( .A(n13087), .B(n13088), .Z(n12477) );
  XNOR U13331 ( .A(n13089), .B(n13090), .Z(n13085) );
  XOR U13332 ( .A(key[710]), .B(n12803), .Z(n13090) );
  IV U13333 ( .A(n13073), .Z(n13070) );
  XOR U13334 ( .A(n13091), .B(n13092), .Z(n13073) );
  XOR U13335 ( .A(n12455), .B(n13093), .Z(n13092) );
  XOR U13336 ( .A(n13094), .B(n13095), .Z(n12455) );
  XOR U13337 ( .A(key[709]), .B(n13096), .Z(n13091) );
  XOR U13338 ( .A(n13097), .B(n13098), .Z(n13074) );
  XNOR U13339 ( .A(n13084), .B(n13082), .Z(n13098) );
  XNOR U13340 ( .A(n13099), .B(n13100), .Z(n13082) );
  XNOR U13341 ( .A(n13088), .B(n12462), .Z(n13100) );
  XNOR U13342 ( .A(n13101), .B(n13102), .Z(n12462) );
  XNOR U13343 ( .A(n13103), .B(n13104), .Z(n13088) );
  XOR U13344 ( .A(key[711]), .B(n13105), .Z(n13099) );
  XNOR U13345 ( .A(n13106), .B(n13107), .Z(n13084) );
  XNOR U13346 ( .A(n12447), .B(n12445), .Z(n13107) );
  XNOR U13347 ( .A(n13108), .B(n13109), .Z(n12445) );
  XNOR U13348 ( .A(n13110), .B(n13096), .Z(n12447) );
  XNOR U13349 ( .A(n13111), .B(n13112), .Z(n13106) );
  XOR U13350 ( .A(key[708]), .B(n13113), .Z(n13112) );
  XNOR U13351 ( .A(n12803), .B(n13067), .Z(n13097) );
  XOR U13352 ( .A(n13114), .B(n13115), .Z(n13067) );
  XNOR U13353 ( .A(n12490), .B(n13116), .Z(n13115) );
  XNOR U13354 ( .A(n13072), .B(n12492), .Z(n13116) );
  XNOR U13355 ( .A(n13110), .B(n13113), .Z(n12492) );
  XOR U13356 ( .A(n13117), .B(n13118), .Z(n13072) );
  XNOR U13357 ( .A(n13119), .B(n13120), .Z(n13118) );
  XOR U13358 ( .A(key[705]), .B(n13121), .Z(n13117) );
  XNOR U13359 ( .A(n12469), .B(n13122), .Z(n13114) );
  XNOR U13360 ( .A(key[707]), .B(n13123), .Z(n13122) );
  XNOR U13361 ( .A(n13124), .B(n13125), .Z(n12803) );
  XNOR U13362 ( .A(n13126), .B(n12463), .Z(n13125) );
  XNOR U13363 ( .A(key[704]), .B(n13127), .Z(n13124) );
  IV U13364 ( .A(n9306), .Z(n12762) );
  XOR U13365 ( .A(n12845), .B(n12790), .Z(n9306) );
  XNOR U13366 ( .A(n12851), .B(n13128), .Z(n12790) );
  XNOR U13367 ( .A(n12848), .B(n13129), .Z(n13128) );
  NANDN U13368 ( .A(n13130), .B(n12823), .Z(n13129) );
  NANDN U13369 ( .A(n13131), .B(n12904), .Z(n12848) );
  XNOR U13370 ( .A(n12850), .B(n12823), .Z(n12904) );
  IV U13371 ( .A(n12952), .Z(n12845) );
  XOR U13372 ( .A(n13133), .B(n12815), .Z(n13132) );
  OR U13373 ( .A(n12961), .B(n13134), .Z(n12815) );
  XNOR U13374 ( .A(n12818), .B(n12957), .Z(n12961) );
  ANDN U13375 ( .B(n12957), .A(n13135), .Z(n13133) );
  XNOR U13376 ( .A(n13136), .B(n12853), .Z(n12851) );
  OR U13377 ( .A(n12969), .B(n13137), .Z(n12853) );
  XNOR U13378 ( .A(n12971), .B(n12967), .Z(n12969) );
  IV U13379 ( .A(n12855), .Z(n12967) );
  XNOR U13380 ( .A(n12957), .B(n12823), .Z(n12855) );
  XOR U13381 ( .A(n13138), .B(n13139), .Z(n12823) );
  NANDN U13382 ( .A(n13140), .B(n13141), .Z(n13139) );
  XOR U13383 ( .A(n13142), .B(n13143), .Z(n12957) );
  NANDN U13384 ( .A(n13140), .B(n13144), .Z(n13143) );
  AND U13385 ( .A(n13145), .B(n12971), .Z(n13136) );
  XNOR U13386 ( .A(n12850), .B(n12818), .Z(n12971) );
  XNOR U13387 ( .A(n13146), .B(n13142), .Z(n12818) );
  NANDN U13388 ( .A(n13147), .B(n13148), .Z(n13142) );
  XOR U13389 ( .A(n13144), .B(n13149), .Z(n13148) );
  ANDN U13390 ( .B(n13149), .A(n13150), .Z(n13146) );
  NANDN U13391 ( .A(n13147), .B(n13152), .Z(n13138) );
  XOR U13392 ( .A(n13153), .B(n13141), .Z(n13152) );
  XNOR U13393 ( .A(n13154), .B(n13155), .Z(n13140) );
  XOR U13394 ( .A(n13156), .B(n13157), .Z(n13155) );
  XNOR U13395 ( .A(n13158), .B(n13159), .Z(n13154) );
  XNOR U13396 ( .A(n13160), .B(n13161), .Z(n13159) );
  ANDN U13397 ( .B(n13153), .A(n13157), .Z(n13160) );
  ANDN U13398 ( .B(n13153), .A(n13150), .Z(n13151) );
  XNOR U13399 ( .A(n13156), .B(n13162), .Z(n13150) );
  XOR U13400 ( .A(n13163), .B(n13161), .Z(n13162) );
  NAND U13401 ( .A(n13164), .B(n13165), .Z(n13161) );
  XNOR U13402 ( .A(n13158), .B(n13141), .Z(n13165) );
  IV U13403 ( .A(n13153), .Z(n13158) );
  XNOR U13404 ( .A(n13144), .B(n13157), .Z(n13164) );
  IV U13405 ( .A(n13149), .Z(n13157) );
  XOR U13406 ( .A(n13166), .B(n13167), .Z(n13149) );
  XNOR U13407 ( .A(n13168), .B(n13169), .Z(n13167) );
  XNOR U13408 ( .A(n13170), .B(n13171), .Z(n13166) );
  ANDN U13409 ( .B(n12849), .A(n12905), .Z(n13170) );
  AND U13410 ( .A(n13141), .B(n13144), .Z(n13163) );
  XNOR U13411 ( .A(n13141), .B(n13144), .Z(n13156) );
  XNOR U13412 ( .A(n13172), .B(n13173), .Z(n13144) );
  XNOR U13413 ( .A(n13174), .B(n13169), .Z(n13173) );
  XOR U13414 ( .A(n13175), .B(n13176), .Z(n13172) );
  XNOR U13415 ( .A(n13177), .B(n13171), .Z(n13176) );
  OR U13416 ( .A(n12903), .B(n13131), .Z(n13171) );
  XNOR U13417 ( .A(n12849), .B(n13208), .Z(n13131) );
  XNOR U13418 ( .A(n12905), .B(n12824), .Z(n12903) );
  ANDN U13419 ( .B(n13178), .A(n13130), .Z(n13177) );
  XNOR U13420 ( .A(n13179), .B(n13180), .Z(n13141) );
  XNOR U13421 ( .A(n13169), .B(n13181), .Z(n13180) );
  XNOR U13422 ( .A(n12960), .B(n13175), .Z(n13181) );
  XNOR U13423 ( .A(n12905), .B(n12849), .Z(n13169) );
  XOR U13424 ( .A(n12817), .B(n13182), .Z(n13179) );
  XNOR U13425 ( .A(n13183), .B(n13184), .Z(n13182) );
  ANDN U13426 ( .B(n13185), .A(n13135), .Z(n13183) );
  XNOR U13427 ( .A(n13186), .B(n13187), .Z(n13153) );
  XNOR U13428 ( .A(n13174), .B(n13188), .Z(n13187) );
  XNOR U13429 ( .A(n13189), .B(n13168), .Z(n13188) );
  XOR U13430 ( .A(n13175), .B(n13190), .Z(n13168) );
  XNOR U13431 ( .A(n13191), .B(n13192), .Z(n13190) );
  NANDN U13432 ( .A(n12966), .B(n12856), .Z(n13192) );
  XNOR U13433 ( .A(n13193), .B(n13191), .Z(n13175) );
  OR U13434 ( .A(n13137), .B(n12970), .Z(n13191) );
  XOR U13435 ( .A(n13194), .B(n12966), .Z(n12970) );
  XNOR U13436 ( .A(n13178), .B(n13185), .Z(n12966) );
  IV U13437 ( .A(n12824), .Z(n13178) );
  XNOR U13438 ( .A(n13145), .B(n12856), .Z(n13137) );
  XNOR U13439 ( .A(n13135), .B(n13208), .Z(n12856) );
  ANDN U13440 ( .B(n13145), .A(n12972), .Z(n13193) );
  IV U13441 ( .A(n13194), .Z(n12972) );
  XOR U13442 ( .A(n13195), .B(n12960), .Z(n13194) );
  XOR U13443 ( .A(n12824), .B(n13130), .Z(n13174) );
  XOR U13444 ( .A(n13196), .B(n13197), .Z(n13130) );
  XOR U13445 ( .A(n13198), .B(n13199), .Z(n12824) );
  XOR U13446 ( .A(n13200), .B(n13197), .Z(n13199) );
  XNOR U13447 ( .A(n12956), .B(n13201), .Z(n13186) );
  XNOR U13448 ( .A(n13202), .B(n13184), .Z(n13201) );
  OR U13449 ( .A(n12962), .B(n13134), .Z(n13184) );
  XNOR U13450 ( .A(n12817), .B(n13135), .Z(n13134) );
  IV U13451 ( .A(n13189), .Z(n13135) );
  XOR U13452 ( .A(n13203), .B(n13204), .Z(n13189) );
  XNOR U13453 ( .A(n13205), .B(n13206), .Z(n13204) );
  XNOR U13454 ( .A(n12817), .B(n13207), .Z(n13203) );
  XNOR U13455 ( .A(n12960), .B(n13185), .Z(n12962) );
  IV U13456 ( .A(n12956), .Z(n13185) );
  ANDN U13457 ( .B(n12960), .A(n12817), .Z(n13202) );
  XOR U13458 ( .A(n13205), .B(n13208), .Z(n12960) );
  XOR U13459 ( .A(n13209), .B(n13210), .Z(n13205) );
  XOR U13460 ( .A(n13211), .B(n13212), .Z(n13210) );
  XNOR U13461 ( .A(n13213), .B(n13214), .Z(n13209) );
  XNOR U13462 ( .A(key[700]), .B(n12587), .Z(n13214) );
  XOR U13463 ( .A(n13215), .B(n13216), .Z(n12587) );
  XNOR U13464 ( .A(n13217), .B(n13218), .Z(n12956) );
  XOR U13465 ( .A(n12905), .B(n13198), .Z(n13218) );
  IV U13466 ( .A(n13195), .Z(n12905) );
  XOR U13467 ( .A(n13207), .B(n13208), .Z(n13195) );
  XNOR U13468 ( .A(n13196), .B(n13197), .Z(n13208) );
  IV U13469 ( .A(n13200), .Z(n13196) );
  XNOR U13470 ( .A(n13219), .B(n13220), .Z(n13200) );
  XOR U13471 ( .A(n13221), .B(n13222), .Z(n13220) );
  XOR U13472 ( .A(n13223), .B(n13224), .Z(n13219) );
  XNOR U13473 ( .A(key[701]), .B(n13225), .Z(n13224) );
  XOR U13474 ( .A(n13226), .B(n13227), .Z(n13207) );
  XOR U13475 ( .A(n13228), .B(n13229), .Z(n13227) );
  XNOR U13476 ( .A(key[703]), .B(n13230), .Z(n13226) );
  XNOR U13477 ( .A(n12817), .B(n12849), .Z(n13145) );
  XNOR U13478 ( .A(n13206), .B(n13231), .Z(n12849) );
  XNOR U13479 ( .A(n13197), .B(n13217), .Z(n13231) );
  XOR U13480 ( .A(n13232), .B(n13233), .Z(n13217) );
  XOR U13481 ( .A(n13234), .B(n13235), .Z(n13233) );
  XOR U13482 ( .A(n12623), .B(n13236), .Z(n13232) );
  XOR U13483 ( .A(key[698]), .B(n13237), .Z(n13236) );
  XOR U13484 ( .A(n13238), .B(n13239), .Z(n13197) );
  XOR U13485 ( .A(n12615), .B(n13240), .Z(n13239) );
  XNOR U13486 ( .A(n12598), .B(n13241), .Z(n12615) );
  XOR U13487 ( .A(n12817), .B(n13242), .Z(n13238) );
  XNOR U13488 ( .A(key[702]), .B(n13243), .Z(n13242) );
  XOR U13489 ( .A(n13244), .B(n13245), .Z(n13206) );
  XNOR U13490 ( .A(n12631), .B(n13246), .Z(n13245) );
  XNOR U13491 ( .A(n13247), .B(n13248), .Z(n13246) );
  XNOR U13492 ( .A(n12628), .B(n13249), .Z(n13244) );
  XOR U13493 ( .A(key[699]), .B(n13198), .Z(n13249) );
  XNOR U13494 ( .A(n13250), .B(n13251), .Z(n13198) );
  XNOR U13495 ( .A(n13252), .B(n12611), .Z(n13251) );
  XOR U13496 ( .A(n13253), .B(n13254), .Z(n13250) );
  XNOR U13497 ( .A(key[697]), .B(n13255), .Z(n13254) );
  XNOR U13498 ( .A(n12598), .B(n13256), .Z(n12628) );
  XNOR U13499 ( .A(n13257), .B(n13258), .Z(n12817) );
  XOR U13500 ( .A(n13259), .B(n13260), .Z(n13258) );
  XOR U13501 ( .A(n12612), .B(n13261), .Z(n13257) );
  XNOR U13502 ( .A(key[696]), .B(n12598), .Z(n13261) );
  IV U13503 ( .A(n13216), .Z(n12598) );
  XOR U13504 ( .A(n12917), .B(n12878), .Z(n10206) );
  XOR U13505 ( .A(n12923), .B(n13262), .Z(n12917) );
  XOR U13506 ( .A(n13263), .B(n12874), .Z(n13262) );
  OR U13507 ( .A(n13264), .B(n13265), .Z(n12874) );
  NOR U13508 ( .A(n13266), .B(n13267), .Z(n13263) );
  XOR U13509 ( .A(key[818]), .B(n11155), .Z(n12996) );
  XOR U13510 ( .A(n10164), .B(n9263), .Z(n11155) );
  XOR U13511 ( .A(n13268), .B(n13269), .Z(n9263) );
  XNOR U13512 ( .A(n12886), .B(n12836), .Z(n13269) );
  XNOR U13513 ( .A(n13270), .B(n13271), .Z(n12836) );
  XNOR U13514 ( .A(n13272), .B(n12770), .Z(n13271) );
  ANDN U13515 ( .B(n13273), .A(n13274), .Z(n12770) );
  NOR U13516 ( .A(n13275), .B(n12989), .Z(n13272) );
  IV U13517 ( .A(n12842), .Z(n12886) );
  XOR U13518 ( .A(n12978), .B(n13276), .Z(n12842) );
  XOR U13519 ( .A(n12987), .B(n13277), .Z(n13276) );
  NANDN U13520 ( .A(n13278), .B(n12772), .Z(n13277) );
  XNOR U13521 ( .A(n12989), .B(n12772), .Z(n13273) );
  IV U13522 ( .A(n12990), .Z(n12978) );
  XNOR U13523 ( .A(n13280), .B(n12992), .Z(n12990) );
  OR U13524 ( .A(n13281), .B(n13282), .Z(n12992) );
  ANDN U13525 ( .B(n13283), .A(n13284), .Z(n13280) );
  XNOR U13526 ( .A(n12844), .B(n12894), .Z(n13268) );
  XNOR U13527 ( .A(n12766), .B(n13285), .Z(n12894) );
  XNOR U13528 ( .A(n13286), .B(n13287), .Z(n13285) );
  NANDN U13529 ( .A(n13288), .B(n12983), .Z(n13287) );
  XNOR U13530 ( .A(n13286), .B(n13290), .Z(n13289) );
  NANDN U13531 ( .A(n13291), .B(n12892), .Z(n13290) );
  OR U13532 ( .A(n12982), .B(n13292), .Z(n13286) );
  XNOR U13533 ( .A(n12892), .B(n12983), .Z(n12982) );
  XNOR U13534 ( .A(n12766), .B(n13293), .Z(n13270) );
  XNOR U13535 ( .A(n13294), .B(n13295), .Z(n13293) );
  NAND U13536 ( .A(n13296), .B(n12994), .Z(n13295) );
  XOR U13537 ( .A(n13297), .B(n13294), .Z(n12766) );
  NANDN U13538 ( .A(n13281), .B(n13298), .Z(n13294) );
  XNOR U13539 ( .A(n13283), .B(n12994), .Z(n13281) );
  XOR U13540 ( .A(n12983), .B(n12772), .Z(n12994) );
  XOR U13541 ( .A(n13299), .B(n13300), .Z(n12772) );
  NANDN U13542 ( .A(n13301), .B(n13302), .Z(n13300) );
  XOR U13543 ( .A(n13303), .B(n13304), .Z(n12983) );
  NANDN U13544 ( .A(n13301), .B(n13305), .Z(n13304) );
  IV U13545 ( .A(n13306), .Z(n13283) );
  ANDN U13546 ( .B(n13307), .A(n13306), .Z(n13297) );
  XOR U13547 ( .A(n12989), .B(n12892), .Z(n13306) );
  XNOR U13548 ( .A(n13308), .B(n13303), .Z(n12892) );
  NANDN U13549 ( .A(n13309), .B(n13310), .Z(n13303) );
  XOR U13550 ( .A(n13305), .B(n13311), .Z(n13310) );
  ANDN U13551 ( .B(n13311), .A(n13312), .Z(n13308) );
  XOR U13552 ( .A(n13313), .B(n13299), .Z(n12989) );
  NANDN U13553 ( .A(n13309), .B(n13314), .Z(n13299) );
  XOR U13554 ( .A(n13315), .B(n13302), .Z(n13314) );
  XNOR U13555 ( .A(n13316), .B(n13317), .Z(n13301) );
  XOR U13556 ( .A(n13318), .B(n13319), .Z(n13317) );
  XNOR U13557 ( .A(n13320), .B(n13321), .Z(n13316) );
  XNOR U13558 ( .A(n13322), .B(n13323), .Z(n13321) );
  ANDN U13559 ( .B(n13315), .A(n13319), .Z(n13322) );
  ANDN U13560 ( .B(n13315), .A(n13312), .Z(n13313) );
  XNOR U13561 ( .A(n13318), .B(n13324), .Z(n13312) );
  XOR U13562 ( .A(n13325), .B(n13323), .Z(n13324) );
  NAND U13563 ( .A(n13326), .B(n13327), .Z(n13323) );
  XNOR U13564 ( .A(n13320), .B(n13302), .Z(n13327) );
  IV U13565 ( .A(n13315), .Z(n13320) );
  XNOR U13566 ( .A(n13305), .B(n13319), .Z(n13326) );
  IV U13567 ( .A(n13311), .Z(n13319) );
  XOR U13568 ( .A(n13328), .B(n13329), .Z(n13311) );
  XNOR U13569 ( .A(n13330), .B(n13331), .Z(n13329) );
  XNOR U13570 ( .A(n13332), .B(n13333), .Z(n13328) );
  ANDN U13571 ( .B(n12988), .A(n13275), .Z(n13332) );
  AND U13572 ( .A(n13302), .B(n13305), .Z(n13325) );
  XNOR U13573 ( .A(n13302), .B(n13305), .Z(n13318) );
  XNOR U13574 ( .A(n13334), .B(n13335), .Z(n13305) );
  XNOR U13575 ( .A(n13336), .B(n13331), .Z(n13335) );
  XOR U13576 ( .A(n13337), .B(n13338), .Z(n13334) );
  XNOR U13577 ( .A(n13339), .B(n13333), .Z(n13338) );
  OR U13578 ( .A(n13274), .B(n13279), .Z(n13333) );
  XNOR U13579 ( .A(n12988), .B(n13340), .Z(n13279) );
  XNOR U13580 ( .A(n13275), .B(n12773), .Z(n13274) );
  ANDN U13581 ( .B(n13341), .A(n13278), .Z(n13339) );
  XNOR U13582 ( .A(n13342), .B(n13343), .Z(n13302) );
  XNOR U13583 ( .A(n13331), .B(n13344), .Z(n13343) );
  XOR U13584 ( .A(n13291), .B(n13337), .Z(n13344) );
  XNOR U13585 ( .A(n12988), .B(n13275), .Z(n13331) );
  XOR U13586 ( .A(n12891), .B(n13345), .Z(n13342) );
  XNOR U13587 ( .A(n13346), .B(n13347), .Z(n13345) );
  ANDN U13588 ( .B(n13348), .A(n12984), .Z(n13346) );
  XNOR U13589 ( .A(n13349), .B(n13350), .Z(n13315) );
  XNOR U13590 ( .A(n13336), .B(n13351), .Z(n13350) );
  XNOR U13591 ( .A(n13288), .B(n13330), .Z(n13351) );
  XOR U13592 ( .A(n13337), .B(n13352), .Z(n13330) );
  XNOR U13593 ( .A(n13353), .B(n13354), .Z(n13352) );
  NAND U13594 ( .A(n12995), .B(n13296), .Z(n13354) );
  XNOR U13595 ( .A(n13355), .B(n13353), .Z(n13337) );
  NANDN U13596 ( .A(n13282), .B(n13298), .Z(n13353) );
  XOR U13597 ( .A(n13307), .B(n13296), .Z(n13298) );
  XNOR U13598 ( .A(n13348), .B(n12773), .Z(n13296) );
  XOR U13599 ( .A(n13284), .B(n12995), .Z(n13282) );
  XNOR U13600 ( .A(n12984), .B(n13340), .Z(n12995) );
  ANDN U13601 ( .B(n13307), .A(n13284), .Z(n13355) );
  XOR U13602 ( .A(n12891), .B(n12988), .Z(n13284) );
  XNOR U13603 ( .A(n13356), .B(n13357), .Z(n12988) );
  XNOR U13604 ( .A(n13358), .B(n13359), .Z(n13357) );
  XOR U13605 ( .A(n13340), .B(n13341), .Z(n13336) );
  IV U13606 ( .A(n12773), .Z(n13341) );
  XOR U13607 ( .A(n13360), .B(n13361), .Z(n12773) );
  XNOR U13608 ( .A(n13362), .B(n13359), .Z(n13361) );
  IV U13609 ( .A(n13278), .Z(n13340) );
  XOR U13610 ( .A(n13359), .B(n13363), .Z(n13278) );
  XNOR U13611 ( .A(n13364), .B(n13365), .Z(n13349) );
  XNOR U13612 ( .A(n13366), .B(n13347), .Z(n13365) );
  OR U13613 ( .A(n13292), .B(n12981), .Z(n13347) );
  XNOR U13614 ( .A(n12891), .B(n12984), .Z(n12981) );
  IV U13615 ( .A(n13364), .Z(n12984) );
  XOR U13616 ( .A(n13291), .B(n13348), .Z(n13292) );
  IV U13617 ( .A(n13288), .Z(n13348) );
  XOR U13618 ( .A(n13367), .B(n13368), .Z(n13288) );
  XNOR U13619 ( .A(n13362), .B(n13356), .Z(n13368) );
  XOR U13620 ( .A(n13369), .B(n13370), .Z(n13356) );
  XNOR U13621 ( .A(n12297), .B(n13371), .Z(n13370) );
  XNOR U13622 ( .A(key[658]), .B(n12288), .Z(n13369) );
  NOR U13623 ( .A(n13291), .B(n12891), .Z(n13366) );
  XOR U13624 ( .A(n13372), .B(n13373), .Z(n13364) );
  XNOR U13625 ( .A(n13374), .B(n13375), .Z(n13373) );
  XNOR U13626 ( .A(n12891), .B(n13358), .Z(n13372) );
  XOR U13627 ( .A(n13376), .B(n13377), .Z(n13358) );
  XNOR U13628 ( .A(n12291), .B(n13378), .Z(n13377) );
  XOR U13629 ( .A(n13362), .B(n13379), .Z(n13378) );
  XOR U13630 ( .A(n13380), .B(n13381), .Z(n13362) );
  XOR U13631 ( .A(n13382), .B(n12286), .Z(n13381) );
  XOR U13632 ( .A(key[657]), .B(n13383), .Z(n13380) );
  XNOR U13633 ( .A(n12300), .B(n13384), .Z(n13376) );
  XNOR U13634 ( .A(key[659]), .B(n12293), .Z(n13384) );
  XNOR U13635 ( .A(n13385), .B(n13386), .Z(n12293) );
  IV U13636 ( .A(n13275), .Z(n13367) );
  XOR U13637 ( .A(n13360), .B(n13387), .Z(n13275) );
  XOR U13638 ( .A(n13359), .B(n13375), .Z(n13387) );
  XNOR U13639 ( .A(n13388), .B(n13389), .Z(n13375) );
  XOR U13640 ( .A(n13390), .B(n12269), .Z(n13389) );
  XNOR U13641 ( .A(n13391), .B(n13392), .Z(n12269) );
  XNOR U13642 ( .A(key[663]), .B(n13393), .Z(n13388) );
  XOR U13643 ( .A(n13360), .B(n13394), .Z(n13291) );
  XOR U13644 ( .A(n13359), .B(n13374), .Z(n13394) );
  XNOR U13645 ( .A(n13395), .B(n13396), .Z(n13374) );
  XOR U13646 ( .A(n12257), .B(n13397), .Z(n13396) );
  XOR U13647 ( .A(n13398), .B(n13399), .Z(n12257) );
  XNOR U13648 ( .A(n13400), .B(n13401), .Z(n13399) );
  XNOR U13649 ( .A(n13402), .B(n13403), .Z(n13398) );
  XNOR U13650 ( .A(key[660]), .B(n13386), .Z(n13395) );
  XOR U13651 ( .A(n13404), .B(n13405), .Z(n13359) );
  XNOR U13652 ( .A(n13406), .B(n12306), .Z(n13405) );
  XNOR U13653 ( .A(n13390), .B(n13407), .Z(n12306) );
  XNOR U13654 ( .A(n13402), .B(n13408), .Z(n13390) );
  XNOR U13655 ( .A(n12277), .B(n13409), .Z(n13404) );
  XOR U13656 ( .A(key[662]), .B(n12891), .Z(n13409) );
  XNOR U13657 ( .A(n13410), .B(n13411), .Z(n12891) );
  XOR U13658 ( .A(n13412), .B(n12270), .Z(n13411) );
  XOR U13659 ( .A(key[656]), .B(n13413), .Z(n13410) );
  IV U13660 ( .A(n13363), .Z(n13360) );
  XOR U13661 ( .A(n13414), .B(n13415), .Z(n13363) );
  XOR U13662 ( .A(n12274), .B(n13416), .Z(n13415) );
  XOR U13663 ( .A(n13417), .B(n13418), .Z(n12274) );
  XNOR U13664 ( .A(key[661]), .B(n13403), .Z(n13414) );
  XOR U13665 ( .A(n13419), .B(n13420), .Z(n10164) );
  XOR U13666 ( .A(n12975), .B(n12883), .Z(n13420) );
  XNOR U13667 ( .A(n13421), .B(n13422), .Z(n12883) );
  XNOR U13668 ( .A(n13423), .B(n12831), .Z(n13422) );
  ANDN U13669 ( .B(n13424), .A(n13425), .Z(n12831) );
  NOR U13670 ( .A(n13426), .B(n12922), .Z(n13423) );
  XOR U13671 ( .A(n12827), .B(n13427), .Z(n12975) );
  XNOR U13672 ( .A(n13428), .B(n13429), .Z(n13427) );
  NANDN U13673 ( .A(n13267), .B(n13430), .Z(n13429) );
  XNOR U13674 ( .A(n12878), .B(n12974), .Z(n13419) );
  IV U13675 ( .A(n12879), .Z(n12974) );
  XOR U13676 ( .A(n13421), .B(n13431), .Z(n12879) );
  XNOR U13677 ( .A(n13428), .B(n13432), .Z(n13431) );
  OR U13678 ( .A(n12876), .B(n13433), .Z(n13432) );
  OR U13679 ( .A(n13265), .B(n13434), .Z(n13428) );
  XNOR U13680 ( .A(n12876), .B(n13267), .Z(n13265) );
  XNOR U13681 ( .A(n12827), .B(n13435), .Z(n13421) );
  XNOR U13682 ( .A(n13436), .B(n13437), .Z(n13435) );
  NAND U13683 ( .A(n13438), .B(n12927), .Z(n13437) );
  XOR U13684 ( .A(n13439), .B(n13436), .Z(n12827) );
  NANDN U13685 ( .A(n13440), .B(n13441), .Z(n13436) );
  AND U13686 ( .A(n13442), .B(n13443), .Z(n13439) );
  XOR U13687 ( .A(n12923), .B(n13444), .Z(n12878) );
  XOR U13688 ( .A(n12920), .B(n13445), .Z(n13444) );
  NAND U13689 ( .A(n13446), .B(n12833), .Z(n13445) );
  XNOR U13690 ( .A(n12922), .B(n12833), .Z(n13424) );
  XOR U13691 ( .A(n13448), .B(n12925), .Z(n12923) );
  OR U13692 ( .A(n13440), .B(n13449), .Z(n12925) );
  XNOR U13693 ( .A(n13442), .B(n12927), .Z(n13440) );
  XNOR U13694 ( .A(n13267), .B(n12833), .Z(n12927) );
  XOR U13695 ( .A(n13450), .B(n13451), .Z(n12833) );
  NANDN U13696 ( .A(n13452), .B(n13453), .Z(n13451) );
  XNOR U13697 ( .A(n13454), .B(n13455), .Z(n13267) );
  OR U13698 ( .A(n13452), .B(n13456), .Z(n13455) );
  ANDN U13699 ( .B(n13442), .A(n13457), .Z(n13448) );
  XOR U13700 ( .A(n12876), .B(n12922), .Z(n13442) );
  XOR U13701 ( .A(n13458), .B(n13450), .Z(n12922) );
  NANDN U13702 ( .A(n13459), .B(n13460), .Z(n13450) );
  ANDN U13703 ( .B(n13461), .A(n13462), .Z(n13458) );
  NANDN U13704 ( .A(n13459), .B(n13464), .Z(n13454) );
  XOR U13705 ( .A(n13465), .B(n13452), .Z(n13459) );
  XNOR U13706 ( .A(n13466), .B(n13467), .Z(n13452) );
  XOR U13707 ( .A(n13468), .B(n13461), .Z(n13467) );
  XNOR U13708 ( .A(n13469), .B(n13470), .Z(n13466) );
  XNOR U13709 ( .A(n13471), .B(n13472), .Z(n13470) );
  ANDN U13710 ( .B(n13461), .A(n13473), .Z(n13471) );
  IV U13711 ( .A(n13474), .Z(n13461) );
  ANDN U13712 ( .B(n13465), .A(n13473), .Z(n13463) );
  IV U13713 ( .A(n13469), .Z(n13473) );
  IV U13714 ( .A(n13462), .Z(n13465) );
  XNOR U13715 ( .A(n13468), .B(n13475), .Z(n13462) );
  XOR U13716 ( .A(n13476), .B(n13472), .Z(n13475) );
  NAND U13717 ( .A(n13464), .B(n13460), .Z(n13472) );
  XNOR U13718 ( .A(n13453), .B(n13474), .Z(n13460) );
  XOR U13719 ( .A(n13477), .B(n13478), .Z(n13474) );
  XOR U13720 ( .A(n13479), .B(n13480), .Z(n13478) );
  XNOR U13721 ( .A(n13430), .B(n13481), .Z(n13480) );
  XNOR U13722 ( .A(n13482), .B(n13483), .Z(n13477) );
  XNOR U13723 ( .A(n13484), .B(n13485), .Z(n13483) );
  ANDN U13724 ( .B(n13486), .A(n12877), .Z(n13484) );
  XNOR U13725 ( .A(n13469), .B(n13456), .Z(n13464) );
  XOR U13726 ( .A(n13487), .B(n13488), .Z(n13469) );
  XNOR U13727 ( .A(n13489), .B(n13481), .Z(n13488) );
  XOR U13728 ( .A(n13490), .B(n13491), .Z(n13481) );
  XNOR U13729 ( .A(n13492), .B(n13493), .Z(n13491) );
  NAND U13730 ( .A(n12928), .B(n13438), .Z(n13493) );
  XNOR U13731 ( .A(n13494), .B(n13495), .Z(n13487) );
  ANDN U13732 ( .B(n13496), .A(n12921), .Z(n13494) );
  ANDN U13733 ( .B(n13453), .A(n13456), .Z(n13476) );
  XOR U13734 ( .A(n13456), .B(n13453), .Z(n13468) );
  XNOR U13735 ( .A(n13497), .B(n13498), .Z(n13453) );
  XNOR U13736 ( .A(n13490), .B(n13499), .Z(n13498) );
  XOR U13737 ( .A(n13489), .B(n13433), .Z(n13499) );
  XOR U13738 ( .A(n12877), .B(n13500), .Z(n13497) );
  XNOR U13739 ( .A(n13501), .B(n13485), .Z(n13500) );
  OR U13740 ( .A(n13434), .B(n13264), .Z(n13485) );
  XNOR U13741 ( .A(n12877), .B(n13266), .Z(n13264) );
  XOR U13742 ( .A(n13433), .B(n13430), .Z(n13434) );
  ANDN U13743 ( .B(n13430), .A(n13266), .Z(n13501) );
  XOR U13744 ( .A(n13502), .B(n13503), .Z(n13456) );
  XOR U13745 ( .A(n13490), .B(n13479), .Z(n13503) );
  XOR U13746 ( .A(n13446), .B(n12834), .Z(n13479) );
  XOR U13747 ( .A(n13504), .B(n13492), .Z(n13490) );
  NANDN U13748 ( .A(n13449), .B(n13441), .Z(n13492) );
  XOR U13749 ( .A(n13443), .B(n13438), .Z(n13441) );
  XNOR U13750 ( .A(n13496), .B(n13505), .Z(n13430) );
  XNOR U13751 ( .A(n13506), .B(n13507), .Z(n13505) );
  XOR U13752 ( .A(n13457), .B(n12928), .Z(n13449) );
  XNOR U13753 ( .A(n13266), .B(n13446), .Z(n12928) );
  IV U13754 ( .A(n13482), .Z(n13266) );
  XOR U13755 ( .A(n13508), .B(n13509), .Z(n13482) );
  XOR U13756 ( .A(n13510), .B(n13511), .Z(n13509) );
  XNOR U13757 ( .A(n12877), .B(n13512), .Z(n13508) );
  ANDN U13758 ( .B(n13443), .A(n13457), .Z(n13504) );
  XNOR U13759 ( .A(n12877), .B(n12921), .Z(n13457) );
  XOR U13760 ( .A(n13496), .B(n13486), .Z(n13443) );
  IV U13761 ( .A(n13433), .Z(n13486) );
  XOR U13762 ( .A(n13513), .B(n13514), .Z(n13433) );
  XOR U13763 ( .A(n13515), .B(n13511), .Z(n13514) );
  XNOR U13764 ( .A(n13516), .B(n13517), .Z(n13511) );
  XOR U13765 ( .A(n13518), .B(n13519), .Z(n13517) );
  XNOR U13766 ( .A(n12127), .B(n13520), .Z(n13516) );
  XNOR U13767 ( .A(key[748]), .B(n13521), .Z(n13520) );
  XOR U13768 ( .A(n12138), .B(n13522), .Z(n12127) );
  IV U13769 ( .A(n13426), .Z(n13496) );
  XOR U13770 ( .A(n13489), .B(n13523), .Z(n13502) );
  XNOR U13771 ( .A(n13524), .B(n13495), .Z(n13523) );
  OR U13772 ( .A(n13425), .B(n13447), .Z(n13495) );
  XNOR U13773 ( .A(n13525), .B(n13446), .Z(n13447) );
  XNOR U13774 ( .A(n13426), .B(n12834), .Z(n13425) );
  ANDN U13775 ( .B(n13446), .A(n12834), .Z(n13524) );
  XOR U13776 ( .A(n13513), .B(n13526), .Z(n12834) );
  XOR U13777 ( .A(n13506), .B(n13527), .Z(n13526) );
  XOR U13778 ( .A(n13515), .B(n13513), .Z(n13446) );
  XNOR U13779 ( .A(n12921), .B(n13426), .Z(n13489) );
  XOR U13780 ( .A(n13513), .B(n13528), .Z(n13426) );
  XNOR U13781 ( .A(n13515), .B(n13510), .Z(n13528) );
  XOR U13782 ( .A(n13529), .B(n13530), .Z(n13510) );
  XOR U13783 ( .A(n13531), .B(n13532), .Z(n13530) );
  XNOR U13784 ( .A(key[751]), .B(n13533), .Z(n13529) );
  XNOR U13785 ( .A(n13534), .B(n13535), .Z(n13513) );
  XOR U13786 ( .A(n13536), .B(n13537), .Z(n13535) );
  XNOR U13787 ( .A(n13538), .B(n13539), .Z(n13534) );
  XOR U13788 ( .A(key[749]), .B(n13540), .Z(n13539) );
  IV U13789 ( .A(n13525), .Z(n12921) );
  XNOR U13790 ( .A(n13507), .B(n13541), .Z(n13525) );
  XOR U13791 ( .A(n13512), .B(n13527), .Z(n13541) );
  IV U13792 ( .A(n13515), .Z(n13527) );
  XOR U13793 ( .A(n13542), .B(n13543), .Z(n13515) );
  XNOR U13794 ( .A(n13544), .B(n13545), .Z(n13543) );
  XNOR U13795 ( .A(n12173), .B(n13546), .Z(n13542) );
  XOR U13796 ( .A(key[750]), .B(n12877), .Z(n13546) );
  XNOR U13797 ( .A(n13547), .B(n13548), .Z(n12877) );
  XOR U13798 ( .A(n13549), .B(n13550), .Z(n13548) );
  XOR U13799 ( .A(n12170), .B(n13551), .Z(n13547) );
  XNOR U13800 ( .A(key[744]), .B(n13552), .Z(n13551) );
  XNOR U13801 ( .A(n12138), .B(n13553), .Z(n12173) );
  XOR U13802 ( .A(n13554), .B(n13555), .Z(n13512) );
  XNOR U13803 ( .A(n12155), .B(n13556), .Z(n13555) );
  XNOR U13804 ( .A(n13506), .B(n13557), .Z(n13556) );
  XOR U13805 ( .A(n13558), .B(n13559), .Z(n13506) );
  XNOR U13806 ( .A(n12169), .B(n13560), .Z(n13559) );
  XNOR U13807 ( .A(n13561), .B(n13562), .Z(n13558) );
  XOR U13808 ( .A(key[745]), .B(n13563), .Z(n13562) );
  XNOR U13809 ( .A(n12138), .B(n13564), .Z(n12155) );
  IV U13810 ( .A(n13550), .Z(n12138) );
  XNOR U13811 ( .A(n13565), .B(n13566), .Z(n13554) );
  XNOR U13812 ( .A(key[747]), .B(n12162), .Z(n13566) );
  XOR U13813 ( .A(n13567), .B(n13568), .Z(n13507) );
  XOR U13814 ( .A(n13569), .B(n13570), .Z(n13568) );
  XOR U13815 ( .A(n12152), .B(n13571), .Z(n13567) );
  XNOR U13816 ( .A(key[746]), .B(n13572), .Z(n13571) );
  XOR U13817 ( .A(key[976]), .B(n6290), .Z(n11724) );
  XNOR U13818 ( .A(n8355), .B(n8385), .Z(n6290) );
  XOR U13819 ( .A(n11556), .B(n11602), .Z(n8385) );
  XNOR U13820 ( .A(n11596), .B(n13573), .Z(n11602) );
  XNOR U13821 ( .A(n12637), .B(n13574), .Z(n13573) );
  OR U13822 ( .A(n11712), .B(n13575), .Z(n13574) );
  NANDN U13823 ( .A(n13576), .B(n11710), .Z(n12637) );
  XOR U13824 ( .A(n11712), .B(n11607), .Z(n11710) );
  XNOR U13825 ( .A(n12635), .B(n13577), .Z(n11596) );
  XNOR U13826 ( .A(n13578), .B(n13579), .Z(n13577) );
  NAND U13827 ( .A(n12648), .B(n13580), .Z(n13579) );
  IV U13828 ( .A(n11702), .Z(n11556) );
  XNOR U13829 ( .A(n12635), .B(n13581), .Z(n11702) );
  XOR U13830 ( .A(n13582), .B(n11598), .Z(n13581) );
  OR U13831 ( .A(n13583), .B(n12653), .Z(n11598) );
  XNOR U13832 ( .A(n11600), .B(n12651), .Z(n12653) );
  NOR U13833 ( .A(n13584), .B(n12651), .Z(n13582) );
  XOR U13834 ( .A(n13585), .B(n13578), .Z(n12635) );
  OR U13835 ( .A(n12656), .B(n13586), .Z(n13578) );
  XNOR U13836 ( .A(n12658), .B(n12648), .Z(n12656) );
  XOR U13837 ( .A(n12651), .B(n11607), .Z(n12648) );
  XNOR U13838 ( .A(n13587), .B(n13588), .Z(n11607) );
  NANDN U13839 ( .A(n13589), .B(n13590), .Z(n13588) );
  XNOR U13840 ( .A(n13591), .B(n13592), .Z(n12651) );
  OR U13841 ( .A(n13589), .B(n13593), .Z(n13592) );
  ANDN U13842 ( .B(n12658), .A(n13594), .Z(n13585) );
  XOR U13843 ( .A(n11600), .B(n11712), .Z(n12658) );
  XNOR U13844 ( .A(n13587), .B(n13595), .Z(n11712) );
  NANDN U13845 ( .A(n13596), .B(n13597), .Z(n13595) );
  NANDN U13846 ( .A(n13598), .B(n13599), .Z(n13587) );
  OR U13847 ( .A(n13601), .B(n13598), .Z(n13591) );
  XOR U13848 ( .A(n13602), .B(n13589), .Z(n13598) );
  XNOR U13849 ( .A(n13603), .B(n13604), .Z(n13589) );
  XOR U13850 ( .A(n13605), .B(n13597), .Z(n13604) );
  XNOR U13851 ( .A(n13606), .B(n13607), .Z(n13603) );
  XNOR U13852 ( .A(n13608), .B(n13609), .Z(n13607) );
  ANDN U13853 ( .B(n13597), .A(n13610), .Z(n13608) );
  IV U13854 ( .A(n13611), .Z(n13597) );
  ANDN U13855 ( .B(n13602), .A(n13610), .Z(n13600) );
  IV U13856 ( .A(n13596), .Z(n13602) );
  XNOR U13857 ( .A(n13605), .B(n13612), .Z(n13596) );
  XNOR U13858 ( .A(n13609), .B(n13613), .Z(n13612) );
  NANDN U13859 ( .A(n13593), .B(n13590), .Z(n13613) );
  NANDN U13860 ( .A(n13601), .B(n13599), .Z(n13609) );
  XNOR U13861 ( .A(n13590), .B(n13611), .Z(n13599) );
  XOR U13862 ( .A(n13614), .B(n13615), .Z(n13611) );
  XOR U13863 ( .A(n13616), .B(n13617), .Z(n13615) );
  XNOR U13864 ( .A(n12652), .B(n13618), .Z(n13617) );
  XNOR U13865 ( .A(n13619), .B(n13620), .Z(n13614) );
  XNOR U13866 ( .A(n13621), .B(n13622), .Z(n13620) );
  ANDN U13867 ( .B(n12643), .A(n11601), .Z(n13621) );
  XNOR U13868 ( .A(n13610), .B(n13593), .Z(n13601) );
  IV U13869 ( .A(n13606), .Z(n13610) );
  XOR U13870 ( .A(n13623), .B(n13624), .Z(n13606) );
  XNOR U13871 ( .A(n13625), .B(n13618), .Z(n13624) );
  XOR U13872 ( .A(n13626), .B(n13627), .Z(n13618) );
  XNOR U13873 ( .A(n13628), .B(n13629), .Z(n13627) );
  NAND U13874 ( .A(n13580), .B(n12647), .Z(n13629) );
  XNOR U13875 ( .A(n13630), .B(n13631), .Z(n13623) );
  ANDN U13876 ( .B(n13632), .A(n13575), .Z(n13630) );
  XOR U13877 ( .A(n13593), .B(n13590), .Z(n13605) );
  XNOR U13878 ( .A(n13633), .B(n13634), .Z(n13590) );
  XNOR U13879 ( .A(n13626), .B(n13635), .Z(n13634) );
  XNOR U13880 ( .A(n13625), .B(n12643), .Z(n13635) );
  XNOR U13881 ( .A(n13636), .B(n13637), .Z(n13633) );
  XNOR U13882 ( .A(n13638), .B(n13622), .Z(n13637) );
  OR U13883 ( .A(n12654), .B(n13583), .Z(n13622) );
  XNOR U13884 ( .A(n13636), .B(n13619), .Z(n13583) );
  XNOR U13885 ( .A(n12643), .B(n12652), .Z(n12654) );
  ANDN U13886 ( .B(n12652), .A(n13584), .Z(n13638) );
  XOR U13887 ( .A(n13639), .B(n13640), .Z(n13593) );
  XOR U13888 ( .A(n13626), .B(n13616), .Z(n13640) );
  XOR U13889 ( .A(n13641), .B(n11606), .Z(n13616) );
  XOR U13890 ( .A(n13642), .B(n13628), .Z(n13626) );
  NANDN U13891 ( .A(n13586), .B(n12657), .Z(n13628) );
  XOR U13892 ( .A(n12659), .B(n12647), .Z(n12657) );
  XOR U13893 ( .A(n11606), .B(n12652), .Z(n12647) );
  XNOR U13894 ( .A(n13632), .B(n13643), .Z(n12652) );
  XOR U13895 ( .A(n13644), .B(n13645), .Z(n13643) );
  XOR U13896 ( .A(n13594), .B(n13580), .Z(n13586) );
  XNOR U13897 ( .A(n13584), .B(n12639), .Z(n13580) );
  IV U13898 ( .A(n13619), .Z(n13584) );
  XOR U13899 ( .A(n13646), .B(n13647), .Z(n13619) );
  XOR U13900 ( .A(n13648), .B(n13649), .Z(n13647) );
  XOR U13901 ( .A(n13636), .B(n13650), .Z(n13646) );
  ANDN U13902 ( .B(n12659), .A(n13594), .Z(n13642) );
  XNOR U13903 ( .A(n13636), .B(n13651), .Z(n13594) );
  XOR U13904 ( .A(n13632), .B(n12643), .Z(n12659) );
  XNOR U13905 ( .A(n13652), .B(n13653), .Z(n12643) );
  XOR U13906 ( .A(n13654), .B(n13649), .Z(n13653) );
  XNOR U13907 ( .A(n13655), .B(n13656), .Z(n13649) );
  XOR U13908 ( .A(n11243), .B(n10037), .Z(n13656) );
  XOR U13909 ( .A(n13658), .B(n11281), .Z(n11243) );
  XNOR U13910 ( .A(key[780]), .B(n9129), .Z(n13655) );
  XOR U13911 ( .A(n13659), .B(n13660), .Z(n9129) );
  XNOR U13912 ( .A(n11245), .B(n11277), .Z(n13660) );
  XOR U13913 ( .A(n13661), .B(n10055), .Z(n11277) );
  XOR U13914 ( .A(n9135), .B(n13662), .Z(n13659) );
  XOR U13915 ( .A(n13663), .B(n13664), .Z(n9135) );
  XNOR U13916 ( .A(n13665), .B(n13666), .Z(n13664) );
  XNOR U13917 ( .A(n13667), .B(n13668), .Z(n13663) );
  XNOR U13918 ( .A(n13669), .B(n13670), .Z(n13668) );
  ANDN U13919 ( .B(n13671), .A(n13672), .Z(n13670) );
  XOR U13920 ( .A(n13625), .B(n13673), .Z(n13639) );
  XNOR U13921 ( .A(n13674), .B(n13631), .Z(n13673) );
  OR U13922 ( .A(n11709), .B(n13576), .Z(n13631) );
  XNOR U13923 ( .A(n13651), .B(n12639), .Z(n13576) );
  IV U13924 ( .A(n13641), .Z(n12639) );
  XNOR U13925 ( .A(n13632), .B(n11606), .Z(n11709) );
  IV U13926 ( .A(n11711), .Z(n13632) );
  ANDN U13927 ( .B(n11606), .A(n13641), .Z(n13674) );
  XNOR U13928 ( .A(n13675), .B(n13676), .Z(n13641) );
  XNOR U13929 ( .A(n13652), .B(n13677), .Z(n11606) );
  XNOR U13930 ( .A(n13645), .B(n13675), .Z(n13677) );
  XNOR U13931 ( .A(n13575), .B(n11711), .Z(n13625) );
  XOR U13932 ( .A(n13652), .B(n13678), .Z(n11711) );
  XNOR U13933 ( .A(n13654), .B(n13648), .Z(n13678) );
  XOR U13934 ( .A(n13679), .B(n13680), .Z(n13648) );
  XNOR U13935 ( .A(n9171), .B(n9141), .Z(n13680) );
  XNOR U13936 ( .A(n11271), .B(n11257), .Z(n9141) );
  XNOR U13937 ( .A(n13681), .B(n13682), .Z(n11271) );
  XNOR U13938 ( .A(n13683), .B(n13684), .Z(n13681) );
  XOR U13939 ( .A(n10076), .B(n13657), .Z(n9171) );
  IV U13940 ( .A(n13662), .Z(n10076) );
  XNOR U13941 ( .A(key[783]), .B(n11255), .Z(n13679) );
  XOR U13942 ( .A(n13685), .B(n13686), .Z(n11255) );
  XOR U13943 ( .A(n13687), .B(n13688), .Z(n13686) );
  XOR U13944 ( .A(n13689), .B(n13690), .Z(n13685) );
  IV U13945 ( .A(n13676), .Z(n13652) );
  XOR U13946 ( .A(n13691), .B(n13692), .Z(n13676) );
  XNOR U13947 ( .A(n13693), .B(n11247), .Z(n13692) );
  XNOR U13948 ( .A(n13694), .B(n13695), .Z(n11247) );
  XOR U13949 ( .A(n13658), .B(n13688), .Z(n13695) );
  XNOR U13950 ( .A(n13696), .B(n13697), .Z(n13688) );
  XNOR U13951 ( .A(n13698), .B(n13699), .Z(n13697) );
  NANDN U13952 ( .A(n13700), .B(n13701), .Z(n13699) );
  XOR U13953 ( .A(n13702), .B(n13703), .Z(n13694) );
  XNOR U13954 ( .A(n13704), .B(n13705), .Z(n13703) );
  ANDN U13955 ( .B(n13706), .A(n13707), .Z(n13705) );
  XNOR U13956 ( .A(n9136), .B(n13708), .Z(n13691) );
  XNOR U13957 ( .A(key[781]), .B(n9154), .Z(n13708) );
  XOR U13958 ( .A(n13709), .B(n13710), .Z(n9154) );
  XOR U13959 ( .A(n11260), .B(n11244), .Z(n9136) );
  IV U13960 ( .A(n10046), .Z(n11244) );
  XNOR U13961 ( .A(n13711), .B(n13712), .Z(n10046) );
  XNOR U13962 ( .A(n13661), .B(n13683), .Z(n13712) );
  XNOR U13963 ( .A(n13713), .B(n13714), .Z(n13683) );
  XNOR U13964 ( .A(n13715), .B(n13716), .Z(n13714) );
  OR U13965 ( .A(n13717), .B(n13718), .Z(n13716) );
  XNOR U13966 ( .A(n13719), .B(n13720), .Z(n13711) );
  XOR U13967 ( .A(n13721), .B(n13722), .Z(n13720) );
  ANDN U13968 ( .B(n13723), .A(n13724), .Z(n13722) );
  XNOR U13969 ( .A(n13725), .B(n13726), .Z(n11260) );
  XNOR U13970 ( .A(n13727), .B(n13728), .Z(n13726) );
  XNOR U13971 ( .A(n13729), .B(n13730), .Z(n13725) );
  XOR U13972 ( .A(n13731), .B(n13732), .Z(n13730) );
  ANDN U13973 ( .B(n13733), .A(n13734), .Z(n13732) );
  IV U13974 ( .A(n13651), .Z(n13575) );
  XOR U13975 ( .A(n13675), .B(n13735), .Z(n13651) );
  XNOR U13976 ( .A(n13644), .B(n13650), .Z(n13735) );
  XOR U13977 ( .A(n13736), .B(n13737), .Z(n13650) );
  XOR U13978 ( .A(n13645), .B(n13738), .Z(n13737) );
  XOR U13979 ( .A(n9157), .B(n10066), .Z(n13738) );
  XOR U13980 ( .A(n13657), .B(n11245), .Z(n10066) );
  XOR U13981 ( .A(n13727), .B(n11292), .Z(n11245) );
  IV U13982 ( .A(n10051), .Z(n13657) );
  XNOR U13983 ( .A(n13662), .B(n9130), .Z(n9157) );
  XNOR U13984 ( .A(n13665), .B(n9148), .Z(n9130) );
  XNOR U13985 ( .A(n13739), .B(n13740), .Z(n13645) );
  XOR U13986 ( .A(n11292), .B(n10075), .Z(n13740) );
  XNOR U13987 ( .A(n10069), .B(n11280), .Z(n10075) );
  XOR U13988 ( .A(n13741), .B(n13742), .Z(n10069) );
  XNOR U13989 ( .A(n13684), .B(n13743), .Z(n13742) );
  XNOR U13990 ( .A(n9148), .B(n13744), .Z(n13739) );
  XNOR U13991 ( .A(key[777]), .B(n11268), .Z(n13744) );
  XOR U13992 ( .A(n13687), .B(n13745), .Z(n11268) );
  XOR U13993 ( .A(n13746), .B(n13690), .Z(n13745) );
  XOR U13994 ( .A(n13747), .B(n13748), .Z(n9148) );
  XNOR U13995 ( .A(n9159), .B(n13749), .Z(n13736) );
  XOR U13996 ( .A(key[779]), .B(n11290), .Z(n13749) );
  XNOR U13997 ( .A(n13750), .B(n13751), .Z(n11290) );
  XNOR U13998 ( .A(n13690), .B(n13687), .Z(n13751) );
  XNOR U13999 ( .A(n13752), .B(n13753), .Z(n13687) );
  XNOR U14000 ( .A(n13754), .B(n13755), .Z(n13753) );
  NANDN U14001 ( .A(n13756), .B(n13701), .Z(n13755) );
  XOR U14002 ( .A(n13757), .B(n13758), .Z(n13750) );
  XOR U14003 ( .A(n11284), .B(n10070), .Z(n9159) );
  XNOR U14004 ( .A(n13759), .B(n13682), .Z(n10070) );
  XOR U14005 ( .A(n13743), .B(n13741), .Z(n13682) );
  XOR U14006 ( .A(n13760), .B(n13761), .Z(n13743) );
  XNOR U14007 ( .A(n13762), .B(n13763), .Z(n13761) );
  NANDN U14008 ( .A(n13717), .B(n13764), .Z(n13763) );
  XNOR U14009 ( .A(n13765), .B(n13766), .Z(n13759) );
  XOR U14010 ( .A(n13767), .B(n13768), .Z(n13644) );
  XNOR U14011 ( .A(n9147), .B(n11284), .Z(n13768) );
  XOR U14012 ( .A(n13769), .B(n13770), .Z(n11284) );
  XNOR U14013 ( .A(n13771), .B(n13772), .Z(n13769) );
  XNOR U14014 ( .A(n11292), .B(n10055), .Z(n9147) );
  XNOR U14015 ( .A(n13773), .B(n13741), .Z(n10055) );
  XNOR U14016 ( .A(n13774), .B(n13775), .Z(n13741) );
  XNOR U14017 ( .A(n13776), .B(n13777), .Z(n13775) );
  NANDN U14018 ( .A(n13778), .B(n13723), .Z(n13777) );
  XNOR U14019 ( .A(n13779), .B(n13780), .Z(n11292) );
  XOR U14020 ( .A(n11287), .B(n13781), .Z(n13767) );
  XOR U14021 ( .A(key[778]), .B(n11281), .Z(n13781) );
  XOR U14022 ( .A(n13782), .B(n13690), .Z(n11281) );
  XOR U14023 ( .A(n13783), .B(n13784), .Z(n13690) );
  XNOR U14024 ( .A(n13785), .B(n13786), .Z(n13784) );
  NANDN U14025 ( .A(n13787), .B(n13706), .Z(n13786) );
  XNOR U14026 ( .A(n13788), .B(n13789), .Z(n11287) );
  XNOR U14027 ( .A(n13790), .B(n13710), .Z(n13788) );
  XNOR U14028 ( .A(n13791), .B(n13792), .Z(n13710) );
  XOR U14029 ( .A(n13793), .B(n13669), .Z(n13792) );
  NANDN U14030 ( .A(n13794), .B(n13795), .Z(n13669) );
  NOR U14031 ( .A(n13796), .B(n13797), .Z(n13793) );
  IV U14032 ( .A(n13654), .Z(n13675) );
  XOR U14033 ( .A(n13798), .B(n13799), .Z(n13654) );
  XOR U14034 ( .A(n10058), .B(n11601), .Z(n13799) );
  IV U14035 ( .A(n13636), .Z(n11601) );
  XOR U14036 ( .A(n13800), .B(n13801), .Z(n13636) );
  XNOR U14037 ( .A(n11280), .B(n10074), .Z(n13801) );
  XOR U14038 ( .A(n9142), .B(n9172), .Z(n10074) );
  XOR U14039 ( .A(n13661), .B(n13802), .Z(n9172) );
  XNOR U14040 ( .A(n13713), .B(n13803), .Z(n13661) );
  XOR U14041 ( .A(n13804), .B(n13776), .Z(n13803) );
  OR U14042 ( .A(n13805), .B(n13806), .Z(n13776) );
  ANDN U14043 ( .B(n13807), .A(n13808), .Z(n13804) );
  XNOR U14044 ( .A(n13774), .B(n13809), .Z(n13713) );
  XNOR U14045 ( .A(n13810), .B(n13811), .Z(n13809) );
  NAND U14046 ( .A(n13812), .B(n13813), .Z(n13811) );
  XOR U14047 ( .A(n13782), .B(n13658), .Z(n9142) );
  XOR U14048 ( .A(n13696), .B(n13814), .Z(n13658) );
  XOR U14049 ( .A(n13815), .B(n13785), .Z(n13814) );
  NANDN U14050 ( .A(n13816), .B(n13817), .Z(n13785) );
  ANDN U14051 ( .B(n13818), .A(n13819), .Z(n13815) );
  XNOR U14052 ( .A(n13783), .B(n13820), .Z(n13696) );
  XNOR U14053 ( .A(n13821), .B(n13822), .Z(n13820) );
  NAND U14054 ( .A(n13823), .B(n13824), .Z(n13822) );
  XNOR U14055 ( .A(n13780), .B(n13825), .Z(n11280) );
  XNOR U14056 ( .A(n13826), .B(n13827), .Z(n13825) );
  XNOR U14057 ( .A(n10051), .B(n13828), .Z(n13800) );
  XOR U14058 ( .A(key[776]), .B(n11283), .Z(n13828) );
  IV U14059 ( .A(n9167), .Z(n11283) );
  XNOR U14060 ( .A(n13748), .B(n13829), .Z(n9167) );
  XNOR U14061 ( .A(n13709), .B(n13830), .Z(n13829) );
  XNOR U14062 ( .A(n10051), .B(n11257), .Z(n10058) );
  XOR U14063 ( .A(n13831), .B(n13770), .Z(n11257) );
  XOR U14064 ( .A(n13827), .B(n13780), .Z(n13770) );
  XNOR U14065 ( .A(n13832), .B(n13833), .Z(n13780) );
  XOR U14066 ( .A(n13834), .B(n13835), .Z(n13833) );
  NANDN U14067 ( .A(n13836), .B(n13733), .Z(n13835) );
  XOR U14068 ( .A(n13837), .B(n13838), .Z(n13827) );
  XNOR U14069 ( .A(n13839), .B(n13840), .Z(n13838) );
  NANDN U14070 ( .A(n13841), .B(n13842), .Z(n13840) );
  XNOR U14071 ( .A(n13728), .B(n13826), .Z(n13831) );
  XNOR U14072 ( .A(n13843), .B(n13844), .Z(n13728) );
  XNOR U14073 ( .A(n13845), .B(n13846), .Z(n13844) );
  OR U14074 ( .A(n13841), .B(n13847), .Z(n13846) );
  XOR U14075 ( .A(n13727), .B(n13848), .Z(n10051) );
  XNOR U14076 ( .A(n13843), .B(n13849), .Z(n13727) );
  XNOR U14077 ( .A(n13850), .B(n13834), .Z(n13849) );
  ANDN U14078 ( .B(n13853), .A(n13854), .Z(n13850) );
  XNOR U14079 ( .A(n13832), .B(n13855), .Z(n13843) );
  XNOR U14080 ( .A(n13856), .B(n13857), .Z(n13855) );
  NAND U14081 ( .A(n13858), .B(n13859), .Z(n13857) );
  XOR U14082 ( .A(n9151), .B(n13860), .Z(n13798) );
  XNOR U14083 ( .A(key[782]), .B(n11262), .Z(n13860) );
  XNOR U14084 ( .A(n13746), .B(n13758), .Z(n11262) );
  XOR U14085 ( .A(n13752), .B(n13861), .Z(n13758) );
  XOR U14086 ( .A(n13862), .B(n13704), .Z(n13861) );
  NANDN U14087 ( .A(n13863), .B(n13817), .Z(n13704) );
  XNOR U14088 ( .A(n13819), .B(n13706), .Z(n13817) );
  NOR U14089 ( .A(n13864), .B(n13819), .Z(n13862) );
  XNOR U14090 ( .A(n13702), .B(n13865), .Z(n13752) );
  XNOR U14091 ( .A(n13866), .B(n13867), .Z(n13865) );
  NAND U14092 ( .A(n13868), .B(n13823), .Z(n13867) );
  IV U14093 ( .A(n13689), .Z(n13746) );
  XNOR U14094 ( .A(n13782), .B(n13757), .Z(n13689) );
  XNOR U14095 ( .A(n13754), .B(n13870), .Z(n13869) );
  NANDN U14096 ( .A(n13871), .B(n13872), .Z(n13870) );
  OR U14097 ( .A(n13873), .B(n13874), .Z(n13754) );
  XNOR U14098 ( .A(n13875), .B(n13866), .Z(n13702) );
  NANDN U14099 ( .A(n13876), .B(n13877), .Z(n13866) );
  ANDN U14100 ( .B(n13878), .A(n13879), .Z(n13875) );
  XOR U14101 ( .A(n13783), .B(n13880), .Z(n13782) );
  XOR U14102 ( .A(n13881), .B(n13698), .Z(n13880) );
  OR U14103 ( .A(n13873), .B(n13882), .Z(n13698) );
  XNOR U14104 ( .A(n13701), .B(n13872), .Z(n13873) );
  ANDN U14105 ( .B(n13883), .A(n13884), .Z(n13881) );
  XOR U14106 ( .A(n13885), .B(n13821), .Z(n13783) );
  OR U14107 ( .A(n13876), .B(n13886), .Z(n13821) );
  XNOR U14108 ( .A(n13887), .B(n13823), .Z(n13876) );
  XOR U14109 ( .A(n13872), .B(n13706), .Z(n13823) );
  XOR U14110 ( .A(n13888), .B(n13889), .Z(n13706) );
  NANDN U14111 ( .A(n13890), .B(n13891), .Z(n13889) );
  IV U14112 ( .A(n13884), .Z(n13872) );
  XNOR U14113 ( .A(n13892), .B(n13893), .Z(n13884) );
  NANDN U14114 ( .A(n13890), .B(n13894), .Z(n13893) );
  ANDN U14115 ( .B(n13887), .A(n13895), .Z(n13885) );
  IV U14116 ( .A(n13879), .Z(n13887) );
  XOR U14117 ( .A(n13819), .B(n13701), .Z(n13879) );
  XNOR U14118 ( .A(n13896), .B(n13892), .Z(n13701) );
  NANDN U14119 ( .A(n13897), .B(n13898), .Z(n13892) );
  XOR U14120 ( .A(n13894), .B(n13899), .Z(n13898) );
  ANDN U14121 ( .B(n13899), .A(n13900), .Z(n13896) );
  XOR U14122 ( .A(n13901), .B(n13888), .Z(n13819) );
  NANDN U14123 ( .A(n13897), .B(n13902), .Z(n13888) );
  XOR U14124 ( .A(n13903), .B(n13891), .Z(n13902) );
  XNOR U14125 ( .A(n13904), .B(n13905), .Z(n13890) );
  XOR U14126 ( .A(n13906), .B(n13907), .Z(n13905) );
  XNOR U14127 ( .A(n13908), .B(n13909), .Z(n13904) );
  XNOR U14128 ( .A(n13910), .B(n13911), .Z(n13909) );
  ANDN U14129 ( .B(n13903), .A(n13907), .Z(n13910) );
  ANDN U14130 ( .B(n13903), .A(n13900), .Z(n13901) );
  XNOR U14131 ( .A(n13906), .B(n13912), .Z(n13900) );
  XOR U14132 ( .A(n13913), .B(n13911), .Z(n13912) );
  NAND U14133 ( .A(n13914), .B(n13915), .Z(n13911) );
  XNOR U14134 ( .A(n13908), .B(n13891), .Z(n13915) );
  IV U14135 ( .A(n13903), .Z(n13908) );
  XNOR U14136 ( .A(n13894), .B(n13907), .Z(n13914) );
  IV U14137 ( .A(n13899), .Z(n13907) );
  XOR U14138 ( .A(n13916), .B(n13917), .Z(n13899) );
  XNOR U14139 ( .A(n13918), .B(n13919), .Z(n13917) );
  XNOR U14140 ( .A(n13920), .B(n13921), .Z(n13916) );
  ANDN U14141 ( .B(n13818), .A(n13864), .Z(n13920) );
  AND U14142 ( .A(n13891), .B(n13894), .Z(n13913) );
  XNOR U14143 ( .A(n13891), .B(n13894), .Z(n13906) );
  XNOR U14144 ( .A(n13922), .B(n13923), .Z(n13894) );
  XNOR U14145 ( .A(n13924), .B(n13919), .Z(n13923) );
  XOR U14146 ( .A(n13925), .B(n13926), .Z(n13922) );
  XNOR U14147 ( .A(n13927), .B(n13921), .Z(n13926) );
  OR U14148 ( .A(n13863), .B(n13816), .Z(n13921) );
  XNOR U14149 ( .A(n13818), .B(n13928), .Z(n13816) );
  XNOR U14150 ( .A(n13864), .B(n13707), .Z(n13863) );
  ANDN U14151 ( .B(n13929), .A(n13787), .Z(n13927) );
  XNOR U14152 ( .A(n13930), .B(n13931), .Z(n13891) );
  XNOR U14153 ( .A(n13919), .B(n13932), .Z(n13931) );
  XOR U14154 ( .A(n13756), .B(n13925), .Z(n13932) );
  XNOR U14155 ( .A(n13818), .B(n13864), .Z(n13919) );
  XNOR U14156 ( .A(n13933), .B(n13934), .Z(n13930) );
  XNOR U14157 ( .A(n13935), .B(n13936), .Z(n13934) );
  ANDN U14158 ( .B(n13883), .A(n13871), .Z(n13935) );
  XNOR U14159 ( .A(n13937), .B(n13938), .Z(n13903) );
  XNOR U14160 ( .A(n13924), .B(n13939), .Z(n13938) );
  XNOR U14161 ( .A(n13871), .B(n13918), .Z(n13939) );
  XOR U14162 ( .A(n13925), .B(n13940), .Z(n13918) );
  XNOR U14163 ( .A(n13941), .B(n13942), .Z(n13940) );
  NAND U14164 ( .A(n13824), .B(n13868), .Z(n13942) );
  XNOR U14165 ( .A(n13943), .B(n13941), .Z(n13925) );
  NANDN U14166 ( .A(n13886), .B(n13877), .Z(n13941) );
  XOR U14167 ( .A(n13878), .B(n13868), .Z(n13877) );
  XNOR U14168 ( .A(n13944), .B(n13707), .Z(n13868) );
  XOR U14169 ( .A(n13895), .B(n13824), .Z(n13886) );
  XOR U14170 ( .A(n13883), .B(n13928), .Z(n13824) );
  ANDN U14171 ( .B(n13878), .A(n13895), .Z(n13943) );
  XNOR U14172 ( .A(n13933), .B(n13818), .Z(n13895) );
  XNOR U14173 ( .A(n13945), .B(n13946), .Z(n13818) );
  XNOR U14174 ( .A(n13947), .B(n13948), .Z(n13946) );
  XOR U14175 ( .A(n13949), .B(n13950), .Z(n13878) );
  XOR U14176 ( .A(n13928), .B(n13929), .Z(n13924) );
  IV U14177 ( .A(n13707), .Z(n13929) );
  XOR U14178 ( .A(n13951), .B(n13952), .Z(n13707) );
  XNOR U14179 ( .A(n13953), .B(n13948), .Z(n13952) );
  IV U14180 ( .A(n13787), .Z(n13928) );
  XOR U14181 ( .A(n13948), .B(n13954), .Z(n13787) );
  XNOR U14182 ( .A(n13883), .B(n13955), .Z(n13937) );
  XNOR U14183 ( .A(n13956), .B(n13936), .Z(n13955) );
  OR U14184 ( .A(n13874), .B(n13882), .Z(n13936) );
  XNOR U14185 ( .A(n13933), .B(n13883), .Z(n13882) );
  XOR U14186 ( .A(n13756), .B(n13944), .Z(n13874) );
  IV U14187 ( .A(n13871), .Z(n13944) );
  XOR U14188 ( .A(n13950), .B(n13957), .Z(n13871) );
  XNOR U14189 ( .A(n13953), .B(n13945), .Z(n13957) );
  XOR U14190 ( .A(n13958), .B(n13959), .Z(n13945) );
  XOR U14191 ( .A(n12152), .B(n12149), .Z(n13959) );
  XOR U14192 ( .A(n13960), .B(n12160), .Z(n12152) );
  XOR U14193 ( .A(key[754]), .B(n13563), .Z(n13958) );
  IV U14194 ( .A(n13864), .Z(n13950) );
  XOR U14195 ( .A(n13951), .B(n13961), .Z(n13864) );
  XOR U14196 ( .A(n13948), .B(n13962), .Z(n13961) );
  ANDN U14197 ( .B(n13949), .A(n13700), .Z(n13956) );
  IV U14198 ( .A(n13756), .Z(n13949) );
  XOR U14199 ( .A(n13951), .B(n13963), .Z(n13756) );
  XOR U14200 ( .A(n13948), .B(n13964), .Z(n13963) );
  XOR U14201 ( .A(n13965), .B(n13966), .Z(n13948) );
  XNOR U14202 ( .A(n13967), .B(n13700), .Z(n13966) );
  IV U14203 ( .A(n13933), .Z(n13700) );
  XOR U14204 ( .A(n13968), .B(n13969), .Z(n13965) );
  XNOR U14205 ( .A(key[758]), .B(n13545), .Z(n13969) );
  XOR U14206 ( .A(n12143), .B(n13970), .Z(n13545) );
  XNOR U14207 ( .A(n13540), .B(n13971), .Z(n12143) );
  IV U14208 ( .A(n13954), .Z(n13951) );
  XOR U14209 ( .A(n13972), .B(n13973), .Z(n13954) );
  XNOR U14210 ( .A(n13538), .B(n13974), .Z(n13973) );
  XNOR U14211 ( .A(n13522), .B(n13975), .Z(n13538) );
  XNOR U14212 ( .A(key[757]), .B(n13976), .Z(n13972) );
  XOR U14213 ( .A(n13977), .B(n13978), .Z(n13883) );
  XNOR U14214 ( .A(n13964), .B(n13962), .Z(n13978) );
  XNOR U14215 ( .A(n13979), .B(n13980), .Z(n13962) );
  XOR U14216 ( .A(n13970), .B(n13533), .Z(n13980) );
  XOR U14217 ( .A(n13553), .B(n13981), .Z(n13533) );
  XOR U14218 ( .A(n13982), .B(n13983), .Z(n13970) );
  XOR U14219 ( .A(key[759]), .B(n13984), .Z(n13979) );
  XNOR U14220 ( .A(n13985), .B(n13986), .Z(n13964) );
  XNOR U14221 ( .A(n13519), .B(n13987), .Z(n13986) );
  XOR U14222 ( .A(n13988), .B(n12125), .Z(n13519) );
  XNOR U14223 ( .A(n13521), .B(n13989), .Z(n13985) );
  XNOR U14224 ( .A(key[756]), .B(n13990), .Z(n13989) );
  XOR U14225 ( .A(n13982), .B(n13976), .Z(n13521) );
  XOR U14226 ( .A(n13933), .B(n13947), .Z(n13977) );
  XOR U14227 ( .A(n13991), .B(n13992), .Z(n13947) );
  XNOR U14228 ( .A(n13953), .B(n13993), .Z(n13992) );
  XNOR U14229 ( .A(n13569), .B(n13994), .Z(n13993) );
  XOR U14230 ( .A(n13995), .B(n13996), .Z(n13953) );
  XOR U14231 ( .A(n12169), .B(n13997), .Z(n13996) );
  XNOR U14232 ( .A(n13549), .B(n12154), .Z(n12169) );
  XOR U14233 ( .A(key[753]), .B(n13998), .Z(n13995) );
  XNOR U14234 ( .A(n13565), .B(n13999), .Z(n13991) );
  XNOR U14235 ( .A(key[755]), .B(n12162), .Z(n13999) );
  XOR U14236 ( .A(n13572), .B(n12157), .Z(n12162) );
  XNOR U14237 ( .A(n12168), .B(n13990), .Z(n13565) );
  IV U14238 ( .A(n13982), .Z(n12168) );
  XOR U14239 ( .A(n14000), .B(n14001), .Z(n13933) );
  XOR U14240 ( .A(key[752]), .B(n14002), .Z(n14000) );
  XOR U14241 ( .A(n10044), .B(n9140), .Z(n9151) );
  XOR U14242 ( .A(n13662), .B(n11256), .Z(n9140) );
  XNOR U14243 ( .A(n14003), .B(n13789), .Z(n11256) );
  XOR U14244 ( .A(n13830), .B(n13748), .Z(n13789) );
  XOR U14245 ( .A(n14004), .B(n14005), .Z(n13748) );
  XNOR U14246 ( .A(n14006), .B(n14007), .Z(n14005) );
  NANDN U14247 ( .A(n14008), .B(n13671), .Z(n14007) );
  XOR U14248 ( .A(n13791), .B(n14009), .Z(n13830) );
  XNOR U14249 ( .A(n14010), .B(n14011), .Z(n14009) );
  NANDN U14250 ( .A(n14012), .B(n14013), .Z(n14011) );
  XNOR U14251 ( .A(n13667), .B(n14014), .Z(n13791) );
  XNOR U14252 ( .A(n14015), .B(n14016), .Z(n14014) );
  NAND U14253 ( .A(n14017), .B(n14018), .Z(n14016) );
  XNOR U14254 ( .A(n13709), .B(n13666), .Z(n14003) );
  XNOR U14255 ( .A(n14019), .B(n14020), .Z(n13666) );
  XNOR U14256 ( .A(n14021), .B(n14022), .Z(n14020) );
  NANDN U14257 ( .A(n14023), .B(n14013), .Z(n14022) );
  XOR U14258 ( .A(n13747), .B(n13790), .Z(n13709) );
  XOR U14259 ( .A(n13667), .B(n14024), .Z(n13790) );
  XNOR U14260 ( .A(n14010), .B(n14025), .Z(n14024) );
  NANDN U14261 ( .A(n14026), .B(n14027), .Z(n14025) );
  OR U14262 ( .A(n14028), .B(n14029), .Z(n14010) );
  XOR U14263 ( .A(n14030), .B(n14015), .Z(n13667) );
  NANDN U14264 ( .A(n14031), .B(n14032), .Z(n14015) );
  ANDN U14265 ( .B(n14033), .A(n14034), .Z(n14030) );
  XOR U14266 ( .A(n13747), .B(n13665), .Z(n13662) );
  XNOR U14267 ( .A(n14019), .B(n14035), .Z(n13665) );
  XOR U14268 ( .A(n14036), .B(n14006), .Z(n14035) );
  NANDN U14269 ( .A(n14037), .B(n13795), .Z(n14006) );
  XNOR U14270 ( .A(n13797), .B(n13671), .Z(n13795) );
  ANDN U14271 ( .B(n14038), .A(n13797), .Z(n14036) );
  XOR U14272 ( .A(n14004), .B(n14039), .Z(n14019) );
  XNOR U14273 ( .A(n14040), .B(n14041), .Z(n14039) );
  NAND U14274 ( .A(n14018), .B(n14042), .Z(n14041) );
  XOR U14275 ( .A(n14044), .B(n14021), .Z(n14043) );
  OR U14276 ( .A(n14045), .B(n14028), .Z(n14021) );
  XNOR U14277 ( .A(n14013), .B(n14027), .Z(n14028) );
  ANDN U14278 ( .B(n14046), .A(n14047), .Z(n14044) );
  XNOR U14279 ( .A(n14048), .B(n14040), .Z(n14004) );
  OR U14280 ( .A(n14031), .B(n14049), .Z(n14040) );
  XNOR U14281 ( .A(n14050), .B(n14018), .Z(n14031) );
  XOR U14282 ( .A(n14027), .B(n13671), .Z(n14018) );
  XOR U14283 ( .A(n14051), .B(n14052), .Z(n13671) );
  NANDN U14284 ( .A(n14053), .B(n14054), .Z(n14052) );
  IV U14285 ( .A(n14047), .Z(n14027) );
  XNOR U14286 ( .A(n14055), .B(n14056), .Z(n14047) );
  NANDN U14287 ( .A(n14053), .B(n14057), .Z(n14056) );
  ANDN U14288 ( .B(n14050), .A(n14058), .Z(n14048) );
  IV U14289 ( .A(n14034), .Z(n14050) );
  XOR U14290 ( .A(n13797), .B(n14013), .Z(n14034) );
  XNOR U14291 ( .A(n14059), .B(n14055), .Z(n14013) );
  NANDN U14292 ( .A(n14060), .B(n14061), .Z(n14055) );
  XOR U14293 ( .A(n14057), .B(n14062), .Z(n14061) );
  ANDN U14294 ( .B(n14062), .A(n14063), .Z(n14059) );
  XOR U14295 ( .A(n14064), .B(n14051), .Z(n13797) );
  NANDN U14296 ( .A(n14060), .B(n14065), .Z(n14051) );
  XOR U14297 ( .A(n14066), .B(n14054), .Z(n14065) );
  XNOR U14298 ( .A(n14067), .B(n14068), .Z(n14053) );
  XOR U14299 ( .A(n14069), .B(n14070), .Z(n14068) );
  XNOR U14300 ( .A(n14071), .B(n14072), .Z(n14067) );
  XNOR U14301 ( .A(n14073), .B(n14074), .Z(n14072) );
  ANDN U14302 ( .B(n14066), .A(n14070), .Z(n14073) );
  ANDN U14303 ( .B(n14066), .A(n14063), .Z(n14064) );
  XNOR U14304 ( .A(n14069), .B(n14075), .Z(n14063) );
  XOR U14305 ( .A(n14076), .B(n14074), .Z(n14075) );
  NAND U14306 ( .A(n14077), .B(n14078), .Z(n14074) );
  XNOR U14307 ( .A(n14071), .B(n14054), .Z(n14078) );
  IV U14308 ( .A(n14066), .Z(n14071) );
  XNOR U14309 ( .A(n14057), .B(n14070), .Z(n14077) );
  IV U14310 ( .A(n14062), .Z(n14070) );
  XOR U14311 ( .A(n14079), .B(n14080), .Z(n14062) );
  XNOR U14312 ( .A(n14081), .B(n14082), .Z(n14080) );
  XNOR U14313 ( .A(n14083), .B(n14084), .Z(n14079) );
  ANDN U14314 ( .B(n14038), .A(n13796), .Z(n14083) );
  AND U14315 ( .A(n14054), .B(n14057), .Z(n14076) );
  XNOR U14316 ( .A(n14054), .B(n14057), .Z(n14069) );
  XNOR U14317 ( .A(n14085), .B(n14086), .Z(n14057) );
  XNOR U14318 ( .A(n14087), .B(n14082), .Z(n14086) );
  XOR U14319 ( .A(n14088), .B(n14089), .Z(n14085) );
  XNOR U14320 ( .A(n14090), .B(n14084), .Z(n14089) );
  OR U14321 ( .A(n13794), .B(n14037), .Z(n14084) );
  XNOR U14322 ( .A(n14038), .B(n14091), .Z(n14037) );
  XNOR U14323 ( .A(n13796), .B(n13672), .Z(n13794) );
  ANDN U14324 ( .B(n14092), .A(n14008), .Z(n14090) );
  XNOR U14325 ( .A(n14093), .B(n14094), .Z(n14054) );
  XNOR U14326 ( .A(n14082), .B(n14095), .Z(n14094) );
  XOR U14327 ( .A(n14012), .B(n14088), .Z(n14095) );
  XNOR U14328 ( .A(n14038), .B(n13796), .Z(n14082) );
  XNOR U14329 ( .A(n14096), .B(n14097), .Z(n14093) );
  XNOR U14330 ( .A(n14098), .B(n14099), .Z(n14097) );
  ANDN U14331 ( .B(n14046), .A(n14026), .Z(n14098) );
  XNOR U14332 ( .A(n14100), .B(n14101), .Z(n14066) );
  XNOR U14333 ( .A(n14087), .B(n14102), .Z(n14101) );
  XNOR U14334 ( .A(n14026), .B(n14081), .Z(n14102) );
  XOR U14335 ( .A(n14088), .B(n14103), .Z(n14081) );
  XNOR U14336 ( .A(n14104), .B(n14105), .Z(n14103) );
  NAND U14337 ( .A(n14042), .B(n14017), .Z(n14105) );
  XNOR U14338 ( .A(n14106), .B(n14104), .Z(n14088) );
  NANDN U14339 ( .A(n14049), .B(n14032), .Z(n14104) );
  XOR U14340 ( .A(n14033), .B(n14017), .Z(n14032) );
  XNOR U14341 ( .A(n14107), .B(n13672), .Z(n14017) );
  XOR U14342 ( .A(n14058), .B(n14042), .Z(n14049) );
  XOR U14343 ( .A(n14046), .B(n14091), .Z(n14042) );
  ANDN U14344 ( .B(n14033), .A(n14058), .Z(n14106) );
  XNOR U14345 ( .A(n14096), .B(n14038), .Z(n14058) );
  XNOR U14346 ( .A(n14108), .B(n14109), .Z(n14038) );
  XNOR U14347 ( .A(n14110), .B(n14111), .Z(n14109) );
  XOR U14348 ( .A(n14112), .B(n14113), .Z(n14033) );
  XOR U14349 ( .A(n14091), .B(n14092), .Z(n14087) );
  IV U14350 ( .A(n13672), .Z(n14092) );
  XOR U14351 ( .A(n14114), .B(n14115), .Z(n13672) );
  XNOR U14352 ( .A(n14116), .B(n14111), .Z(n14115) );
  IV U14353 ( .A(n14008), .Z(n14091) );
  XOR U14354 ( .A(n14111), .B(n14117), .Z(n14008) );
  XNOR U14355 ( .A(n14046), .B(n14118), .Z(n14100) );
  XNOR U14356 ( .A(n14119), .B(n14099), .Z(n14118) );
  OR U14357 ( .A(n14029), .B(n14045), .Z(n14099) );
  XNOR U14358 ( .A(n14096), .B(n14046), .Z(n14045) );
  XOR U14359 ( .A(n14012), .B(n14107), .Z(n14029) );
  IV U14360 ( .A(n14026), .Z(n14107) );
  XOR U14361 ( .A(n14113), .B(n14120), .Z(n14026) );
  XNOR U14362 ( .A(n14116), .B(n14108), .Z(n14120) );
  XOR U14363 ( .A(n14121), .B(n14122), .Z(n14108) );
  XOR U14364 ( .A(n12482), .B(n14123), .Z(n14122) );
  XOR U14365 ( .A(n14124), .B(n14125), .Z(n14121) );
  XOR U14366 ( .A(key[714]), .B(n14126), .Z(n14125) );
  IV U14367 ( .A(n13796), .Z(n14113) );
  XOR U14368 ( .A(n14114), .B(n14127), .Z(n13796) );
  XOR U14369 ( .A(n14111), .B(n14128), .Z(n14127) );
  ANDN U14370 ( .B(n14112), .A(n14023), .Z(n14119) );
  IV U14371 ( .A(n14012), .Z(n14112) );
  XOR U14372 ( .A(n14114), .B(n14129), .Z(n14012) );
  XOR U14373 ( .A(n14111), .B(n14130), .Z(n14129) );
  XOR U14374 ( .A(n14131), .B(n14132), .Z(n14111) );
  XNOR U14375 ( .A(n14133), .B(n14023), .Z(n14132) );
  IV U14376 ( .A(n14096), .Z(n14023) );
  XNOR U14377 ( .A(n12458), .B(n14134), .Z(n14131) );
  XNOR U14378 ( .A(key[718]), .B(n13089), .Z(n14134) );
  XNOR U14379 ( .A(n13105), .B(n14135), .Z(n13089) );
  IV U14380 ( .A(n14117), .Z(n14114) );
  XOR U14381 ( .A(n14136), .B(n14137), .Z(n14117) );
  XNOR U14382 ( .A(n12475), .B(n14138), .Z(n14137) );
  XNOR U14383 ( .A(n13094), .B(n14139), .Z(n14136) );
  XNOR U14384 ( .A(key[717]), .B(n14140), .Z(n14139) );
  XOR U14385 ( .A(n14141), .B(n14142), .Z(n14046) );
  XNOR U14386 ( .A(n14130), .B(n14128), .Z(n14142) );
  XNOR U14387 ( .A(n14143), .B(n14144), .Z(n14128) );
  XOR U14388 ( .A(n12496), .B(n14145), .Z(n14144) );
  XNOR U14389 ( .A(key[719]), .B(n13101), .Z(n14143) );
  XNOR U14390 ( .A(n14146), .B(n14147), .Z(n14130) );
  XNOR U14391 ( .A(n13108), .B(n14148), .Z(n14146) );
  XNOR U14392 ( .A(key[716]), .B(n13111), .Z(n14148) );
  XNOR U14393 ( .A(n13105), .B(n14149), .Z(n13111) );
  XOR U14394 ( .A(n14096), .B(n14110), .Z(n14141) );
  XOR U14395 ( .A(n14150), .B(n14151), .Z(n14110) );
  XNOR U14396 ( .A(n14116), .B(n14152), .Z(n14151) );
  XOR U14397 ( .A(n14153), .B(n14154), .Z(n14152) );
  XOR U14398 ( .A(n14155), .B(n14156), .Z(n14116) );
  XNOR U14399 ( .A(n14157), .B(n14158), .Z(n14156) );
  XOR U14400 ( .A(n12471), .B(n14159), .Z(n14155) );
  XNOR U14401 ( .A(n12467), .B(n14160), .Z(n14150) );
  XNOR U14402 ( .A(key[715]), .B(n13123), .Z(n14160) );
  XOR U14403 ( .A(n13105), .B(n12449), .Z(n13123) );
  XOR U14404 ( .A(n14161), .B(n14162), .Z(n14096) );
  XNOR U14405 ( .A(n13105), .B(n14163), .Z(n14162) );
  XOR U14406 ( .A(n12463), .B(n14164), .Z(n14161) );
  XOR U14407 ( .A(key[712]), .B(n14165), .Z(n14164) );
  XOR U14408 ( .A(n13110), .B(n12497), .Z(n12463) );
  IV U14409 ( .A(n13103), .Z(n13110) );
  XOR U14410 ( .A(n10061), .B(n11272), .Z(n10044) );
  IV U14411 ( .A(n13693), .Z(n11272) );
  XNOR U14412 ( .A(n13826), .B(n13772), .Z(n13693) );
  XNOR U14413 ( .A(n13837), .B(n14166), .Z(n13772) );
  XNOR U14414 ( .A(n14167), .B(n13731), .Z(n14166) );
  ANDN U14415 ( .B(n13852), .A(n14168), .Z(n13731) );
  XNOR U14416 ( .A(n13854), .B(n13733), .Z(n13852) );
  NOR U14417 ( .A(n13854), .B(n14169), .Z(n14167) );
  XNOR U14418 ( .A(n13729), .B(n14170), .Z(n13837) );
  XNOR U14419 ( .A(n14171), .B(n14172), .Z(n14170) );
  NAND U14420 ( .A(n14173), .B(n13858), .Z(n14172) );
  XNOR U14421 ( .A(n13779), .B(n13771), .Z(n13826) );
  XOR U14422 ( .A(n13729), .B(n14174), .Z(n13771) );
  XNOR U14423 ( .A(n13839), .B(n14175), .Z(n14174) );
  NANDN U14424 ( .A(n14176), .B(n14177), .Z(n14175) );
  OR U14425 ( .A(n14178), .B(n14179), .Z(n13839) );
  XOR U14426 ( .A(n14180), .B(n14171), .Z(n13729) );
  OR U14427 ( .A(n14181), .B(n14182), .Z(n14171) );
  ANDN U14428 ( .B(n14183), .A(n14184), .Z(n14180) );
  IV U14429 ( .A(n13848), .Z(n13779) );
  XOR U14430 ( .A(n13832), .B(n14185), .Z(n13848) );
  XOR U14431 ( .A(n14186), .B(n13845), .Z(n14185) );
  OR U14432 ( .A(n14187), .B(n14178), .Z(n13845) );
  XNOR U14433 ( .A(n13841), .B(n14176), .Z(n14178) );
  NOR U14434 ( .A(n14188), .B(n14176), .Z(n14186) );
  XOR U14435 ( .A(n14189), .B(n13856), .Z(n13832) );
  OR U14436 ( .A(n14181), .B(n14190), .Z(n13856) );
  XNOR U14437 ( .A(n14183), .B(n13858), .Z(n14181) );
  XNOR U14438 ( .A(n14176), .B(n13733), .Z(n13858) );
  XOR U14439 ( .A(n14191), .B(n14192), .Z(n13733) );
  NANDN U14440 ( .A(n14193), .B(n14194), .Z(n14192) );
  XNOR U14441 ( .A(n14195), .B(n14196), .Z(n14176) );
  OR U14442 ( .A(n14193), .B(n14197), .Z(n14196) );
  XOR U14443 ( .A(n13841), .B(n13854), .Z(n14183) );
  XOR U14444 ( .A(n14199), .B(n14191), .Z(n13854) );
  NANDN U14445 ( .A(n14200), .B(n14201), .Z(n14191) );
  ANDN U14446 ( .B(n14202), .A(n14203), .Z(n14199) );
  NANDN U14447 ( .A(n14200), .B(n14205), .Z(n14195) );
  XOR U14448 ( .A(n14206), .B(n14193), .Z(n14200) );
  XNOR U14449 ( .A(n14207), .B(n14208), .Z(n14193) );
  XOR U14450 ( .A(n14209), .B(n14202), .Z(n14208) );
  XNOR U14451 ( .A(n14210), .B(n14211), .Z(n14207) );
  XNOR U14452 ( .A(n14212), .B(n14213), .Z(n14211) );
  ANDN U14453 ( .B(n14202), .A(n14214), .Z(n14212) );
  IV U14454 ( .A(n14215), .Z(n14202) );
  ANDN U14455 ( .B(n14206), .A(n14214), .Z(n14204) );
  IV U14456 ( .A(n14210), .Z(n14214) );
  IV U14457 ( .A(n14203), .Z(n14206) );
  XNOR U14458 ( .A(n14209), .B(n14216), .Z(n14203) );
  XOR U14459 ( .A(n14217), .B(n14213), .Z(n14216) );
  NAND U14460 ( .A(n14205), .B(n14201), .Z(n14213) );
  XNOR U14461 ( .A(n14194), .B(n14215), .Z(n14201) );
  XOR U14462 ( .A(n14218), .B(n14219), .Z(n14215) );
  XOR U14463 ( .A(n14220), .B(n14221), .Z(n14219) );
  XOR U14464 ( .A(n14222), .B(n14223), .Z(n14221) );
  XOR U14465 ( .A(n14177), .B(n14224), .Z(n14218) );
  XNOR U14466 ( .A(n14225), .B(n14226), .Z(n14224) );
  ANDN U14467 ( .B(n13842), .A(n13847), .Z(n14225) );
  XNOR U14468 ( .A(n14210), .B(n14197), .Z(n14205) );
  XOR U14469 ( .A(n14227), .B(n14228), .Z(n14210) );
  XNOR U14470 ( .A(n14229), .B(n14223), .Z(n14228) );
  XOR U14471 ( .A(n14230), .B(n14231), .Z(n14223) );
  XNOR U14472 ( .A(n14232), .B(n14233), .Z(n14231) );
  NAND U14473 ( .A(n13859), .B(n14173), .Z(n14233) );
  XNOR U14474 ( .A(n14234), .B(n14235), .Z(n14227) );
  ANDN U14475 ( .B(n13853), .A(n14169), .Z(n14234) );
  ANDN U14476 ( .B(n14194), .A(n14197), .Z(n14217) );
  XOR U14477 ( .A(n14197), .B(n14194), .Z(n14209) );
  XNOR U14478 ( .A(n14236), .B(n14237), .Z(n14194) );
  XNOR U14479 ( .A(n14230), .B(n14238), .Z(n14237) );
  XNOR U14480 ( .A(n13842), .B(n14229), .Z(n14238) );
  XNOR U14481 ( .A(n14239), .B(n14240), .Z(n14236) );
  XNOR U14482 ( .A(n14241), .B(n14226), .Z(n14240) );
  OR U14483 ( .A(n14179), .B(n14187), .Z(n14226) );
  XNOR U14484 ( .A(n14239), .B(n14222), .Z(n14187) );
  XNOR U14485 ( .A(n13842), .B(n14177), .Z(n14179) );
  ANDN U14486 ( .B(n14177), .A(n14188), .Z(n14241) );
  IV U14487 ( .A(n14222), .Z(n14188) );
  XOR U14488 ( .A(n14242), .B(n14243), .Z(n14197) );
  XOR U14489 ( .A(n14230), .B(n14220), .Z(n14243) );
  XOR U14490 ( .A(n14244), .B(n13836), .Z(n14220) );
  XOR U14491 ( .A(n14245), .B(n14232), .Z(n14230) );
  OR U14492 ( .A(n14190), .B(n14182), .Z(n14232) );
  XOR U14493 ( .A(n14184), .B(n14173), .Z(n14182) );
  XOR U14494 ( .A(n14244), .B(n14177), .Z(n14173) );
  XOR U14495 ( .A(n14246), .B(n14247), .Z(n14177) );
  XNOR U14496 ( .A(n14169), .B(n14248), .Z(n14247) );
  XNOR U14497 ( .A(n14198), .B(n13859), .Z(n14190) );
  XNOR U14498 ( .A(n13836), .B(n14222), .Z(n13859) );
  XOR U14499 ( .A(n14249), .B(n14250), .Z(n14222) );
  XNOR U14500 ( .A(n14251), .B(n14252), .Z(n14250) );
  XOR U14501 ( .A(n14239), .B(n14253), .Z(n14249) );
  ANDN U14502 ( .B(n14198), .A(n14184), .Z(n14245) );
  XOR U14503 ( .A(n14169), .B(n13842), .Z(n14184) );
  XOR U14504 ( .A(n14251), .B(n14254), .Z(n13842) );
  XOR U14505 ( .A(n14255), .B(n14256), .Z(n14254) );
  XOR U14506 ( .A(n14257), .B(n14258), .Z(n14251) );
  XNOR U14507 ( .A(n14259), .B(n14260), .Z(n14258) );
  XOR U14508 ( .A(n13212), .B(n14261), .Z(n14257) );
  XNOR U14509 ( .A(key[676]), .B(n13213), .Z(n14261) );
  XNOR U14510 ( .A(n14262), .B(n14263), .Z(n13213) );
  XOR U14511 ( .A(n14264), .B(n12585), .Z(n13212) );
  XOR U14512 ( .A(n14229), .B(n14265), .Z(n14242) );
  XNOR U14513 ( .A(n14266), .B(n14235), .Z(n14265) );
  OR U14514 ( .A(n13851), .B(n14168), .Z(n14235) );
  XOR U14515 ( .A(n14169), .B(n14244), .Z(n14168) );
  XNOR U14516 ( .A(n13853), .B(n14268), .Z(n13851) );
  ANDN U14517 ( .B(n14244), .A(n13836), .Z(n14266) );
  XOR U14518 ( .A(n14267), .B(n14256), .Z(n13836) );
  IV U14519 ( .A(n13734), .Z(n14244) );
  XNOR U14520 ( .A(n14248), .B(n14268), .Z(n13734) );
  XOR U14521 ( .A(n14169), .B(n13853), .Z(n14229) );
  XNOR U14522 ( .A(n14253), .B(n14268), .Z(n14169) );
  XNOR U14523 ( .A(n14267), .B(n14256), .Z(n14268) );
  IV U14524 ( .A(n14255), .Z(n14267) );
  XNOR U14525 ( .A(n14269), .B(n14270), .Z(n14255) );
  XOR U14526 ( .A(n14263), .B(n14271), .Z(n14270) );
  XNOR U14527 ( .A(key[677]), .B(n13221), .Z(n14269) );
  XNOR U14528 ( .A(n13215), .B(n12603), .Z(n13221) );
  XOR U14529 ( .A(n14272), .B(n14273), .Z(n14253) );
  XNOR U14530 ( .A(n14274), .B(n13230), .Z(n14273) );
  XOR U14531 ( .A(n13241), .B(n14275), .Z(n13230) );
  XNOR U14532 ( .A(key[679]), .B(n14276), .Z(n14272) );
  XOR U14533 ( .A(n14239), .B(n13853), .Z(n14198) );
  XNOR U14534 ( .A(n14252), .B(n14277), .Z(n13853) );
  XNOR U14535 ( .A(n14256), .B(n14246), .Z(n14277) );
  XOR U14536 ( .A(n14278), .B(n14279), .Z(n14246) );
  XOR U14537 ( .A(n12623), .B(n12620), .Z(n14279) );
  XNOR U14538 ( .A(n13255), .B(n12633), .Z(n12623) );
  XOR U14539 ( .A(key[674]), .B(n13253), .Z(n14278) );
  XOR U14540 ( .A(n14280), .B(n14281), .Z(n14256) );
  XOR U14541 ( .A(n14282), .B(n13847), .Z(n14281) );
  IV U14542 ( .A(n14239), .Z(n13847) );
  XOR U14543 ( .A(n13240), .B(n14283), .Z(n14280) );
  XNOR U14544 ( .A(key[678]), .B(n14284), .Z(n14283) );
  XOR U14545 ( .A(n12601), .B(n14274), .Z(n13240) );
  XOR U14546 ( .A(n12610), .B(n14285), .Z(n14274) );
  XNOR U14547 ( .A(n14286), .B(n12613), .Z(n12601) );
  XOR U14548 ( .A(n14287), .B(n14288), .Z(n14252) );
  XNOR U14549 ( .A(n14248), .B(n14289), .Z(n14288) );
  XNOR U14550 ( .A(n12631), .B(n14290), .Z(n14289) );
  XOR U14551 ( .A(n13234), .B(n12626), .Z(n12631) );
  XOR U14552 ( .A(n14291), .B(n14292), .Z(n14248) );
  XOR U14553 ( .A(n12611), .B(n12632), .Z(n14292) );
  XOR U14554 ( .A(n13259), .B(n12625), .Z(n12611) );
  XNOR U14555 ( .A(key[673]), .B(n14293), .Z(n14291) );
  XNOR U14556 ( .A(n13247), .B(n14294), .Z(n14287) );
  XOR U14557 ( .A(key[675]), .B(n13235), .Z(n14294) );
  XNOR U14558 ( .A(n14262), .B(n14259), .Z(n13247) );
  XOR U14559 ( .A(n14295), .B(n14296), .Z(n14239) );
  XOR U14560 ( .A(n13229), .B(n12624), .Z(n14296) );
  XOR U14561 ( .A(key[672]), .B(n14297), .Z(n14295) );
  XNOR U14562 ( .A(n13684), .B(n13766), .Z(n10061) );
  XNOR U14563 ( .A(n13760), .B(n14298), .Z(n13766) );
  XNOR U14564 ( .A(n14299), .B(n13721), .Z(n14298) );
  NOR U14565 ( .A(n13806), .B(n14300), .Z(n13721) );
  XNOR U14566 ( .A(n14301), .B(n13723), .Z(n13806) );
  NOR U14567 ( .A(n13808), .B(n14302), .Z(n14299) );
  IV U14568 ( .A(n14301), .Z(n13808) );
  XNOR U14569 ( .A(n13719), .B(n14303), .Z(n13760) );
  XNOR U14570 ( .A(n14304), .B(n14305), .Z(n14303) );
  NAND U14571 ( .A(n14306), .B(n13812), .Z(n14305) );
  XNOR U14572 ( .A(n13773), .B(n13765), .Z(n13684) );
  XOR U14573 ( .A(n13719), .B(n14307), .Z(n13765) );
  XNOR U14574 ( .A(n13762), .B(n14308), .Z(n14307) );
  NANDN U14575 ( .A(n14309), .B(n14310), .Z(n14308) );
  OR U14576 ( .A(n14311), .B(n14312), .Z(n13762) );
  XOR U14577 ( .A(n14313), .B(n14304), .Z(n13719) );
  OR U14578 ( .A(n14314), .B(n14315), .Z(n14304) );
  IV U14579 ( .A(n13802), .Z(n13773) );
  XOR U14580 ( .A(n13774), .B(n14318), .Z(n13802) );
  XOR U14581 ( .A(n14319), .B(n13715), .Z(n14318) );
  OR U14582 ( .A(n14320), .B(n14311), .Z(n13715) );
  XNOR U14583 ( .A(n13717), .B(n14309), .Z(n14311) );
  NOR U14584 ( .A(n14321), .B(n14309), .Z(n14319) );
  XOR U14585 ( .A(n14322), .B(n13810), .Z(n13774) );
  NANDN U14586 ( .A(n14314), .B(n14323), .Z(n13810) );
  XOR U14587 ( .A(n14317), .B(n13812), .Z(n14314) );
  XNOR U14588 ( .A(n14309), .B(n13723), .Z(n13812) );
  XOR U14589 ( .A(n14324), .B(n14325), .Z(n13723) );
  NANDN U14590 ( .A(n14326), .B(n14327), .Z(n14325) );
  XNOR U14591 ( .A(n14328), .B(n14329), .Z(n14309) );
  OR U14592 ( .A(n14326), .B(n14330), .Z(n14329) );
  ANDN U14593 ( .B(n14331), .A(n14317), .Z(n14322) );
  XOR U14594 ( .A(n13717), .B(n14301), .Z(n14317) );
  XNOR U14595 ( .A(n14332), .B(n14324), .Z(n14301) );
  NANDN U14596 ( .A(n14333), .B(n14334), .Z(n14324) );
  ANDN U14597 ( .B(n14335), .A(n14336), .Z(n14332) );
  NANDN U14598 ( .A(n14333), .B(n14338), .Z(n14328) );
  XOR U14599 ( .A(n14339), .B(n14326), .Z(n14333) );
  XNOR U14600 ( .A(n14340), .B(n14341), .Z(n14326) );
  XOR U14601 ( .A(n14342), .B(n14335), .Z(n14341) );
  XNOR U14602 ( .A(n14343), .B(n14344), .Z(n14340) );
  XNOR U14603 ( .A(n14345), .B(n14346), .Z(n14344) );
  ANDN U14604 ( .B(n14335), .A(n14347), .Z(n14345) );
  IV U14605 ( .A(n14348), .Z(n14335) );
  ANDN U14606 ( .B(n14339), .A(n14347), .Z(n14337) );
  IV U14607 ( .A(n14343), .Z(n14347) );
  IV U14608 ( .A(n14336), .Z(n14339) );
  XNOR U14609 ( .A(n14342), .B(n14349), .Z(n14336) );
  XOR U14610 ( .A(n14350), .B(n14346), .Z(n14349) );
  NAND U14611 ( .A(n14338), .B(n14334), .Z(n14346) );
  XNOR U14612 ( .A(n14327), .B(n14348), .Z(n14334) );
  XOR U14613 ( .A(n14351), .B(n14352), .Z(n14348) );
  XOR U14614 ( .A(n14353), .B(n14354), .Z(n14352) );
  XOR U14615 ( .A(n14355), .B(n14356), .Z(n14354) );
  XOR U14616 ( .A(n14310), .B(n14357), .Z(n14351) );
  XNOR U14617 ( .A(n14358), .B(n14359), .Z(n14357) );
  ANDN U14618 ( .B(n13764), .A(n13718), .Z(n14358) );
  XNOR U14619 ( .A(n14343), .B(n14330), .Z(n14338) );
  XOR U14620 ( .A(n14360), .B(n14361), .Z(n14343) );
  XNOR U14621 ( .A(n14362), .B(n14356), .Z(n14361) );
  XOR U14622 ( .A(n14363), .B(n14364), .Z(n14356) );
  XNOR U14623 ( .A(n14365), .B(n14366), .Z(n14364) );
  NAND U14624 ( .A(n13813), .B(n14306), .Z(n14366) );
  XNOR U14625 ( .A(n14367), .B(n14368), .Z(n14360) );
  ANDN U14626 ( .B(n13807), .A(n14302), .Z(n14367) );
  ANDN U14627 ( .B(n14327), .A(n14330), .Z(n14350) );
  XOR U14628 ( .A(n14330), .B(n14327), .Z(n14342) );
  XNOR U14629 ( .A(n14369), .B(n14370), .Z(n14327) );
  XNOR U14630 ( .A(n14363), .B(n14371), .Z(n14370) );
  XNOR U14631 ( .A(n13764), .B(n14362), .Z(n14371) );
  XNOR U14632 ( .A(n14372), .B(n14373), .Z(n14369) );
  XNOR U14633 ( .A(n14374), .B(n14359), .Z(n14373) );
  OR U14634 ( .A(n14312), .B(n14320), .Z(n14359) );
  XNOR U14635 ( .A(n14372), .B(n14355), .Z(n14320) );
  XNOR U14636 ( .A(n13764), .B(n14310), .Z(n14312) );
  ANDN U14637 ( .B(n14310), .A(n14321), .Z(n14374) );
  IV U14638 ( .A(n14355), .Z(n14321) );
  XOR U14639 ( .A(n14375), .B(n14376), .Z(n14330) );
  XOR U14640 ( .A(n14363), .B(n14353), .Z(n14376) );
  XOR U14641 ( .A(n14377), .B(n13778), .Z(n14353) );
  XOR U14642 ( .A(n14378), .B(n14365), .Z(n14363) );
  NANDN U14643 ( .A(n14315), .B(n14323), .Z(n14365) );
  XOR U14644 ( .A(n14331), .B(n13813), .Z(n14323) );
  XNOR U14645 ( .A(n13778), .B(n14355), .Z(n13813) );
  XOR U14646 ( .A(n14379), .B(n14380), .Z(n14355) );
  XNOR U14647 ( .A(n14381), .B(n14382), .Z(n14380) );
  XOR U14648 ( .A(n14372), .B(n14383), .Z(n14379) );
  XOR U14649 ( .A(n14316), .B(n14306), .Z(n14315) );
  XOR U14650 ( .A(n14377), .B(n14310), .Z(n14306) );
  XOR U14651 ( .A(n14384), .B(n14385), .Z(n14310) );
  XNOR U14652 ( .A(n14302), .B(n14386), .Z(n14385) );
  ANDN U14653 ( .B(n14331), .A(n14316), .Z(n14378) );
  XOR U14654 ( .A(n14302), .B(n13764), .Z(n14316) );
  XOR U14655 ( .A(n14381), .B(n14387), .Z(n13764) );
  XOR U14656 ( .A(n14388), .B(n14389), .Z(n14387) );
  XOR U14657 ( .A(n14390), .B(n14391), .Z(n14381) );
  XOR U14658 ( .A(n13397), .B(n14392), .Z(n14390) );
  XNOR U14659 ( .A(key[668]), .B(n13400), .Z(n14392) );
  XOR U14660 ( .A(n14393), .B(n12273), .Z(n13397) );
  XOR U14661 ( .A(n14362), .B(n14394), .Z(n14375) );
  XNOR U14662 ( .A(n14395), .B(n14368), .Z(n14394) );
  OR U14663 ( .A(n13805), .B(n14300), .Z(n14368) );
  XOR U14664 ( .A(n14302), .B(n14377), .Z(n14300) );
  XNOR U14665 ( .A(n13807), .B(n14397), .Z(n13805) );
  ANDN U14666 ( .B(n14377), .A(n13778), .Z(n14395) );
  XOR U14667 ( .A(n14396), .B(n14389), .Z(n13778) );
  IV U14668 ( .A(n13724), .Z(n14377) );
  XNOR U14669 ( .A(n14386), .B(n14397), .Z(n13724) );
  XOR U14670 ( .A(n14302), .B(n13807), .Z(n14362) );
  XNOR U14671 ( .A(n14383), .B(n14397), .Z(n14302) );
  XNOR U14672 ( .A(n14396), .B(n14389), .Z(n14397) );
  IV U14673 ( .A(n14388), .Z(n14396) );
  XNOR U14674 ( .A(n14398), .B(n14399), .Z(n14388) );
  XNOR U14675 ( .A(n14400), .B(n14401), .Z(n14399) );
  XNOR U14676 ( .A(n13417), .B(n14402), .Z(n14398) );
  XOR U14677 ( .A(key[669]), .B(n14403), .Z(n14402) );
  XOR U14678 ( .A(n14404), .B(n14405), .Z(n14383) );
  XOR U14679 ( .A(n12310), .B(n14406), .Z(n14405) );
  XNOR U14680 ( .A(key[671]), .B(n13391), .Z(n14404) );
  XOR U14681 ( .A(n14372), .B(n13807), .Z(n14331) );
  XNOR U14682 ( .A(n14382), .B(n14407), .Z(n13807) );
  XNOR U14683 ( .A(n14389), .B(n14384), .Z(n14407) );
  XOR U14684 ( .A(n14408), .B(n14409), .Z(n14384) );
  XOR U14685 ( .A(n12287), .B(n12283), .Z(n14409) );
  XOR U14686 ( .A(n14410), .B(n14411), .Z(n14408) );
  XOR U14687 ( .A(key[666]), .B(n13382), .Z(n14411) );
  XOR U14688 ( .A(n14412), .B(n14413), .Z(n14389) );
  XNOR U14689 ( .A(n14414), .B(n13718), .Z(n14413) );
  IV U14690 ( .A(n14372), .Z(n13718) );
  XNOR U14691 ( .A(n12275), .B(n14415), .Z(n14412) );
  XNOR U14692 ( .A(key[670]), .B(n13406), .Z(n14415) );
  XNOR U14693 ( .A(n13393), .B(n12268), .Z(n13406) );
  XOR U14694 ( .A(n14416), .B(n14417), .Z(n14382) );
  XNOR U14695 ( .A(n14386), .B(n14418), .Z(n14417) );
  XOR U14696 ( .A(n13371), .B(n14419), .Z(n14418) );
  XOR U14697 ( .A(n14420), .B(n14421), .Z(n14386) );
  XNOR U14698 ( .A(n14422), .B(n14423), .Z(n14421) );
  XNOR U14699 ( .A(n12298), .B(n14424), .Z(n14420) );
  XNOR U14700 ( .A(n12296), .B(n14425), .Z(n14416) );
  XOR U14701 ( .A(key[667]), .B(n13379), .Z(n14425) );
  XOR U14702 ( .A(n14393), .B(n12259), .Z(n13379) );
  XOR U14703 ( .A(n14426), .B(n14427), .Z(n14372) );
  XOR U14704 ( .A(n14428), .B(n13393), .Z(n14427) );
  IV U14705 ( .A(n14393), .Z(n13393) );
  XOR U14706 ( .A(n12270), .B(n14429), .Z(n14426) );
  XOR U14707 ( .A(key[664]), .B(n14430), .Z(n14429) );
  XOR U14708 ( .A(n13402), .B(n12311), .Z(n12270) );
  IV U14709 ( .A(n13385), .Z(n13402) );
  XOR U14710 ( .A(n11518), .B(n11532), .Z(n8355) );
  XNOR U14711 ( .A(n11565), .B(n14431), .Z(n11532) );
  XNOR U14712 ( .A(n14432), .B(n11677), .Z(n14431) );
  ANDN U14713 ( .B(n11691), .A(n14433), .Z(n11677) );
  XOR U14714 ( .A(n11689), .B(n11536), .Z(n11691) );
  ANDN U14715 ( .B(n11689), .A(n14434), .Z(n14432) );
  XNOR U14716 ( .A(n11675), .B(n14435), .Z(n11565) );
  XNOR U14717 ( .A(n14436), .B(n14437), .Z(n14435) );
  NANDN U14718 ( .A(n11695), .B(n14438), .Z(n14437) );
  XNOR U14719 ( .A(n11675), .B(n14439), .Z(n11518) );
  XOR U14720 ( .A(n14440), .B(n11567), .Z(n14439) );
  OR U14721 ( .A(n14441), .B(n11682), .Z(n11567) );
  XOR U14722 ( .A(n11569), .B(n11685), .Z(n11682) );
  ANDN U14723 ( .B(n11685), .A(n14442), .Z(n14440) );
  XOR U14724 ( .A(n14443), .B(n14436), .Z(n11675) );
  OR U14725 ( .A(n11698), .B(n14444), .Z(n14436) );
  XOR U14726 ( .A(n14445), .B(n11695), .Z(n11698) );
  XNOR U14727 ( .A(n11685), .B(n11536), .Z(n11695) );
  XOR U14728 ( .A(n14446), .B(n14447), .Z(n11536) );
  NANDN U14729 ( .A(n14448), .B(n14449), .Z(n14447) );
  XOR U14730 ( .A(n14450), .B(n14451), .Z(n11685) );
  OR U14731 ( .A(n14448), .B(n14452), .Z(n14451) );
  ANDN U14732 ( .B(n14445), .A(n14453), .Z(n14443) );
  IV U14733 ( .A(n11701), .Z(n14445) );
  XOR U14734 ( .A(n11569), .B(n11689), .Z(n11701) );
  XNOR U14735 ( .A(n14454), .B(n14446), .Z(n11689) );
  NANDN U14736 ( .A(n14455), .B(n14456), .Z(n14446) );
  ANDN U14737 ( .B(n14457), .A(n14458), .Z(n14454) );
  NANDN U14738 ( .A(n14455), .B(n14460), .Z(n14450) );
  XOR U14739 ( .A(n14461), .B(n14448), .Z(n14455) );
  XNOR U14740 ( .A(n14462), .B(n14463), .Z(n14448) );
  XOR U14741 ( .A(n14464), .B(n14457), .Z(n14463) );
  XNOR U14742 ( .A(n14465), .B(n14466), .Z(n14462) );
  XNOR U14743 ( .A(n14467), .B(n14468), .Z(n14466) );
  ANDN U14744 ( .B(n14457), .A(n14469), .Z(n14467) );
  IV U14745 ( .A(n14470), .Z(n14457) );
  ANDN U14746 ( .B(n14461), .A(n14469), .Z(n14459) );
  IV U14747 ( .A(n14465), .Z(n14469) );
  IV U14748 ( .A(n14458), .Z(n14461) );
  XNOR U14749 ( .A(n14464), .B(n14471), .Z(n14458) );
  XOR U14750 ( .A(n14472), .B(n14468), .Z(n14471) );
  NAND U14751 ( .A(n14460), .B(n14456), .Z(n14468) );
  XNOR U14752 ( .A(n14449), .B(n14470), .Z(n14456) );
  XOR U14753 ( .A(n14473), .B(n14474), .Z(n14470) );
  XOR U14754 ( .A(n14475), .B(n14476), .Z(n14474) );
  XNOR U14755 ( .A(n11684), .B(n14477), .Z(n14476) );
  XNOR U14756 ( .A(n14478), .B(n14479), .Z(n14473) );
  XNOR U14757 ( .A(n14480), .B(n14481), .Z(n14479) );
  ANDN U14758 ( .B(n11674), .A(n11570), .Z(n14480) );
  XNOR U14759 ( .A(n14465), .B(n14452), .Z(n14460) );
  XOR U14760 ( .A(n14482), .B(n14483), .Z(n14465) );
  XNOR U14761 ( .A(n14484), .B(n14477), .Z(n14483) );
  XOR U14762 ( .A(n14485), .B(n14486), .Z(n14477) );
  XNOR U14763 ( .A(n14487), .B(n14488), .Z(n14486) );
  NAND U14764 ( .A(n14438), .B(n11696), .Z(n14488) );
  XNOR U14765 ( .A(n14489), .B(n14490), .Z(n14482) );
  ANDN U14766 ( .B(n14491), .A(n14434), .Z(n14489) );
  ANDN U14767 ( .B(n14449), .A(n14452), .Z(n14472) );
  XOR U14768 ( .A(n14452), .B(n14449), .Z(n14464) );
  XNOR U14769 ( .A(n14492), .B(n14493), .Z(n14449) );
  XNOR U14770 ( .A(n14485), .B(n14494), .Z(n14493) );
  XNOR U14771 ( .A(n14484), .B(n11674), .Z(n14494) );
  XNOR U14772 ( .A(n14495), .B(n14496), .Z(n14492) );
  XNOR U14773 ( .A(n14497), .B(n14481), .Z(n14496) );
  OR U14774 ( .A(n11683), .B(n14441), .Z(n14481) );
  XNOR U14775 ( .A(n14495), .B(n14478), .Z(n14441) );
  XNOR U14776 ( .A(n11674), .B(n11684), .Z(n11683) );
  ANDN U14777 ( .B(n11684), .A(n14442), .Z(n14497) );
  XOR U14778 ( .A(n14498), .B(n14499), .Z(n14452) );
  XOR U14779 ( .A(n14485), .B(n14475), .Z(n14499) );
  XOR U14780 ( .A(n11679), .B(n11537), .Z(n14475) );
  XOR U14781 ( .A(n14500), .B(n14487), .Z(n14485) );
  NANDN U14782 ( .A(n14444), .B(n11699), .Z(n14487) );
  XOR U14783 ( .A(n11700), .B(n11696), .Z(n11699) );
  XNOR U14784 ( .A(n14491), .B(n14501), .Z(n11684) );
  XOR U14785 ( .A(n14502), .B(n14503), .Z(n14501) );
  XOR U14786 ( .A(n14453), .B(n14438), .Z(n14444) );
  XNOR U14787 ( .A(n14442), .B(n11679), .Z(n14438) );
  IV U14788 ( .A(n14478), .Z(n14442) );
  XOR U14789 ( .A(n14504), .B(n14505), .Z(n14478) );
  XOR U14790 ( .A(n14506), .B(n14507), .Z(n14505) );
  XOR U14791 ( .A(n14495), .B(n14508), .Z(n14504) );
  ANDN U14792 ( .B(n11700), .A(n14453), .Z(n14500) );
  XNOR U14793 ( .A(n14495), .B(n14509), .Z(n14453) );
  XOR U14794 ( .A(n14491), .B(n11674), .Z(n11700) );
  XNOR U14795 ( .A(n14510), .B(n14511), .Z(n11674) );
  XOR U14796 ( .A(n14512), .B(n14507), .Z(n14511) );
  XNOR U14797 ( .A(n14513), .B(n10472), .Z(n14507) );
  XNOR U14798 ( .A(n14514), .B(n14515), .Z(n10472) );
  XOR U14799 ( .A(n11408), .B(n9580), .Z(n14515) );
  XNOR U14800 ( .A(n14516), .B(n9634), .Z(n9580) );
  XNOR U14801 ( .A(n14517), .B(n9626), .Z(n11408) );
  XOR U14802 ( .A(n11419), .B(n11394), .Z(n14514) );
  XNOR U14803 ( .A(n9579), .B(n14518), .Z(n14513) );
  XOR U14804 ( .A(key[868]), .B(n11406), .Z(n14518) );
  XOR U14805 ( .A(n9612), .B(n10489), .Z(n9579) );
  XOR U14806 ( .A(n14519), .B(n14520), .Z(n10489) );
  XNOR U14807 ( .A(n14521), .B(n14522), .Z(n14520) );
  XNOR U14808 ( .A(n14523), .B(n14524), .Z(n14519) );
  XOR U14809 ( .A(n14525), .B(n14526), .Z(n14524) );
  ANDN U14810 ( .B(n14527), .A(n14528), .Z(n14526) );
  IV U14811 ( .A(n11688), .Z(n14491) );
  XOR U14812 ( .A(n14484), .B(n14529), .Z(n14498) );
  XNOR U14813 ( .A(n14530), .B(n14490), .Z(n14529) );
  OR U14814 ( .A(n11690), .B(n14433), .Z(n14490) );
  XNOR U14815 ( .A(n14509), .B(n11679), .Z(n14433) );
  XNOR U14816 ( .A(n11688), .B(n11537), .Z(n11690) );
  ANDN U14817 ( .B(n11679), .A(n11537), .Z(n14530) );
  XOR U14818 ( .A(n14510), .B(n14531), .Z(n11537) );
  XNOR U14819 ( .A(n14503), .B(n14532), .Z(n14531) );
  XOR U14820 ( .A(n14512), .B(n14510), .Z(n11679) );
  XNOR U14821 ( .A(n14434), .B(n11688), .Z(n14484) );
  XOR U14822 ( .A(n14510), .B(n14533), .Z(n11688) );
  XNOR U14823 ( .A(n14512), .B(n14506), .Z(n14533) );
  XOR U14824 ( .A(n14534), .B(n14535), .Z(n14506) );
  XNOR U14825 ( .A(n14536), .B(n10485), .Z(n14535) );
  XNOR U14826 ( .A(n11402), .B(n9591), .Z(n10485) );
  XOR U14827 ( .A(n14537), .B(n14538), .Z(n9591) );
  XOR U14828 ( .A(n14539), .B(n14540), .Z(n14538) );
  XNOR U14829 ( .A(n14541), .B(n14542), .Z(n14537) );
  XOR U14830 ( .A(n14543), .B(n14544), .Z(n11402) );
  XNOR U14831 ( .A(n14545), .B(n14546), .Z(n14544) );
  XNOR U14832 ( .A(n14547), .B(n14548), .Z(n14543) );
  XOR U14833 ( .A(key[871]), .B(n9612), .Z(n14534) );
  XNOR U14834 ( .A(n14549), .B(n14550), .Z(n14510) );
  XOR U14835 ( .A(n11394), .B(n10490), .Z(n14550) );
  XOR U14836 ( .A(n11395), .B(n9596), .Z(n10490) );
  XNOR U14837 ( .A(n14551), .B(n14552), .Z(n9596) );
  XOR U14838 ( .A(n14553), .B(n14540), .Z(n14552) );
  XNOR U14839 ( .A(n14554), .B(n14555), .Z(n14540) );
  XNOR U14840 ( .A(n14556), .B(n14557), .Z(n14555) );
  NANDN U14841 ( .A(n14558), .B(n14559), .Z(n14557) );
  XNOR U14842 ( .A(n14516), .B(n14560), .Z(n14551) );
  XOR U14843 ( .A(n14561), .B(n14562), .Z(n14560) );
  ANDN U14844 ( .B(n14563), .A(n14564), .Z(n14562) );
  XOR U14845 ( .A(n14565), .B(n14566), .Z(n11395) );
  XNOR U14846 ( .A(n14517), .B(n14546), .Z(n14566) );
  XNOR U14847 ( .A(n14567), .B(n14568), .Z(n14546) );
  XNOR U14848 ( .A(n14569), .B(n14570), .Z(n14568) );
  NANDN U14849 ( .A(n14571), .B(n14572), .Z(n14570) );
  XNOR U14850 ( .A(n14573), .B(n14574), .Z(n14565) );
  XOR U14851 ( .A(n14575), .B(n14576), .Z(n14574) );
  ANDN U14852 ( .B(n14577), .A(n14578), .Z(n14576) );
  XNOR U14853 ( .A(n14579), .B(n14580), .Z(n11394) );
  XNOR U14854 ( .A(n14581), .B(n14582), .Z(n14580) );
  XNOR U14855 ( .A(n14583), .B(n14584), .Z(n14579) );
  XOR U14856 ( .A(n14585), .B(n14586), .Z(n14584) );
  ANDN U14857 ( .B(n14587), .A(n14588), .Z(n14586) );
  XNOR U14858 ( .A(key[869]), .B(n11389), .Z(n14549) );
  XNOR U14859 ( .A(n9600), .B(n10493), .Z(n11389) );
  XOR U14860 ( .A(n14589), .B(n14590), .Z(n9600) );
  IV U14861 ( .A(n14509), .Z(n14434) );
  XOR U14862 ( .A(n14532), .B(n14591), .Z(n14509) );
  XNOR U14863 ( .A(n14502), .B(n14508), .Z(n14591) );
  XOR U14864 ( .A(n14592), .B(n14593), .Z(n14508) );
  XOR U14865 ( .A(n14503), .B(n14594), .Z(n14593) );
  XNOR U14866 ( .A(n10516), .B(n10507), .Z(n14594) );
  XOR U14867 ( .A(n9627), .B(n9632), .Z(n10507) );
  XNOR U14868 ( .A(n14595), .B(n14596), .Z(n9632) );
  XNOR U14869 ( .A(n14545), .B(n14597), .Z(n14596) );
  XOR U14870 ( .A(n14547), .B(n14598), .Z(n14595) );
  IV U14871 ( .A(n10523), .Z(n9627) );
  XNOR U14872 ( .A(n14599), .B(n14600), .Z(n10523) );
  XOR U14873 ( .A(n14542), .B(n14601), .Z(n14600) );
  XOR U14874 ( .A(n14541), .B(n14602), .Z(n14599) );
  XOR U14875 ( .A(n11419), .B(n11406), .Z(n10516) );
  XNOR U14876 ( .A(n14583), .B(n10512), .Z(n11406) );
  XNOR U14877 ( .A(n14603), .B(n14604), .Z(n14503) );
  XOR U14878 ( .A(n11381), .B(n10513), .Z(n14604) );
  XOR U14879 ( .A(n9614), .B(n9624), .Z(n10513) );
  XNOR U14880 ( .A(n14539), .B(n14605), .Z(n9624) );
  XNOR U14881 ( .A(n14541), .B(n14606), .Z(n14605) );
  XNOR U14882 ( .A(n14607), .B(n14608), .Z(n14541) );
  XNOR U14883 ( .A(n14609), .B(n14610), .Z(n14608) );
  NANDN U14884 ( .A(n14611), .B(n14559), .Z(n14610) );
  XOR U14885 ( .A(n14547), .B(n14548), .Z(n14612) );
  XNOR U14886 ( .A(n14614), .B(n14615), .Z(n14613) );
  NAND U14887 ( .A(n14616), .B(n14572), .Z(n14615) );
  XOR U14888 ( .A(n9622), .B(n10512), .Z(n11381) );
  XNOR U14889 ( .A(key[865]), .B(n10502), .Z(n14603) );
  XNOR U14890 ( .A(n9617), .B(n14618), .Z(n14592) );
  XNOR U14891 ( .A(key[867]), .B(n10520), .Z(n14618) );
  XOR U14892 ( .A(n9612), .B(n11405), .Z(n9617) );
  IV U14893 ( .A(n10475), .Z(n11405) );
  XNOR U14894 ( .A(n14523), .B(n9622), .Z(n10475) );
  XOR U14895 ( .A(n14619), .B(n14620), .Z(n9622) );
  XOR U14896 ( .A(n14621), .B(n14622), .Z(n14502) );
  XNOR U14897 ( .A(n10512), .B(n11414), .Z(n14622) );
  IV U14898 ( .A(n10521), .Z(n11414) );
  XOR U14899 ( .A(n9626), .B(n9634), .Z(n10521) );
  XOR U14900 ( .A(n14623), .B(n14606), .Z(n9634) );
  IV U14901 ( .A(n14542), .Z(n14606) );
  XNOR U14902 ( .A(n14624), .B(n14625), .Z(n14542) );
  XNOR U14903 ( .A(n14626), .B(n14627), .Z(n14625) );
  NANDN U14904 ( .A(n14628), .B(n14563), .Z(n14627) );
  XNOR U14905 ( .A(n14629), .B(n14545), .Z(n9626) );
  XOR U14906 ( .A(n14630), .B(n14631), .Z(n14545) );
  XNOR U14907 ( .A(n14632), .B(n14633), .Z(n14631) );
  NANDN U14908 ( .A(n14634), .B(n14577), .Z(n14633) );
  XNOR U14909 ( .A(n14635), .B(n14636), .Z(n10512) );
  XOR U14910 ( .A(key[866]), .B(n9619), .Z(n14621) );
  XNOR U14911 ( .A(n10520), .B(n9636), .Z(n9619) );
  XNOR U14912 ( .A(n14637), .B(n14638), .Z(n9636) );
  XNOR U14913 ( .A(n14639), .B(n14590), .Z(n14638) );
  XNOR U14914 ( .A(n14640), .B(n14641), .Z(n14590) );
  XNOR U14915 ( .A(n14642), .B(n14525), .Z(n14641) );
  ANDN U14916 ( .B(n14643), .A(n14644), .Z(n14525) );
  ANDN U14917 ( .B(n14645), .A(n14646), .Z(n14642) );
  XOR U14918 ( .A(n14647), .B(n14648), .Z(n14637) );
  XOR U14919 ( .A(n14649), .B(n14650), .Z(n10520) );
  XOR U14920 ( .A(n14651), .B(n14652), .Z(n14650) );
  IV U14921 ( .A(n14512), .Z(n14532) );
  XOR U14922 ( .A(n14653), .B(n14654), .Z(n14512) );
  XNOR U14923 ( .A(n10498), .B(n11570), .Z(n14654) );
  IV U14924 ( .A(n14495), .Z(n11570) );
  XOR U14925 ( .A(n14655), .B(n14656), .Z(n14495) );
  XNOR U14926 ( .A(n11418), .B(n9623), .Z(n14656) );
  XOR U14927 ( .A(n10515), .B(n10502), .Z(n9623) );
  XNOR U14928 ( .A(n14657), .B(n14658), .Z(n10502) );
  XOR U14929 ( .A(n14636), .B(n14659), .Z(n14658) );
  IV U14930 ( .A(n9610), .Z(n10515) );
  XOR U14931 ( .A(n14620), .B(n14660), .Z(n9610) );
  XNOR U14932 ( .A(n14647), .B(n14589), .Z(n14660) );
  IV U14933 ( .A(n14639), .Z(n14620) );
  IV U14934 ( .A(n11401), .Z(n11418) );
  XOR U14935 ( .A(n14629), .B(n14517), .Z(n11401) );
  XNOR U14936 ( .A(n14567), .B(n14661), .Z(n14517) );
  XOR U14937 ( .A(n14662), .B(n14632), .Z(n14661) );
  OR U14938 ( .A(n14663), .B(n14664), .Z(n14632) );
  XOR U14939 ( .A(n14630), .B(n14667), .Z(n14567) );
  XNOR U14940 ( .A(n14668), .B(n14669), .Z(n14667) );
  NANDN U14941 ( .A(n14670), .B(n14671), .Z(n14669) );
  XNOR U14942 ( .A(key[864]), .B(n10486), .Z(n14655) );
  XOR U14943 ( .A(n10504), .B(n11419), .Z(n10486) );
  XOR U14944 ( .A(n14516), .B(n14672), .Z(n10504) );
  XNOR U14945 ( .A(n14554), .B(n14673), .Z(n14516) );
  XOR U14946 ( .A(n14674), .B(n14626), .Z(n14673) );
  NOR U14947 ( .A(n14677), .B(n14678), .Z(n14674) );
  XNOR U14948 ( .A(n14624), .B(n14679), .Z(n14554) );
  XNOR U14949 ( .A(n14680), .B(n14681), .Z(n14679) );
  NAND U14950 ( .A(n14682), .B(n14683), .Z(n14681) );
  XOR U14951 ( .A(n11393), .B(n14536), .Z(n10498) );
  XOR U14952 ( .A(n11419), .B(n11400), .Z(n14536) );
  XNOR U14953 ( .A(n14649), .B(n14684), .Z(n11400) );
  XNOR U14954 ( .A(n14657), .B(n14582), .Z(n14684) );
  XNOR U14955 ( .A(n14685), .B(n14686), .Z(n14582) );
  XNOR U14956 ( .A(n14687), .B(n14688), .Z(n14686) );
  OR U14957 ( .A(n14689), .B(n14690), .Z(n14688) );
  XNOR U14958 ( .A(n14636), .B(n14659), .Z(n14649) );
  XOR U14959 ( .A(n14691), .B(n14692), .Z(n14659) );
  XNOR U14960 ( .A(n14693), .B(n14694), .Z(n14692) );
  OR U14961 ( .A(n14689), .B(n14695), .Z(n14694) );
  XNOR U14962 ( .A(n14696), .B(n14697), .Z(n14636) );
  XNOR U14963 ( .A(n14698), .B(n14699), .Z(n14697) );
  NAND U14964 ( .A(n14700), .B(n14587), .Z(n14699) );
  XOR U14965 ( .A(n14635), .B(n14583), .Z(n11419) );
  XNOR U14966 ( .A(n14685), .B(n14701), .Z(n14583) );
  XOR U14967 ( .A(n14702), .B(n14698), .Z(n14701) );
  ANDN U14968 ( .B(n14705), .A(n14706), .Z(n14702) );
  XNOR U14969 ( .A(n14696), .B(n14707), .Z(n14685) );
  XNOR U14970 ( .A(n14708), .B(n14709), .Z(n14707) );
  NANDN U14971 ( .A(n14710), .B(n14711), .Z(n14709) );
  XOR U14972 ( .A(n9604), .B(n9598), .Z(n11393) );
  XOR U14973 ( .A(n14548), .B(n14597), .Z(n9598) );
  XNOR U14974 ( .A(n14617), .B(n14712), .Z(n14597) );
  XNOR U14975 ( .A(n14713), .B(n14575), .Z(n14712) );
  NOR U14976 ( .A(n14664), .B(n14714), .Z(n14575) );
  XNOR U14977 ( .A(n14666), .B(n14577), .Z(n14664) );
  ANDN U14978 ( .B(n14666), .A(n14715), .Z(n14713) );
  XNOR U14979 ( .A(n14573), .B(n14716), .Z(n14617) );
  XNOR U14980 ( .A(n14717), .B(n14718), .Z(n14716) );
  OR U14981 ( .A(n14670), .B(n14719), .Z(n14718) );
  XOR U14982 ( .A(n14629), .B(n14598), .Z(n14548) );
  XOR U14983 ( .A(n14573), .B(n14720), .Z(n14598) );
  XNOR U14984 ( .A(n14614), .B(n14721), .Z(n14720) );
  NANDN U14985 ( .A(n14722), .B(n14723), .Z(n14721) );
  OR U14986 ( .A(n14724), .B(n14725), .Z(n14614) );
  XOR U14987 ( .A(n14726), .B(n14717), .Z(n14573) );
  OR U14988 ( .A(n14727), .B(n14728), .Z(n14717) );
  ANDN U14989 ( .B(n14729), .A(n14730), .Z(n14726) );
  XOR U14990 ( .A(n14732), .B(n14569), .Z(n14731) );
  OR U14991 ( .A(n14724), .B(n14733), .Z(n14569) );
  XNOR U14992 ( .A(n14572), .B(n14723), .Z(n14724) );
  ANDN U14993 ( .B(n14723), .A(n14734), .Z(n14732) );
  XNOR U14994 ( .A(n14735), .B(n14668), .Z(n14630) );
  NANDN U14995 ( .A(n14728), .B(n14736), .Z(n14668) );
  XOR U14996 ( .A(n14729), .B(n14670), .Z(n14728) );
  XNOR U14997 ( .A(n14723), .B(n14577), .Z(n14670) );
  XNOR U14998 ( .A(n14737), .B(n14738), .Z(n14577) );
  NANDN U14999 ( .A(n14739), .B(n14740), .Z(n14738) );
  XOR U15000 ( .A(n14741), .B(n14742), .Z(n14723) );
  NANDN U15001 ( .A(n14739), .B(n14743), .Z(n14742) );
  XOR U15002 ( .A(n14666), .B(n14572), .Z(n14729) );
  XNOR U15003 ( .A(n14745), .B(n14741), .Z(n14572) );
  NANDN U15004 ( .A(n14746), .B(n14747), .Z(n14741) );
  XOR U15005 ( .A(n14743), .B(n14748), .Z(n14747) );
  ANDN U15006 ( .B(n14748), .A(n14749), .Z(n14745) );
  XOR U15007 ( .A(n14750), .B(n14737), .Z(n14666) );
  ANDN U15008 ( .B(n14751), .A(n14746), .Z(n14737) );
  XNOR U15009 ( .A(n14752), .B(n14753), .Z(n14739) );
  XOR U15010 ( .A(n14754), .B(n14755), .Z(n14753) );
  XNOR U15011 ( .A(n14756), .B(n14757), .Z(n14752) );
  XNOR U15012 ( .A(n14758), .B(n14759), .Z(n14757) );
  ANDN U15013 ( .B(n14760), .A(n14755), .Z(n14758) );
  XOR U15014 ( .A(n14760), .B(n14740), .Z(n14751) );
  ANDN U15015 ( .B(n14760), .A(n14749), .Z(n14750) );
  XNOR U15016 ( .A(n14754), .B(n14761), .Z(n14749) );
  XOR U15017 ( .A(n14762), .B(n14759), .Z(n14761) );
  NAND U15018 ( .A(n14763), .B(n14764), .Z(n14759) );
  XNOR U15019 ( .A(n14756), .B(n14740), .Z(n14764) );
  IV U15020 ( .A(n14760), .Z(n14756) );
  XNOR U15021 ( .A(n14743), .B(n14755), .Z(n14763) );
  IV U15022 ( .A(n14748), .Z(n14755) );
  XOR U15023 ( .A(n14765), .B(n14766), .Z(n14748) );
  XNOR U15024 ( .A(n14767), .B(n14768), .Z(n14766) );
  XNOR U15025 ( .A(n14769), .B(n14770), .Z(n14765) );
  ANDN U15026 ( .B(n14771), .A(n14772), .Z(n14769) );
  AND U15027 ( .A(n14740), .B(n14743), .Z(n14762) );
  XNOR U15028 ( .A(n14740), .B(n14743), .Z(n14754) );
  XNOR U15029 ( .A(n14773), .B(n14774), .Z(n14743) );
  XNOR U15030 ( .A(n14775), .B(n14768), .Z(n14774) );
  XOR U15031 ( .A(n14776), .B(n14777), .Z(n14773) );
  XNOR U15032 ( .A(n14778), .B(n14770), .Z(n14777) );
  OR U15033 ( .A(n14714), .B(n14663), .Z(n14770) );
  XNOR U15034 ( .A(n14665), .B(n14809), .Z(n14663) );
  XNOR U15035 ( .A(n14715), .B(n14578), .Z(n14714) );
  ANDN U15036 ( .B(n14779), .A(n14634), .Z(n14778) );
  XNOR U15037 ( .A(n14780), .B(n14781), .Z(n14740) );
  XNOR U15038 ( .A(n14768), .B(n14782), .Z(n14781) );
  XNOR U15039 ( .A(n14616), .B(n14776), .Z(n14782) );
  XNOR U15040 ( .A(n14715), .B(n14665), .Z(n14768) );
  XNOR U15041 ( .A(n14783), .B(n14784), .Z(n14780) );
  XNOR U15042 ( .A(n14785), .B(n14786), .Z(n14784) );
  ANDN U15043 ( .B(n14787), .A(n14734), .Z(n14785) );
  XNOR U15044 ( .A(n14788), .B(n14789), .Z(n14760) );
  XNOR U15045 ( .A(n14775), .B(n14790), .Z(n14789) );
  XNOR U15046 ( .A(n14791), .B(n14767), .Z(n14790) );
  XOR U15047 ( .A(n14776), .B(n14792), .Z(n14767) );
  XNOR U15048 ( .A(n14793), .B(n14794), .Z(n14792) );
  NANDN U15049 ( .A(n14719), .B(n14671), .Z(n14794) );
  XNOR U15050 ( .A(n14795), .B(n14793), .Z(n14776) );
  NANDN U15051 ( .A(n14727), .B(n14736), .Z(n14793) );
  XOR U15052 ( .A(n14744), .B(n14671), .Z(n14736) );
  XNOR U15053 ( .A(n14734), .B(n14809), .Z(n14671) );
  IV U15054 ( .A(n14791), .Z(n14734) );
  XOR U15055 ( .A(n14796), .B(n14719), .Z(n14727) );
  XNOR U15056 ( .A(n14779), .B(n14787), .Z(n14719) );
  IV U15057 ( .A(n14578), .Z(n14779) );
  ANDN U15058 ( .B(n14744), .A(n14730), .Z(n14795) );
  IV U15059 ( .A(n14796), .Z(n14730) );
  XOR U15060 ( .A(n14771), .B(n14616), .Z(n14796) );
  XOR U15061 ( .A(n14578), .B(n14634), .Z(n14775) );
  XOR U15062 ( .A(n14797), .B(n14798), .Z(n14634) );
  XOR U15063 ( .A(n14799), .B(n14800), .Z(n14578) );
  XOR U15064 ( .A(n14801), .B(n14798), .Z(n14800) );
  XNOR U15065 ( .A(n14722), .B(n14802), .Z(n14788) );
  XNOR U15066 ( .A(n14803), .B(n14786), .Z(n14802) );
  OR U15067 ( .A(n14725), .B(n14733), .Z(n14786) );
  XNOR U15068 ( .A(n14783), .B(n14791), .Z(n14733) );
  XOR U15069 ( .A(n14804), .B(n14805), .Z(n14791) );
  XNOR U15070 ( .A(n14806), .B(n14807), .Z(n14805) );
  XOR U15071 ( .A(n14783), .B(n14808), .Z(n14804) );
  XNOR U15072 ( .A(n14616), .B(n14787), .Z(n14725) );
  IV U15073 ( .A(n14722), .Z(n14787) );
  ANDN U15074 ( .B(n14616), .A(n14571), .Z(n14803) );
  XOR U15075 ( .A(n14806), .B(n14809), .Z(n14616) );
  XOR U15076 ( .A(n14810), .B(n14811), .Z(n14806) );
  XOR U15077 ( .A(n12584), .B(n14260), .Z(n14811) );
  XOR U15078 ( .A(n13225), .B(n14276), .Z(n14260) );
  XOR U15079 ( .A(n13211), .B(n14259), .Z(n12584) );
  XNOR U15080 ( .A(n14812), .B(n13253), .Z(n14259) );
  XNOR U15081 ( .A(n12583), .B(n14813), .Z(n14810) );
  XNOR U15082 ( .A(key[684]), .B(n13256), .Z(n14813) );
  IV U15083 ( .A(n14264), .Z(n13256) );
  XOR U15084 ( .A(n14814), .B(n13255), .Z(n14264) );
  XOR U15085 ( .A(n14815), .B(n14816), .Z(n12603) );
  XNOR U15086 ( .A(n14817), .B(n14818), .Z(n14816) );
  XNOR U15087 ( .A(n14819), .B(n14820), .Z(n14815) );
  XNOR U15088 ( .A(n14821), .B(n14822), .Z(n14820) );
  ANDN U15089 ( .B(n14823), .A(n14824), .Z(n14822) );
  XNOR U15090 ( .A(n14825), .B(n14826), .Z(n14722) );
  XOR U15091 ( .A(n14715), .B(n14799), .Z(n14826) );
  IV U15092 ( .A(n14771), .Z(n14715) );
  XOR U15093 ( .A(n14808), .B(n14809), .Z(n14771) );
  XNOR U15094 ( .A(n14797), .B(n14798), .Z(n14809) );
  IV U15095 ( .A(n14801), .Z(n14797) );
  XNOR U15096 ( .A(n14827), .B(n14828), .Z(n14801) );
  XOR U15097 ( .A(n12613), .B(n12602), .Z(n14828) );
  XNOR U15098 ( .A(n13225), .B(n14263), .Z(n12602) );
  XNOR U15099 ( .A(n14829), .B(n14830), .Z(n14263) );
  XNOR U15100 ( .A(n14812), .B(n14831), .Z(n14830) );
  XNOR U15101 ( .A(n14832), .B(n14833), .Z(n14829) );
  XOR U15102 ( .A(n14834), .B(n14835), .Z(n14833) );
  ANDN U15103 ( .B(n14836), .A(n14837), .Z(n14835) );
  XOR U15104 ( .A(n14838), .B(n14839), .Z(n13225) );
  XNOR U15105 ( .A(n14840), .B(n14841), .Z(n14839) );
  XNOR U15106 ( .A(n14842), .B(n14843), .Z(n14838) );
  XNOR U15107 ( .A(n14844), .B(n14845), .Z(n14843) );
  ANDN U15108 ( .B(n14846), .A(n14847), .Z(n14845) );
  XOR U15109 ( .A(n14848), .B(n14849), .Z(n12613) );
  XNOR U15110 ( .A(n13243), .B(n14850), .Z(n14827) );
  XNOR U15111 ( .A(key[685]), .B(n13215), .Z(n14850) );
  XOR U15112 ( .A(n14851), .B(n14852), .Z(n13215) );
  XNOR U15113 ( .A(n14814), .B(n14853), .Z(n14852) );
  XNOR U15114 ( .A(n14854), .B(n14855), .Z(n14851) );
  XOR U15115 ( .A(n14856), .B(n14857), .Z(n14855) );
  ANDN U15116 ( .B(n14858), .A(n14859), .Z(n14857) );
  XOR U15117 ( .A(n14860), .B(n14861), .Z(n14808) );
  XNOR U15118 ( .A(n13241), .B(n12597), .Z(n14861) );
  XNOR U15119 ( .A(n14285), .B(n13228), .Z(n12597) );
  XNOR U15120 ( .A(n14862), .B(n14863), .Z(n14285) );
  XNOR U15121 ( .A(n14864), .B(n14831), .Z(n14863) );
  XNOR U15122 ( .A(n14865), .B(n14866), .Z(n14831) );
  XNOR U15123 ( .A(n14867), .B(n14868), .Z(n14866) );
  OR U15124 ( .A(n14869), .B(n14870), .Z(n14868) );
  XNOR U15125 ( .A(n14871), .B(n14872), .Z(n14862) );
  XOR U15126 ( .A(n14873), .B(n14874), .Z(n13241) );
  XNOR U15127 ( .A(n14875), .B(n14853), .Z(n14873) );
  XNOR U15128 ( .A(n14876), .B(n14877), .Z(n14853) );
  XNOR U15129 ( .A(n14878), .B(n14879), .Z(n14877) );
  NANDN U15130 ( .A(n14880), .B(n14881), .Z(n14879) );
  XOR U15131 ( .A(n14882), .B(n14297), .Z(n12612) );
  XOR U15132 ( .A(n14571), .B(n14772), .Z(n14744) );
  IV U15133 ( .A(n14665), .Z(n14772) );
  XNOR U15134 ( .A(n14807), .B(n14883), .Z(n14665) );
  XNOR U15135 ( .A(n14798), .B(n14825), .Z(n14883) );
  XOR U15136 ( .A(n14884), .B(n14885), .Z(n14825) );
  XOR U15137 ( .A(n12626), .B(n12632), .Z(n14885) );
  XNOR U15138 ( .A(n13237), .B(n13253), .Z(n12632) );
  XNOR U15139 ( .A(n14886), .B(n14872), .Z(n13253) );
  XNOR U15140 ( .A(n14887), .B(n14888), .Z(n12626) );
  XOR U15141 ( .A(n14848), .B(n14889), .Z(n14887) );
  XOR U15142 ( .A(n14890), .B(n14891), .Z(n14848) );
  XOR U15143 ( .A(n14892), .B(n14821), .Z(n14891) );
  OR U15144 ( .A(n14893), .B(n14894), .Z(n14821) );
  ANDN U15145 ( .B(n14895), .A(n14896), .Z(n14892) );
  XNOR U15146 ( .A(n13248), .B(n14897), .Z(n14884) );
  XNOR U15147 ( .A(key[682]), .B(n13255), .Z(n14897) );
  XOR U15148 ( .A(n14898), .B(n14899), .Z(n13255) );
  XOR U15149 ( .A(n14900), .B(n14901), .Z(n14798) );
  XOR U15150 ( .A(n14282), .B(n14571), .Z(n14901) );
  XNOR U15151 ( .A(n14882), .B(n13228), .Z(n14282) );
  XNOR U15152 ( .A(n14902), .B(n14903), .Z(n13228) );
  XNOR U15153 ( .A(n14841), .B(n14904), .Z(n14902) );
  XNOR U15154 ( .A(n14905), .B(n14906), .Z(n14841) );
  XNOR U15155 ( .A(n14907), .B(n14908), .Z(n14906) );
  NANDN U15156 ( .A(n14909), .B(n14910), .Z(n14908) );
  IV U15157 ( .A(n14276), .Z(n14882) );
  XOR U15158 ( .A(n12607), .B(n14911), .Z(n14900) );
  XNOR U15159 ( .A(key[686]), .B(n14286), .Z(n14911) );
  IV U15160 ( .A(n13223), .Z(n14286) );
  XNOR U15161 ( .A(n14875), .B(n14912), .Z(n13223) );
  XOR U15162 ( .A(n14271), .B(n12596), .Z(n12607) );
  XNOR U15163 ( .A(n14297), .B(n14275), .Z(n12596) );
  XNOR U15164 ( .A(n14913), .B(n14888), .Z(n14275) );
  XOR U15165 ( .A(n14914), .B(n14915), .Z(n14888) );
  XNOR U15166 ( .A(n14818), .B(n14849), .Z(n14913) );
  XNOR U15167 ( .A(n14916), .B(n14917), .Z(n14818) );
  XNOR U15168 ( .A(n14918), .B(n14919), .Z(n14917) );
  NANDN U15169 ( .A(n14920), .B(n14921), .Z(n14919) );
  XNOR U15170 ( .A(n14284), .B(n13243), .Z(n14271) );
  XOR U15171 ( .A(n14922), .B(n14904), .Z(n13243) );
  IV U15172 ( .A(n13222), .Z(n14284) );
  XNOR U15173 ( .A(n14871), .B(n14923), .Z(n13222) );
  XOR U15174 ( .A(n14924), .B(n14925), .Z(n14807) );
  XNOR U15175 ( .A(n14290), .B(n14926), .Z(n14925) );
  XOR U15176 ( .A(n12618), .B(n14799), .Z(n14926) );
  XNOR U15177 ( .A(n14927), .B(n14928), .Z(n14799) );
  XNOR U15178 ( .A(n12633), .B(n12624), .Z(n14928) );
  XOR U15179 ( .A(n13260), .B(n13252), .Z(n12624) );
  IV U15180 ( .A(n14293), .Z(n13260) );
  XNOR U15181 ( .A(n14864), .B(n14929), .Z(n14293) );
  XNOR U15182 ( .A(n14871), .B(n14930), .Z(n14929) );
  XOR U15183 ( .A(n14931), .B(n14932), .Z(n14871) );
  XNOR U15184 ( .A(n14933), .B(n14934), .Z(n14927) );
  XNOR U15185 ( .A(key[681]), .B(n13259), .Z(n14934) );
  XOR U15186 ( .A(n14935), .B(n14936), .Z(n13259) );
  XNOR U15187 ( .A(n14875), .B(n14937), .Z(n14936) );
  XNOR U15188 ( .A(n14898), .B(n14938), .Z(n14875) );
  XNOR U15189 ( .A(n14297), .B(n12585), .Z(n12618) );
  XNOR U15190 ( .A(n14819), .B(n12633), .Z(n12585) );
  XOR U15191 ( .A(n14939), .B(n14914), .Z(n12633) );
  XNOR U15192 ( .A(n14819), .B(n14939), .Z(n14297) );
  XNOR U15193 ( .A(n14916), .B(n14940), .Z(n14819) );
  XOR U15194 ( .A(n14941), .B(n14942), .Z(n14940) );
  ANDN U15195 ( .B(n14943), .A(n14896), .Z(n14941) );
  IV U15196 ( .A(n14944), .Z(n14896) );
  XNOR U15197 ( .A(n14945), .B(n14946), .Z(n14916) );
  XNOR U15198 ( .A(n14947), .B(n14948), .Z(n14946) );
  NAND U15199 ( .A(n14949), .B(n14950), .Z(n14948) );
  XNOR U15200 ( .A(n14276), .B(n13211), .Z(n14290) );
  XOR U15201 ( .A(n14842), .B(n13237), .Z(n13211) );
  IV U15202 ( .A(n14933), .Z(n13237) );
  XNOR U15203 ( .A(n14951), .B(n14952), .Z(n14933) );
  XNOR U15204 ( .A(n12620), .B(n14953), .Z(n14924) );
  XNOR U15205 ( .A(key[683]), .B(n13234), .Z(n14953) );
  XOR U15206 ( .A(n14954), .B(n14874), .Z(n13234) );
  XOR U15207 ( .A(n14899), .B(n14935), .Z(n14874) );
  XOR U15208 ( .A(n14955), .B(n14956), .Z(n14935) );
  XNOR U15209 ( .A(n14957), .B(n14958), .Z(n14956) );
  NANDN U15210 ( .A(n14959), .B(n14881), .Z(n14958) );
  IV U15211 ( .A(n14937), .Z(n14899) );
  XOR U15212 ( .A(n14960), .B(n14961), .Z(n14937) );
  XOR U15213 ( .A(n14962), .B(n14963), .Z(n14961) );
  NANDN U15214 ( .A(n14964), .B(n14858), .Z(n14963) );
  XOR U15215 ( .A(n14938), .B(n14912), .Z(n14954) );
  XNOR U15216 ( .A(n14955), .B(n14965), .Z(n14912) );
  XNOR U15217 ( .A(n14966), .B(n14856), .Z(n14965) );
  ANDN U15218 ( .B(n14967), .A(n14968), .Z(n14856) );
  NOR U15219 ( .A(n14969), .B(n14970), .Z(n14966) );
  XNOR U15220 ( .A(n14854), .B(n14971), .Z(n14955) );
  XNOR U15221 ( .A(n14972), .B(n14973), .Z(n14971) );
  NANDN U15222 ( .A(n14974), .B(n14975), .Z(n14973) );
  XNOR U15223 ( .A(n14854), .B(n14976), .Z(n14938) );
  XNOR U15224 ( .A(n14957), .B(n14977), .Z(n14976) );
  NANDN U15225 ( .A(n14978), .B(n14979), .Z(n14977) );
  OR U15226 ( .A(n14980), .B(n14981), .Z(n14957) );
  XOR U15227 ( .A(n14982), .B(n14972), .Z(n14854) );
  NANDN U15228 ( .A(n14983), .B(n14984), .Z(n14972) );
  ANDN U15229 ( .B(n14985), .A(n14986), .Z(n14982) );
  XOR U15230 ( .A(n13235), .B(n13248), .Z(n12620) );
  XOR U15231 ( .A(n14987), .B(n14903), .Z(n13248) );
  XNOR U15232 ( .A(n14952), .B(n14988), .Z(n14903) );
  IV U15233 ( .A(n14989), .Z(n14952) );
  XOR U15234 ( .A(n14922), .B(n14990), .Z(n14987) );
  XOR U15235 ( .A(n14991), .B(n14992), .Z(n14922) );
  XOR U15236 ( .A(n14993), .B(n14844), .Z(n14992) );
  OR U15237 ( .A(n14994), .B(n14995), .Z(n14844) );
  ANDN U15238 ( .B(n14996), .A(n14997), .Z(n14993) );
  XNOR U15239 ( .A(n14998), .B(n14999), .Z(n13235) );
  XNOR U15240 ( .A(n14872), .B(n14864), .Z(n14999) );
  XNOR U15241 ( .A(n15000), .B(n15001), .Z(n14864) );
  XNOR U15242 ( .A(n15002), .B(n15003), .Z(n15001) );
  NANDN U15243 ( .A(n14869), .B(n15004), .Z(n15003) );
  IV U15244 ( .A(n14930), .Z(n14872) );
  XOR U15245 ( .A(n15005), .B(n15006), .Z(n14930) );
  XOR U15246 ( .A(n15007), .B(n15008), .Z(n15006) );
  NANDN U15247 ( .A(n15009), .B(n14836), .Z(n15008) );
  XOR U15248 ( .A(n14931), .B(n14923), .Z(n14998) );
  XNOR U15249 ( .A(n15000), .B(n15010), .Z(n14923) );
  XNOR U15250 ( .A(n15011), .B(n14834), .Z(n15010) );
  ANDN U15251 ( .B(n15012), .A(n15013), .Z(n14834) );
  NOR U15252 ( .A(n15014), .B(n15015), .Z(n15011) );
  XNOR U15253 ( .A(n14832), .B(n15016), .Z(n15000) );
  XNOR U15254 ( .A(n15017), .B(n15018), .Z(n15016) );
  NAND U15255 ( .A(n15019), .B(n15020), .Z(n15018) );
  XNOR U15256 ( .A(n14832), .B(n15021), .Z(n14931) );
  XNOR U15257 ( .A(n15002), .B(n15022), .Z(n15021) );
  NANDN U15258 ( .A(n15023), .B(n15024), .Z(n15022) );
  OR U15259 ( .A(n15025), .B(n15026), .Z(n15002) );
  XOR U15260 ( .A(n15027), .B(n15017), .Z(n14832) );
  OR U15261 ( .A(n15028), .B(n15029), .Z(n15017) );
  ANDN U15262 ( .B(n15030), .A(n15031), .Z(n15027) );
  IV U15263 ( .A(n14783), .Z(n14571) );
  XOR U15264 ( .A(n15032), .B(n15033), .Z(n14783) );
  XNOR U15265 ( .A(n14915), .B(n15034), .Z(n12625) );
  XNOR U15266 ( .A(n14849), .B(n14914), .Z(n15034) );
  XOR U15267 ( .A(n14945), .B(n15035), .Z(n14914) );
  XNOR U15268 ( .A(n14942), .B(n15036), .Z(n15035) );
  NANDN U15269 ( .A(n15037), .B(n14823), .Z(n15036) );
  OR U15270 ( .A(n15038), .B(n14893), .Z(n14942) );
  XNOR U15271 ( .A(n14944), .B(n14823), .Z(n14893) );
  XNOR U15272 ( .A(n14939), .B(n14889), .Z(n14849) );
  XNOR U15273 ( .A(n14817), .B(n15039), .Z(n14889) );
  XNOR U15274 ( .A(n15040), .B(n15041), .Z(n15039) );
  NANDN U15275 ( .A(n15042), .B(n15043), .Z(n15041) );
  XOR U15276 ( .A(n14945), .B(n15044), .Z(n14939) );
  XOR U15277 ( .A(n15045), .B(n14918), .Z(n15044) );
  OR U15278 ( .A(n15046), .B(n15047), .Z(n14918) );
  ANDN U15279 ( .B(n15043), .A(n15048), .Z(n15045) );
  XOR U15280 ( .A(n15049), .B(n14947), .Z(n14945) );
  OR U15281 ( .A(n15050), .B(n15051), .Z(n14947) );
  NOR U15282 ( .A(n15052), .B(n15053), .Z(n15049) );
  XOR U15283 ( .A(n14890), .B(n15054), .Z(n14915) );
  XNOR U15284 ( .A(n15040), .B(n15055), .Z(n15054) );
  NANDN U15285 ( .A(n15056), .B(n14921), .Z(n15055) );
  OR U15286 ( .A(n15046), .B(n15057), .Z(n15040) );
  XNOR U15287 ( .A(n14921), .B(n15043), .Z(n15046) );
  XOR U15288 ( .A(n14817), .B(n15058), .Z(n14890) );
  XNOR U15289 ( .A(n15059), .B(n15060), .Z(n15058) );
  NAND U15290 ( .A(n15061), .B(n14949), .Z(n15060) );
  XOR U15291 ( .A(n15062), .B(n15059), .Z(n14817) );
  NANDN U15292 ( .A(n15050), .B(n15063), .Z(n15059) );
  XOR U15293 ( .A(n15052), .B(n14949), .Z(n15050) );
  XOR U15294 ( .A(n15043), .B(n14823), .Z(n14949) );
  XOR U15295 ( .A(n15064), .B(n15065), .Z(n14823) );
  NANDN U15296 ( .A(n15066), .B(n15067), .Z(n15065) );
  XOR U15297 ( .A(n15068), .B(n15069), .Z(n15043) );
  NANDN U15298 ( .A(n15066), .B(n15070), .Z(n15069) );
  ANDN U15299 ( .B(n15071), .A(n15052), .Z(n15062) );
  XNOR U15300 ( .A(n14944), .B(n14921), .Z(n15052) );
  XNOR U15301 ( .A(n15072), .B(n15068), .Z(n14921) );
  NANDN U15302 ( .A(n15073), .B(n15074), .Z(n15068) );
  XOR U15303 ( .A(n15070), .B(n15075), .Z(n15074) );
  ANDN U15304 ( .B(n15075), .A(n15076), .Z(n15072) );
  XNOR U15305 ( .A(n15077), .B(n15064), .Z(n14944) );
  NANDN U15306 ( .A(n15073), .B(n15078), .Z(n15064) );
  XOR U15307 ( .A(n15079), .B(n15067), .Z(n15078) );
  XNOR U15308 ( .A(n15080), .B(n15081), .Z(n15066) );
  XOR U15309 ( .A(n15082), .B(n15083), .Z(n15081) );
  XNOR U15310 ( .A(n15084), .B(n15085), .Z(n15080) );
  XNOR U15311 ( .A(n15086), .B(n15087), .Z(n15085) );
  ANDN U15312 ( .B(n15079), .A(n15083), .Z(n15086) );
  ANDN U15313 ( .B(n15079), .A(n15076), .Z(n15077) );
  XNOR U15314 ( .A(n15082), .B(n15088), .Z(n15076) );
  XOR U15315 ( .A(n15089), .B(n15087), .Z(n15088) );
  NAND U15316 ( .A(n15090), .B(n15091), .Z(n15087) );
  XNOR U15317 ( .A(n15084), .B(n15067), .Z(n15091) );
  IV U15318 ( .A(n15079), .Z(n15084) );
  XNOR U15319 ( .A(n15070), .B(n15083), .Z(n15090) );
  IV U15320 ( .A(n15075), .Z(n15083) );
  XOR U15321 ( .A(n15092), .B(n15093), .Z(n15075) );
  XNOR U15322 ( .A(n15094), .B(n15095), .Z(n15093) );
  XNOR U15323 ( .A(n15096), .B(n15097), .Z(n15092) );
  ANDN U15324 ( .B(n14943), .A(n15098), .Z(n15096) );
  AND U15325 ( .A(n15067), .B(n15070), .Z(n15089) );
  XNOR U15326 ( .A(n15067), .B(n15070), .Z(n15082) );
  XNOR U15327 ( .A(n15099), .B(n15100), .Z(n15070) );
  XNOR U15328 ( .A(n15101), .B(n15095), .Z(n15100) );
  XOR U15329 ( .A(n15102), .B(n15103), .Z(n15099) );
  XNOR U15330 ( .A(n15104), .B(n15097), .Z(n15103) );
  OR U15331 ( .A(n14894), .B(n15038), .Z(n15097) );
  XNOR U15332 ( .A(n14943), .B(n15105), .Z(n15038) );
  XNOR U15333 ( .A(n15098), .B(n14824), .Z(n14894) );
  ANDN U15334 ( .B(n15106), .A(n15037), .Z(n15104) );
  XNOR U15335 ( .A(n15107), .B(n15108), .Z(n15067) );
  XNOR U15336 ( .A(n15095), .B(n15109), .Z(n15108) );
  XOR U15337 ( .A(n15056), .B(n15102), .Z(n15109) );
  XNOR U15338 ( .A(n14943), .B(n15098), .Z(n15095) );
  XOR U15339 ( .A(n14920), .B(n15110), .Z(n15107) );
  XNOR U15340 ( .A(n15111), .B(n15112), .Z(n15110) );
  ANDN U15341 ( .B(n15113), .A(n15048), .Z(n15111) );
  XNOR U15342 ( .A(n15114), .B(n15115), .Z(n15079) );
  XNOR U15343 ( .A(n15101), .B(n15116), .Z(n15115) );
  XNOR U15344 ( .A(n15042), .B(n15094), .Z(n15116) );
  XOR U15345 ( .A(n15102), .B(n15117), .Z(n15094) );
  XNOR U15346 ( .A(n15118), .B(n15119), .Z(n15117) );
  NAND U15347 ( .A(n14950), .B(n15061), .Z(n15119) );
  XNOR U15348 ( .A(n15120), .B(n15118), .Z(n15102) );
  NANDN U15349 ( .A(n15051), .B(n15063), .Z(n15118) );
  XOR U15350 ( .A(n15071), .B(n15061), .Z(n15063) );
  XNOR U15351 ( .A(n15113), .B(n14824), .Z(n15061) );
  XOR U15352 ( .A(n15053), .B(n14950), .Z(n15051) );
  XNOR U15353 ( .A(n15048), .B(n15105), .Z(n14950) );
  ANDN U15354 ( .B(n15071), .A(n15053), .Z(n15120) );
  XOR U15355 ( .A(n14920), .B(n14943), .Z(n15053) );
  XNOR U15356 ( .A(n15121), .B(n15122), .Z(n14943) );
  XNOR U15357 ( .A(n15123), .B(n15124), .Z(n15122) );
  XOR U15358 ( .A(n15105), .B(n15106), .Z(n15101) );
  IV U15359 ( .A(n14824), .Z(n15106) );
  XOR U15360 ( .A(n15125), .B(n15126), .Z(n14824) );
  XNOR U15361 ( .A(n15127), .B(n15124), .Z(n15126) );
  IV U15362 ( .A(n15037), .Z(n15105) );
  XOR U15363 ( .A(n15124), .B(n15128), .Z(n15037) );
  XNOR U15364 ( .A(n15129), .B(n15130), .Z(n15114) );
  XNOR U15365 ( .A(n15131), .B(n15112), .Z(n15130) );
  OR U15366 ( .A(n15057), .B(n15047), .Z(n15112) );
  XNOR U15367 ( .A(n14920), .B(n15048), .Z(n15047) );
  IV U15368 ( .A(n15129), .Z(n15048) );
  XOR U15369 ( .A(n15056), .B(n15113), .Z(n15057) );
  IV U15370 ( .A(n15042), .Z(n15113) );
  XOR U15371 ( .A(n14895), .B(n15132), .Z(n15042) );
  XNOR U15372 ( .A(n15127), .B(n15121), .Z(n15132) );
  XOR U15373 ( .A(n15133), .B(n15134), .Z(n15121) );
  XNOR U15374 ( .A(n15135), .B(n15136), .Z(n15134) );
  XNOR U15375 ( .A(n15137), .B(n15138), .Z(n15133) );
  XNOR U15376 ( .A(key[618]), .B(n15139), .Z(n15138) );
  NOR U15377 ( .A(n15056), .B(n14920), .Z(n15131) );
  XOR U15378 ( .A(n15140), .B(n15141), .Z(n15129) );
  XNOR U15379 ( .A(n15142), .B(n15143), .Z(n15141) );
  XNOR U15380 ( .A(n14920), .B(n15123), .Z(n15140) );
  XOR U15381 ( .A(n15144), .B(n15145), .Z(n15123) );
  XNOR U15382 ( .A(n15146), .B(n15147), .Z(n15145) );
  XOR U15383 ( .A(n15127), .B(n15148), .Z(n15147) );
  XOR U15384 ( .A(n15149), .B(n15150), .Z(n15127) );
  XNOR U15385 ( .A(n15151), .B(n15152), .Z(n15150) );
  XNOR U15386 ( .A(n15153), .B(n15154), .Z(n15149) );
  XOR U15387 ( .A(key[617]), .B(n15155), .Z(n15154) );
  XNOR U15388 ( .A(n15156), .B(n15157), .Z(n15144) );
  XNOR U15389 ( .A(key[619]), .B(n15158), .Z(n15157) );
  IV U15390 ( .A(n15098), .Z(n14895) );
  XOR U15391 ( .A(n15125), .B(n15159), .Z(n15098) );
  XOR U15392 ( .A(n15124), .B(n15143), .Z(n15159) );
  XNOR U15393 ( .A(n15160), .B(n15161), .Z(n15143) );
  XNOR U15394 ( .A(n15162), .B(n15163), .Z(n15161) );
  XOR U15395 ( .A(key[623]), .B(n15164), .Z(n15160) );
  XOR U15396 ( .A(n15125), .B(n15165), .Z(n15056) );
  XOR U15397 ( .A(n15124), .B(n15142), .Z(n15165) );
  XNOR U15398 ( .A(n15166), .B(n15167), .Z(n15142) );
  XNOR U15399 ( .A(n15168), .B(n15169), .Z(n15167) );
  XNOR U15400 ( .A(n15170), .B(n15171), .Z(n15166) );
  XOR U15401 ( .A(key[620]), .B(n15172), .Z(n15171) );
  XOR U15402 ( .A(n15173), .B(n15174), .Z(n15124) );
  XNOR U15403 ( .A(n15175), .B(n15176), .Z(n15174) );
  XNOR U15404 ( .A(n15177), .B(n15178), .Z(n15173) );
  XOR U15405 ( .A(key[622]), .B(n14920), .Z(n15178) );
  XNOR U15406 ( .A(n15179), .B(n15180), .Z(n14920) );
  XNOR U15407 ( .A(n15181), .B(n15182), .Z(n15180) );
  XNOR U15408 ( .A(n15183), .B(n15184), .Z(n15179) );
  XOR U15409 ( .A(key[616]), .B(n15185), .Z(n15184) );
  IV U15410 ( .A(n15128), .Z(n15125) );
  XOR U15411 ( .A(n15186), .B(n15187), .Z(n15128) );
  XNOR U15412 ( .A(n15188), .B(n15189), .Z(n15187) );
  XOR U15413 ( .A(n15190), .B(n15191), .Z(n15186) );
  XOR U15414 ( .A(key[621]), .B(n15192), .Z(n15191) );
  XOR U15415 ( .A(n14988), .B(n15193), .Z(n13252) );
  XNOR U15416 ( .A(n14904), .B(n14989), .Z(n15193) );
  XOR U15417 ( .A(n15194), .B(n15195), .Z(n14989) );
  XNOR U15418 ( .A(n15196), .B(n15197), .Z(n15195) );
  NANDN U15419 ( .A(n15198), .B(n14846), .Z(n15197) );
  XOR U15420 ( .A(n14951), .B(n14990), .Z(n14904) );
  XNOR U15421 ( .A(n14840), .B(n15199), .Z(n14990) );
  XNOR U15422 ( .A(n15200), .B(n15201), .Z(n15199) );
  NANDN U15423 ( .A(n15202), .B(n15203), .Z(n15201) );
  IV U15424 ( .A(n15204), .Z(n14951) );
  XOR U15425 ( .A(n14991), .B(n15205), .Z(n14988) );
  XNOR U15426 ( .A(n15200), .B(n15206), .Z(n15205) );
  NANDN U15427 ( .A(n15207), .B(n14910), .Z(n15206) );
  OR U15428 ( .A(n15208), .B(n15209), .Z(n15200) );
  XOR U15429 ( .A(n14840), .B(n15210), .Z(n14991) );
  XNOR U15430 ( .A(n15211), .B(n15212), .Z(n15210) );
  NAND U15431 ( .A(n15213), .B(n15214), .Z(n15212) );
  XOR U15432 ( .A(n15215), .B(n15211), .Z(n14840) );
  NANDN U15433 ( .A(n15216), .B(n15217), .Z(n15211) );
  ANDN U15434 ( .B(n15218), .A(n15219), .Z(n15215) );
  XNOR U15435 ( .A(n13229), .B(n15220), .Z(n15032) );
  XNOR U15436 ( .A(key[680]), .B(n14276), .Z(n15220) );
  XOR U15437 ( .A(n14842), .B(n15204), .Z(n14276) );
  XOR U15438 ( .A(n15194), .B(n15221), .Z(n15204) );
  XOR U15439 ( .A(n15222), .B(n14907), .Z(n15221) );
  OR U15440 ( .A(n15223), .B(n15208), .Z(n14907) );
  XNOR U15441 ( .A(n14910), .B(n15203), .Z(n15208) );
  ANDN U15442 ( .B(n15203), .A(n15224), .Z(n15222) );
  XNOR U15443 ( .A(n14905), .B(n15225), .Z(n14842) );
  XOR U15444 ( .A(n15226), .B(n15196), .Z(n15225) );
  OR U15445 ( .A(n15227), .B(n14994), .Z(n15196) );
  XNOR U15446 ( .A(n15228), .B(n14846), .Z(n14994) );
  ANDN U15447 ( .B(n15229), .A(n14997), .Z(n15226) );
  IV U15448 ( .A(n15228), .Z(n14997) );
  XNOR U15449 ( .A(n15194), .B(n15230), .Z(n14905) );
  XNOR U15450 ( .A(n15231), .B(n15232), .Z(n15230) );
  NAND U15451 ( .A(n15214), .B(n15233), .Z(n15232) );
  XOR U15452 ( .A(n15234), .B(n15231), .Z(n15194) );
  OR U15453 ( .A(n15235), .B(n15216), .Z(n15231) );
  XOR U15454 ( .A(n15219), .B(n15214), .Z(n15216) );
  XOR U15455 ( .A(n15203), .B(n14846), .Z(n15214) );
  XOR U15456 ( .A(n15236), .B(n15237), .Z(n14846) );
  NANDN U15457 ( .A(n15238), .B(n15239), .Z(n15237) );
  XOR U15458 ( .A(n15240), .B(n15241), .Z(n15203) );
  NANDN U15459 ( .A(n15238), .B(n15242), .Z(n15241) );
  NOR U15460 ( .A(n15219), .B(n15243), .Z(n15234) );
  XNOR U15461 ( .A(n15228), .B(n14910), .Z(n15219) );
  XNOR U15462 ( .A(n15244), .B(n15240), .Z(n14910) );
  NANDN U15463 ( .A(n15245), .B(n15246), .Z(n15240) );
  XOR U15464 ( .A(n15242), .B(n15247), .Z(n15246) );
  ANDN U15465 ( .B(n15247), .A(n15248), .Z(n15244) );
  XNOR U15466 ( .A(n15249), .B(n15236), .Z(n15228) );
  NANDN U15467 ( .A(n15245), .B(n15250), .Z(n15236) );
  XOR U15468 ( .A(n15251), .B(n15239), .Z(n15250) );
  XNOR U15469 ( .A(n15252), .B(n15253), .Z(n15238) );
  XOR U15470 ( .A(n15254), .B(n15255), .Z(n15253) );
  XNOR U15471 ( .A(n15256), .B(n15257), .Z(n15252) );
  XNOR U15472 ( .A(n15258), .B(n15259), .Z(n15257) );
  ANDN U15473 ( .B(n15251), .A(n15255), .Z(n15258) );
  ANDN U15474 ( .B(n15251), .A(n15248), .Z(n15249) );
  XNOR U15475 ( .A(n15254), .B(n15260), .Z(n15248) );
  XOR U15476 ( .A(n15261), .B(n15259), .Z(n15260) );
  NAND U15477 ( .A(n15262), .B(n15263), .Z(n15259) );
  XNOR U15478 ( .A(n15256), .B(n15239), .Z(n15263) );
  IV U15479 ( .A(n15251), .Z(n15256) );
  XNOR U15480 ( .A(n15242), .B(n15255), .Z(n15262) );
  IV U15481 ( .A(n15247), .Z(n15255) );
  XOR U15482 ( .A(n15264), .B(n15265), .Z(n15247) );
  XNOR U15483 ( .A(n15266), .B(n15267), .Z(n15265) );
  XNOR U15484 ( .A(n15268), .B(n15269), .Z(n15264) );
  ANDN U15485 ( .B(n15229), .A(n15270), .Z(n15268) );
  AND U15486 ( .A(n15239), .B(n15242), .Z(n15261) );
  XNOR U15487 ( .A(n15239), .B(n15242), .Z(n15254) );
  XNOR U15488 ( .A(n15271), .B(n15272), .Z(n15242) );
  XNOR U15489 ( .A(n15273), .B(n15267), .Z(n15272) );
  XOR U15490 ( .A(n15274), .B(n15275), .Z(n15271) );
  XNOR U15491 ( .A(n15276), .B(n15269), .Z(n15275) );
  OR U15492 ( .A(n14995), .B(n15227), .Z(n15269) );
  XNOR U15493 ( .A(n15229), .B(n15277), .Z(n15227) );
  XNOR U15494 ( .A(n15270), .B(n14847), .Z(n14995) );
  ANDN U15495 ( .B(n15278), .A(n15198), .Z(n15276) );
  XNOR U15496 ( .A(n15279), .B(n15280), .Z(n15239) );
  XNOR U15497 ( .A(n15267), .B(n15281), .Z(n15280) );
  XOR U15498 ( .A(n15207), .B(n15274), .Z(n15281) );
  XNOR U15499 ( .A(n15229), .B(n15270), .Z(n15267) );
  XOR U15500 ( .A(n14909), .B(n15282), .Z(n15279) );
  XNOR U15501 ( .A(n15283), .B(n15284), .Z(n15282) );
  ANDN U15502 ( .B(n15285), .A(n15224), .Z(n15283) );
  XNOR U15503 ( .A(n15286), .B(n15287), .Z(n15251) );
  XNOR U15504 ( .A(n15273), .B(n15288), .Z(n15287) );
  XNOR U15505 ( .A(n15202), .B(n15266), .Z(n15288) );
  XOR U15506 ( .A(n15274), .B(n15289), .Z(n15266) );
  XNOR U15507 ( .A(n15290), .B(n15291), .Z(n15289) );
  NAND U15508 ( .A(n15233), .B(n15213), .Z(n15291) );
  XNOR U15509 ( .A(n15292), .B(n15290), .Z(n15274) );
  NANDN U15510 ( .A(n15235), .B(n15217), .Z(n15290) );
  XOR U15511 ( .A(n15218), .B(n15213), .Z(n15217) );
  XNOR U15512 ( .A(n15285), .B(n14847), .Z(n15213) );
  XOR U15513 ( .A(n15243), .B(n15233), .Z(n15235) );
  XNOR U15514 ( .A(n15224), .B(n15277), .Z(n15233) );
  ANDN U15515 ( .B(n15218), .A(n15243), .Z(n15292) );
  XOR U15516 ( .A(n14909), .B(n15229), .Z(n15243) );
  XNOR U15517 ( .A(n15293), .B(n15294), .Z(n15229) );
  XNOR U15518 ( .A(n15295), .B(n15296), .Z(n15294) );
  XOR U15519 ( .A(n15277), .B(n15278), .Z(n15273) );
  IV U15520 ( .A(n14847), .Z(n15278) );
  XOR U15521 ( .A(n15297), .B(n15298), .Z(n14847) );
  XNOR U15522 ( .A(n15299), .B(n15296), .Z(n15298) );
  IV U15523 ( .A(n15198), .Z(n15277) );
  XOR U15524 ( .A(n15296), .B(n15300), .Z(n15198) );
  XNOR U15525 ( .A(n15301), .B(n15302), .Z(n15286) );
  XNOR U15526 ( .A(n15303), .B(n15284), .Z(n15302) );
  OR U15527 ( .A(n15209), .B(n15223), .Z(n15284) );
  XNOR U15528 ( .A(n14909), .B(n15224), .Z(n15223) );
  IV U15529 ( .A(n15301), .Z(n15224) );
  XOR U15530 ( .A(n15207), .B(n15285), .Z(n15209) );
  IV U15531 ( .A(n15202), .Z(n15285) );
  XOR U15532 ( .A(n14996), .B(n15304), .Z(n15202) );
  XNOR U15533 ( .A(n15299), .B(n15293), .Z(n15304) );
  XOR U15534 ( .A(n15305), .B(n15306), .Z(n15293) );
  XNOR U15535 ( .A(n15307), .B(n15308), .Z(n15306) );
  XNOR U15536 ( .A(key[578]), .B(n15309), .Z(n15305) );
  IV U15537 ( .A(n15270), .Z(n14996) );
  XOR U15538 ( .A(n15297), .B(n15310), .Z(n15270) );
  XOR U15539 ( .A(n15296), .B(n15311), .Z(n15310) );
  NOR U15540 ( .A(n15207), .B(n14909), .Z(n15303) );
  XOR U15541 ( .A(n15297), .B(n15312), .Z(n15207) );
  XOR U15542 ( .A(n15296), .B(n15313), .Z(n15312) );
  XOR U15543 ( .A(n15314), .B(n15315), .Z(n15296) );
  XNOR U15544 ( .A(n15316), .B(n15317), .Z(n15315) );
  XOR U15545 ( .A(n15318), .B(n15319), .Z(n15314) );
  XOR U15546 ( .A(key[582]), .B(n14909), .Z(n15319) );
  IV U15547 ( .A(n15300), .Z(n15297) );
  XOR U15548 ( .A(n15320), .B(n15321), .Z(n15300) );
  XNOR U15549 ( .A(n15322), .B(n15323), .Z(n15321) );
  XNOR U15550 ( .A(key[581]), .B(n15324), .Z(n15320) );
  XOR U15551 ( .A(n15325), .B(n15326), .Z(n15301) );
  XNOR U15552 ( .A(n15313), .B(n15311), .Z(n15326) );
  XNOR U15553 ( .A(n15327), .B(n15328), .Z(n15311) );
  XNOR U15554 ( .A(n15329), .B(n15330), .Z(n15328) );
  XNOR U15555 ( .A(key[583]), .B(n15331), .Z(n15327) );
  XNOR U15556 ( .A(n15332), .B(n15333), .Z(n15313) );
  XNOR U15557 ( .A(n15334), .B(n15335), .Z(n15333) );
  XNOR U15558 ( .A(n15336), .B(n15337), .Z(n15332) );
  XNOR U15559 ( .A(key[580]), .B(n15338), .Z(n15337) );
  XNOR U15560 ( .A(n14909), .B(n15295), .Z(n15325) );
  XOR U15561 ( .A(n15339), .B(n15340), .Z(n15295) );
  XNOR U15562 ( .A(n15341), .B(n15342), .Z(n15340) );
  XOR U15563 ( .A(n15299), .B(n15343), .Z(n15342) );
  XOR U15564 ( .A(n15344), .B(n15345), .Z(n15299) );
  XOR U15565 ( .A(n15346), .B(n15347), .Z(n15345) );
  XOR U15566 ( .A(key[577]), .B(n15348), .Z(n15344) );
  XOR U15567 ( .A(n15349), .B(n15350), .Z(n15339) );
  XNOR U15568 ( .A(key[579]), .B(n15351), .Z(n15350) );
  XNOR U15569 ( .A(n15352), .B(n15353), .Z(n14909) );
  XNOR U15570 ( .A(n15354), .B(n15355), .Z(n15353) );
  XOR U15571 ( .A(key[576]), .B(n15356), .Z(n15352) );
  XNOR U15572 ( .A(n13216), .B(n14262), .Z(n13229) );
  IV U15573 ( .A(n12610), .Z(n14262) );
  XOR U15574 ( .A(n14886), .B(n14812), .Z(n12610) );
  XNOR U15575 ( .A(n14865), .B(n15357), .Z(n14812) );
  XNOR U15576 ( .A(n15358), .B(n15007), .Z(n15357) );
  XNOR U15577 ( .A(n15014), .B(n14836), .Z(n15012) );
  ANDN U15578 ( .B(n15360), .A(n15014), .Z(n15358) );
  XNOR U15579 ( .A(n15005), .B(n15361), .Z(n14865) );
  XNOR U15580 ( .A(n15362), .B(n15363), .Z(n15361) );
  NAND U15581 ( .A(n15020), .B(n15364), .Z(n15363) );
  IV U15582 ( .A(n14932), .Z(n14886) );
  XNOR U15583 ( .A(n15005), .B(n15365), .Z(n14932) );
  XOR U15584 ( .A(n15366), .B(n14867), .Z(n15365) );
  OR U15585 ( .A(n15367), .B(n15025), .Z(n14867) );
  XNOR U15586 ( .A(n14869), .B(n15023), .Z(n15025) );
  NOR U15587 ( .A(n15368), .B(n15023), .Z(n15366) );
  XOR U15588 ( .A(n15369), .B(n15362), .Z(n15005) );
  OR U15589 ( .A(n15028), .B(n15370), .Z(n15362) );
  XNOR U15590 ( .A(n15030), .B(n15020), .Z(n15028) );
  XNOR U15591 ( .A(n15023), .B(n14836), .Z(n15020) );
  XOR U15592 ( .A(n15371), .B(n15372), .Z(n14836) );
  NANDN U15593 ( .A(n15373), .B(n15374), .Z(n15372) );
  XNOR U15594 ( .A(n15375), .B(n15376), .Z(n15023) );
  OR U15595 ( .A(n15373), .B(n15377), .Z(n15376) );
  XOR U15596 ( .A(n14869), .B(n15014), .Z(n15030) );
  XOR U15597 ( .A(n15379), .B(n15371), .Z(n15014) );
  NANDN U15598 ( .A(n15380), .B(n15381), .Z(n15371) );
  ANDN U15599 ( .B(n15382), .A(n15383), .Z(n15379) );
  NANDN U15600 ( .A(n15380), .B(n15385), .Z(n15375) );
  XOR U15601 ( .A(n15386), .B(n15373), .Z(n15380) );
  XNOR U15602 ( .A(n15387), .B(n15388), .Z(n15373) );
  XOR U15603 ( .A(n15389), .B(n15382), .Z(n15388) );
  XNOR U15604 ( .A(n15390), .B(n15391), .Z(n15387) );
  XNOR U15605 ( .A(n15392), .B(n15393), .Z(n15391) );
  ANDN U15606 ( .B(n15382), .A(n15394), .Z(n15392) );
  IV U15607 ( .A(n15395), .Z(n15382) );
  ANDN U15608 ( .B(n15386), .A(n15394), .Z(n15384) );
  IV U15609 ( .A(n15390), .Z(n15394) );
  IV U15610 ( .A(n15383), .Z(n15386) );
  XNOR U15611 ( .A(n15389), .B(n15396), .Z(n15383) );
  XOR U15612 ( .A(n15397), .B(n15393), .Z(n15396) );
  NAND U15613 ( .A(n15385), .B(n15381), .Z(n15393) );
  XNOR U15614 ( .A(n15374), .B(n15395), .Z(n15381) );
  XOR U15615 ( .A(n15398), .B(n15399), .Z(n15395) );
  XOR U15616 ( .A(n15400), .B(n15401), .Z(n15399) );
  XOR U15617 ( .A(n15402), .B(n15403), .Z(n15401) );
  XOR U15618 ( .A(n15024), .B(n15404), .Z(n15398) );
  XNOR U15619 ( .A(n15405), .B(n15406), .Z(n15404) );
  ANDN U15620 ( .B(n15004), .A(n14870), .Z(n15405) );
  XNOR U15621 ( .A(n15390), .B(n15377), .Z(n15385) );
  XOR U15622 ( .A(n15407), .B(n15408), .Z(n15390) );
  XNOR U15623 ( .A(n15409), .B(n15403), .Z(n15408) );
  XOR U15624 ( .A(n15410), .B(n15411), .Z(n15403) );
  XNOR U15625 ( .A(n15412), .B(n15413), .Z(n15411) );
  NAND U15626 ( .A(n15364), .B(n15019), .Z(n15413) );
  XNOR U15627 ( .A(n15414), .B(n15415), .Z(n15407) );
  ANDN U15628 ( .B(n15360), .A(n15015), .Z(n15414) );
  ANDN U15629 ( .B(n15374), .A(n15377), .Z(n15397) );
  XOR U15630 ( .A(n15377), .B(n15374), .Z(n15389) );
  XNOR U15631 ( .A(n15416), .B(n15417), .Z(n15374) );
  XNOR U15632 ( .A(n15410), .B(n15418), .Z(n15417) );
  XNOR U15633 ( .A(n15004), .B(n15409), .Z(n15418) );
  XNOR U15634 ( .A(n15419), .B(n15420), .Z(n15416) );
  XNOR U15635 ( .A(n15421), .B(n15406), .Z(n15420) );
  OR U15636 ( .A(n15026), .B(n15367), .Z(n15406) );
  XNOR U15637 ( .A(n15419), .B(n15402), .Z(n15367) );
  XNOR U15638 ( .A(n15004), .B(n15024), .Z(n15026) );
  ANDN U15639 ( .B(n15024), .A(n15368), .Z(n15421) );
  IV U15640 ( .A(n15402), .Z(n15368) );
  XOR U15641 ( .A(n15422), .B(n15423), .Z(n15377) );
  XOR U15642 ( .A(n15410), .B(n15400), .Z(n15423) );
  XOR U15643 ( .A(n15424), .B(n15009), .Z(n15400) );
  XOR U15644 ( .A(n15425), .B(n15412), .Z(n15410) );
  OR U15645 ( .A(n15370), .B(n15029), .Z(n15412) );
  XOR U15646 ( .A(n15031), .B(n15019), .Z(n15029) );
  XOR U15647 ( .A(n15424), .B(n15024), .Z(n15019) );
  XOR U15648 ( .A(n15426), .B(n15427), .Z(n15024) );
  XNOR U15649 ( .A(n15015), .B(n15428), .Z(n15427) );
  XNOR U15650 ( .A(n15378), .B(n15364), .Z(n15370) );
  XNOR U15651 ( .A(n15009), .B(n15402), .Z(n15364) );
  XOR U15652 ( .A(n15429), .B(n15430), .Z(n15402) );
  XNOR U15653 ( .A(n15431), .B(n15432), .Z(n15430) );
  XOR U15654 ( .A(n15419), .B(n15433), .Z(n15429) );
  ANDN U15655 ( .B(n15378), .A(n15031), .Z(n15425) );
  XOR U15656 ( .A(n15015), .B(n15004), .Z(n15031) );
  XOR U15657 ( .A(n15431), .B(n15434), .Z(n15004) );
  XOR U15658 ( .A(n15435), .B(n15436), .Z(n15434) );
  XOR U15659 ( .A(n15437), .B(n15438), .Z(n15431) );
  XOR U15660 ( .A(n15439), .B(n15440), .Z(n15438) );
  XNOR U15661 ( .A(n15441), .B(n15442), .Z(n15437) );
  XNOR U15662 ( .A(key[572]), .B(n15443), .Z(n15442) );
  XOR U15663 ( .A(n15409), .B(n15444), .Z(n15422) );
  XNOR U15664 ( .A(n15445), .B(n15415), .Z(n15444) );
  OR U15665 ( .A(n15359), .B(n15013), .Z(n15415) );
  XOR U15666 ( .A(n15015), .B(n15424), .Z(n15013) );
  XNOR U15667 ( .A(n15360), .B(n15447), .Z(n15359) );
  ANDN U15668 ( .B(n15424), .A(n15009), .Z(n15445) );
  XOR U15669 ( .A(n15446), .B(n15436), .Z(n15009) );
  IV U15670 ( .A(n14837), .Z(n15424) );
  XNOR U15671 ( .A(n15428), .B(n15447), .Z(n14837) );
  XOR U15672 ( .A(n15015), .B(n15360), .Z(n15409) );
  XNOR U15673 ( .A(n15433), .B(n15447), .Z(n15015) );
  XNOR U15674 ( .A(n15446), .B(n15436), .Z(n15447) );
  IV U15675 ( .A(n15435), .Z(n15446) );
  XNOR U15676 ( .A(n15448), .B(n15449), .Z(n15435) );
  XNOR U15677 ( .A(n15450), .B(n15451), .Z(n15449) );
  XNOR U15678 ( .A(n15452), .B(n15453), .Z(n15448) );
  XNOR U15679 ( .A(key[573]), .B(n15454), .Z(n15453) );
  XOR U15680 ( .A(n15455), .B(n15456), .Z(n15433) );
  XNOR U15681 ( .A(n15457), .B(n15458), .Z(n15456) );
  XOR U15682 ( .A(key[575]), .B(n15459), .Z(n15455) );
  XOR U15683 ( .A(n15419), .B(n15360), .Z(n15378) );
  XNOR U15684 ( .A(n15432), .B(n15460), .Z(n15360) );
  XNOR U15685 ( .A(n15436), .B(n15426), .Z(n15460) );
  XOR U15686 ( .A(n15461), .B(n15462), .Z(n15426) );
  XNOR U15687 ( .A(n15465), .B(n15466), .Z(n15461) );
  XNOR U15688 ( .A(key[570]), .B(n15467), .Z(n15466) );
  XOR U15689 ( .A(n15468), .B(n15469), .Z(n15436) );
  XOR U15690 ( .A(n15470), .B(n14870), .Z(n15469) );
  IV U15691 ( .A(n15419), .Z(n14870) );
  XNOR U15692 ( .A(n15471), .B(n15472), .Z(n15468) );
  XNOR U15693 ( .A(key[574]), .B(n15473), .Z(n15472) );
  XOR U15694 ( .A(n15474), .B(n15475), .Z(n15432) );
  XNOR U15695 ( .A(n15476), .B(n15477), .Z(n15475) );
  XOR U15696 ( .A(n15478), .B(n15479), .Z(n15477) );
  XNOR U15697 ( .A(n15480), .B(n15481), .Z(n15474) );
  XNOR U15698 ( .A(key[571]), .B(n15428), .Z(n15481) );
  XOR U15699 ( .A(n15482), .B(n15483), .Z(n15428) );
  XNOR U15700 ( .A(n15484), .B(n15485), .Z(n15483) );
  XOR U15701 ( .A(n15486), .B(n15487), .Z(n15482) );
  XNOR U15702 ( .A(key[569]), .B(n15488), .Z(n15487) );
  XOR U15703 ( .A(n15489), .B(n15490), .Z(n15419) );
  XNOR U15704 ( .A(n15491), .B(n15492), .Z(n15490) );
  XOR U15705 ( .A(n15493), .B(n15494), .Z(n15489) );
  XNOR U15706 ( .A(key[568]), .B(n15495), .Z(n15494) );
  XNOR U15707 ( .A(n14898), .B(n14814), .Z(n13216) );
  XNOR U15708 ( .A(n14876), .B(n15496), .Z(n14814) );
  XNOR U15709 ( .A(n15497), .B(n14962), .Z(n15496) );
  XNOR U15710 ( .A(n14970), .B(n14858), .Z(n14967) );
  ANDN U15711 ( .B(n15499), .A(n14970), .Z(n15497) );
  XNOR U15712 ( .A(n14960), .B(n15500), .Z(n14876) );
  XNOR U15713 ( .A(n15501), .B(n15502), .Z(n15500) );
  NANDN U15714 ( .A(n14974), .B(n15503), .Z(n15502) );
  XOR U15715 ( .A(n14960), .B(n15504), .Z(n14898) );
  XOR U15716 ( .A(n15505), .B(n14878), .Z(n15504) );
  OR U15717 ( .A(n15506), .B(n14980), .Z(n14878) );
  XNOR U15718 ( .A(n14881), .B(n14979), .Z(n14980) );
  ANDN U15719 ( .B(n14979), .A(n15507), .Z(n15505) );
  XOR U15720 ( .A(n15508), .B(n15501), .Z(n14960) );
  OR U15721 ( .A(n14983), .B(n15509), .Z(n15501) );
  XOR U15722 ( .A(n15510), .B(n14974), .Z(n14983) );
  XNOR U15723 ( .A(n14979), .B(n14858), .Z(n14974) );
  XOR U15724 ( .A(n15511), .B(n15512), .Z(n14858) );
  NANDN U15725 ( .A(n15513), .B(n15514), .Z(n15512) );
  XOR U15726 ( .A(n15515), .B(n15516), .Z(n14979) );
  NANDN U15727 ( .A(n15513), .B(n15517), .Z(n15516) );
  ANDN U15728 ( .B(n15510), .A(n15518), .Z(n15508) );
  IV U15729 ( .A(n14986), .Z(n15510) );
  XOR U15730 ( .A(n14970), .B(n14881), .Z(n14986) );
  XNOR U15731 ( .A(n15519), .B(n15515), .Z(n14881) );
  NANDN U15732 ( .A(n15520), .B(n15521), .Z(n15515) );
  XOR U15733 ( .A(n15517), .B(n15522), .Z(n15521) );
  ANDN U15734 ( .B(n15522), .A(n15523), .Z(n15519) );
  XOR U15735 ( .A(n15524), .B(n15511), .Z(n14970) );
  NANDN U15736 ( .A(n15520), .B(n15525), .Z(n15511) );
  XOR U15737 ( .A(n15526), .B(n15514), .Z(n15525) );
  XNOR U15738 ( .A(n15527), .B(n15528), .Z(n15513) );
  XOR U15739 ( .A(n15529), .B(n15530), .Z(n15528) );
  XNOR U15740 ( .A(n15531), .B(n15532), .Z(n15527) );
  XNOR U15741 ( .A(n15533), .B(n15534), .Z(n15532) );
  ANDN U15742 ( .B(n15526), .A(n15530), .Z(n15533) );
  ANDN U15743 ( .B(n15526), .A(n15523), .Z(n15524) );
  XNOR U15744 ( .A(n15529), .B(n15535), .Z(n15523) );
  XOR U15745 ( .A(n15536), .B(n15534), .Z(n15535) );
  NAND U15746 ( .A(n15537), .B(n15538), .Z(n15534) );
  XNOR U15747 ( .A(n15531), .B(n15514), .Z(n15538) );
  IV U15748 ( .A(n15526), .Z(n15531) );
  XNOR U15749 ( .A(n15517), .B(n15530), .Z(n15537) );
  IV U15750 ( .A(n15522), .Z(n15530) );
  XOR U15751 ( .A(n15539), .B(n15540), .Z(n15522) );
  XNOR U15752 ( .A(n15541), .B(n15542), .Z(n15540) );
  XNOR U15753 ( .A(n15543), .B(n15544), .Z(n15539) );
  ANDN U15754 ( .B(n15499), .A(n14969), .Z(n15543) );
  AND U15755 ( .A(n15514), .B(n15517), .Z(n15536) );
  XNOR U15756 ( .A(n15514), .B(n15517), .Z(n15529) );
  XNOR U15757 ( .A(n15545), .B(n15546), .Z(n15517) );
  XNOR U15758 ( .A(n15547), .B(n15542), .Z(n15546) );
  XOR U15759 ( .A(n15548), .B(n15549), .Z(n15545) );
  XNOR U15760 ( .A(n15550), .B(n15544), .Z(n15549) );
  OR U15761 ( .A(n14968), .B(n15498), .Z(n15544) );
  XNOR U15762 ( .A(n15499), .B(n15551), .Z(n15498) );
  XNOR U15763 ( .A(n14969), .B(n14859), .Z(n14968) );
  ANDN U15764 ( .B(n15552), .A(n14964), .Z(n15550) );
  XNOR U15765 ( .A(n15553), .B(n15554), .Z(n15514) );
  XNOR U15766 ( .A(n15542), .B(n15555), .Z(n15554) );
  XOR U15767 ( .A(n14959), .B(n15548), .Z(n15555) );
  XNOR U15768 ( .A(n15499), .B(n14969), .Z(n15542) );
  XOR U15769 ( .A(n14880), .B(n15556), .Z(n15553) );
  XNOR U15770 ( .A(n15557), .B(n15558), .Z(n15556) );
  ANDN U15771 ( .B(n15559), .A(n15507), .Z(n15557) );
  XNOR U15772 ( .A(n15560), .B(n15561), .Z(n15526) );
  XNOR U15773 ( .A(n15547), .B(n15562), .Z(n15561) );
  XNOR U15774 ( .A(n14978), .B(n15541), .Z(n15562) );
  XOR U15775 ( .A(n15548), .B(n15563), .Z(n15541) );
  XNOR U15776 ( .A(n15564), .B(n15565), .Z(n15563) );
  NAND U15777 ( .A(n15503), .B(n14975), .Z(n15565) );
  XNOR U15778 ( .A(n15566), .B(n15564), .Z(n15548) );
  NANDN U15779 ( .A(n15509), .B(n14984), .Z(n15564) );
  XOR U15780 ( .A(n14985), .B(n14975), .Z(n14984) );
  XNOR U15781 ( .A(n15559), .B(n14859), .Z(n14975) );
  XOR U15782 ( .A(n15518), .B(n15503), .Z(n15509) );
  XNOR U15783 ( .A(n15507), .B(n15551), .Z(n15503) );
  ANDN U15784 ( .B(n14985), .A(n15518), .Z(n15566) );
  XOR U15785 ( .A(n14880), .B(n15499), .Z(n15518) );
  XNOR U15786 ( .A(n15567), .B(n15568), .Z(n15499) );
  XNOR U15787 ( .A(n15569), .B(n15570), .Z(n15568) );
  XOR U15788 ( .A(n15551), .B(n15552), .Z(n15547) );
  IV U15789 ( .A(n14859), .Z(n15552) );
  XOR U15790 ( .A(n15572), .B(n15573), .Z(n14859) );
  XNOR U15791 ( .A(n15574), .B(n15570), .Z(n15573) );
  IV U15792 ( .A(n14964), .Z(n15551) );
  XOR U15793 ( .A(n15570), .B(n15575), .Z(n14964) );
  XNOR U15794 ( .A(n15576), .B(n15577), .Z(n15560) );
  XNOR U15795 ( .A(n15578), .B(n15558), .Z(n15577) );
  OR U15796 ( .A(n14981), .B(n15506), .Z(n15558) );
  XNOR U15797 ( .A(n14880), .B(n15507), .Z(n15506) );
  IV U15798 ( .A(n15576), .Z(n15507) );
  XOR U15799 ( .A(n14959), .B(n15559), .Z(n14981) );
  IV U15800 ( .A(n14978), .Z(n15559) );
  XOR U15801 ( .A(n15571), .B(n15579), .Z(n14978) );
  XNOR U15802 ( .A(n15574), .B(n15567), .Z(n15579) );
  XOR U15803 ( .A(n15580), .B(n15581), .Z(n15567) );
  XOR U15804 ( .A(n15582), .B(n15583), .Z(n15581) );
  XNOR U15805 ( .A(key[530]), .B(n15584), .Z(n15580) );
  IV U15806 ( .A(n14969), .Z(n15571) );
  XOR U15807 ( .A(n15572), .B(n15585), .Z(n14969) );
  XOR U15808 ( .A(n15570), .B(n15586), .Z(n15585) );
  NOR U15809 ( .A(n14959), .B(n14880), .Z(n15578) );
  XOR U15810 ( .A(n15572), .B(n15587), .Z(n14959) );
  XOR U15811 ( .A(n15570), .B(n15588), .Z(n15587) );
  XOR U15812 ( .A(n15589), .B(n15590), .Z(n15570) );
  XNOR U15813 ( .A(n15591), .B(n15592), .Z(n15590) );
  XOR U15814 ( .A(n15593), .B(n15594), .Z(n15589) );
  XOR U15815 ( .A(key[534]), .B(n14880), .Z(n15594) );
  IV U15816 ( .A(n15575), .Z(n15572) );
  XOR U15817 ( .A(n15595), .B(n15596), .Z(n15575) );
  XNOR U15818 ( .A(n15597), .B(n15598), .Z(n15596) );
  XOR U15819 ( .A(key[533]), .B(n15599), .Z(n15595) );
  XOR U15820 ( .A(n15600), .B(n15601), .Z(n15576) );
  XNOR U15821 ( .A(n15588), .B(n15586), .Z(n15601) );
  XNOR U15822 ( .A(n15602), .B(n15603), .Z(n15586) );
  XNOR U15823 ( .A(n15604), .B(n15605), .Z(n15603) );
  XOR U15824 ( .A(key[535]), .B(n15606), .Z(n15602) );
  XNOR U15825 ( .A(n15607), .B(n15608), .Z(n15588) );
  XNOR U15826 ( .A(n15609), .B(n15610), .Z(n15608) );
  XNOR U15827 ( .A(key[532]), .B(n15611), .Z(n15607) );
  XNOR U15828 ( .A(n14880), .B(n15569), .Z(n15600) );
  XOR U15829 ( .A(n15612), .B(n15613), .Z(n15569) );
  XNOR U15830 ( .A(n15614), .B(n15615), .Z(n15613) );
  XOR U15831 ( .A(n15574), .B(n15616), .Z(n15615) );
  XOR U15832 ( .A(n15617), .B(n15618), .Z(n15574) );
  XNOR U15833 ( .A(n15619), .B(n15620), .Z(n15618) );
  XOR U15834 ( .A(key[529]), .B(n15621), .Z(n15617) );
  XNOR U15835 ( .A(n15622), .B(n15623), .Z(n15612) );
  XOR U15836 ( .A(key[531]), .B(n15624), .Z(n15623) );
  XNOR U15837 ( .A(n15625), .B(n15626), .Z(n14880) );
  XOR U15838 ( .A(n15627), .B(n15628), .Z(n15626) );
  XOR U15839 ( .A(key[528]), .B(n15629), .Z(n15625) );
  IV U15840 ( .A(n10491), .Z(n9604) );
  XOR U15841 ( .A(n14601), .B(n14539), .Z(n10491) );
  XOR U15842 ( .A(n14623), .B(n14602), .Z(n14539) );
  XNOR U15843 ( .A(n14553), .B(n15630), .Z(n14602) );
  XNOR U15844 ( .A(n14609), .B(n15631), .Z(n15630) );
  NANDN U15845 ( .A(n15632), .B(n15633), .Z(n15631) );
  OR U15846 ( .A(n15634), .B(n15635), .Z(n14609) );
  IV U15847 ( .A(n14672), .Z(n14623) );
  XNOR U15848 ( .A(n14624), .B(n15636), .Z(n14672) );
  XOR U15849 ( .A(n15637), .B(n14556), .Z(n15636) );
  OR U15850 ( .A(n15638), .B(n15634), .Z(n14556) );
  XNOR U15851 ( .A(n14559), .B(n15633), .Z(n15634) );
  ANDN U15852 ( .B(n15633), .A(n15639), .Z(n15637) );
  XOR U15853 ( .A(n15640), .B(n14680), .Z(n14624) );
  OR U15854 ( .A(n15641), .B(n15642), .Z(n14680) );
  ANDN U15855 ( .B(n15643), .A(n15644), .Z(n15640) );
  XNOR U15856 ( .A(n14607), .B(n15645), .Z(n14601) );
  XNOR U15857 ( .A(n15646), .B(n14561), .Z(n15645) );
  ANDN U15858 ( .B(n14676), .A(n15647), .Z(n14561) );
  XNOR U15859 ( .A(n14678), .B(n14563), .Z(n14676) );
  NOR U15860 ( .A(n15648), .B(n14678), .Z(n15646) );
  XNOR U15861 ( .A(n14553), .B(n15649), .Z(n14607) );
  XNOR U15862 ( .A(n15650), .B(n15651), .Z(n15649) );
  NAND U15863 ( .A(n15652), .B(n14682), .Z(n15651) );
  XNOR U15864 ( .A(n15653), .B(n15650), .Z(n14553) );
  NANDN U15865 ( .A(n15641), .B(n15654), .Z(n15650) );
  XNOR U15866 ( .A(n15643), .B(n14682), .Z(n15641) );
  XOR U15867 ( .A(n15633), .B(n14563), .Z(n14682) );
  XOR U15868 ( .A(n15655), .B(n15656), .Z(n14563) );
  NANDN U15869 ( .A(n15657), .B(n15658), .Z(n15656) );
  XOR U15870 ( .A(n15659), .B(n15660), .Z(n15633) );
  NANDN U15871 ( .A(n15657), .B(n15661), .Z(n15660) );
  IV U15872 ( .A(n15662), .Z(n15643) );
  ANDN U15873 ( .B(n15663), .A(n15662), .Z(n15653) );
  XOR U15874 ( .A(n14678), .B(n14559), .Z(n15662) );
  XNOR U15875 ( .A(n15664), .B(n15659), .Z(n14559) );
  NANDN U15876 ( .A(n15665), .B(n15666), .Z(n15659) );
  XOR U15877 ( .A(n15661), .B(n15667), .Z(n15666) );
  ANDN U15878 ( .B(n15667), .A(n15668), .Z(n15664) );
  XOR U15879 ( .A(n15669), .B(n15655), .Z(n14678) );
  NANDN U15880 ( .A(n15665), .B(n15670), .Z(n15655) );
  XOR U15881 ( .A(n15671), .B(n15658), .Z(n15670) );
  XNOR U15882 ( .A(n15672), .B(n15673), .Z(n15657) );
  XOR U15883 ( .A(n15674), .B(n15675), .Z(n15673) );
  XNOR U15884 ( .A(n15676), .B(n15677), .Z(n15672) );
  XNOR U15885 ( .A(n15678), .B(n15679), .Z(n15677) );
  ANDN U15886 ( .B(n15671), .A(n15675), .Z(n15678) );
  ANDN U15887 ( .B(n15671), .A(n15668), .Z(n15669) );
  XNOR U15888 ( .A(n15674), .B(n15680), .Z(n15668) );
  XOR U15889 ( .A(n15681), .B(n15679), .Z(n15680) );
  NAND U15890 ( .A(n15682), .B(n15683), .Z(n15679) );
  XNOR U15891 ( .A(n15676), .B(n15658), .Z(n15683) );
  IV U15892 ( .A(n15671), .Z(n15676) );
  XNOR U15893 ( .A(n15661), .B(n15675), .Z(n15682) );
  IV U15894 ( .A(n15667), .Z(n15675) );
  XOR U15895 ( .A(n15684), .B(n15685), .Z(n15667) );
  XNOR U15896 ( .A(n15686), .B(n15687), .Z(n15685) );
  XNOR U15897 ( .A(n15688), .B(n15689), .Z(n15684) );
  NOR U15898 ( .A(n15648), .B(n14677), .Z(n15688) );
  AND U15899 ( .A(n15658), .B(n15661), .Z(n15681) );
  XNOR U15900 ( .A(n15658), .B(n15661), .Z(n15674) );
  XNOR U15901 ( .A(n15690), .B(n15691), .Z(n15661) );
  XNOR U15902 ( .A(n15692), .B(n15687), .Z(n15691) );
  XOR U15903 ( .A(n15693), .B(n15694), .Z(n15690) );
  XNOR U15904 ( .A(n15695), .B(n15689), .Z(n15694) );
  OR U15905 ( .A(n15647), .B(n14675), .Z(n15689) );
  XNOR U15906 ( .A(n14677), .B(n14628), .Z(n14675) );
  XNOR U15907 ( .A(n15648), .B(n14564), .Z(n15647) );
  ANDN U15908 ( .B(n15696), .A(n14628), .Z(n15695) );
  XNOR U15909 ( .A(n15697), .B(n15698), .Z(n15658) );
  XNOR U15910 ( .A(n15687), .B(n15699), .Z(n15698) );
  XOR U15911 ( .A(n14611), .B(n15693), .Z(n15699) );
  XNOR U15912 ( .A(n14677), .B(n15700), .Z(n15687) );
  XOR U15913 ( .A(n14558), .B(n15701), .Z(n15697) );
  XNOR U15914 ( .A(n15702), .B(n15703), .Z(n15701) );
  ANDN U15915 ( .B(n15704), .A(n15639), .Z(n15702) );
  XNOR U15916 ( .A(n15705), .B(n15706), .Z(n15671) );
  XNOR U15917 ( .A(n15692), .B(n15707), .Z(n15706) );
  XNOR U15918 ( .A(n15632), .B(n15686), .Z(n15707) );
  XOR U15919 ( .A(n15693), .B(n15708), .Z(n15686) );
  XNOR U15920 ( .A(n15709), .B(n15710), .Z(n15708) );
  NAND U15921 ( .A(n14683), .B(n15652), .Z(n15710) );
  XNOR U15922 ( .A(n15711), .B(n15709), .Z(n15693) );
  NANDN U15923 ( .A(n15642), .B(n15654), .Z(n15709) );
  XOR U15924 ( .A(n15663), .B(n15652), .Z(n15654) );
  XNOR U15925 ( .A(n15704), .B(n14564), .Z(n15652) );
  XOR U15926 ( .A(n15644), .B(n14683), .Z(n15642) );
  XNOR U15927 ( .A(n15639), .B(n15712), .Z(n14683) );
  ANDN U15928 ( .B(n15663), .A(n15644), .Z(n15711) );
  XNOR U15929 ( .A(n14558), .B(n14677), .Z(n15644) );
  XOR U15930 ( .A(n15713), .B(n15714), .Z(n14677) );
  XNOR U15931 ( .A(n15715), .B(n15716), .Z(n15714) );
  XOR U15932 ( .A(n15712), .B(n15696), .Z(n15692) );
  IV U15933 ( .A(n14564), .Z(n15696) );
  XOR U15934 ( .A(n15717), .B(n15718), .Z(n14564) );
  XOR U15935 ( .A(n15719), .B(n15716), .Z(n15718) );
  IV U15936 ( .A(n14628), .Z(n15712) );
  XOR U15937 ( .A(n15716), .B(n15720), .Z(n14628) );
  XNOR U15938 ( .A(n15721), .B(n15722), .Z(n15705) );
  XNOR U15939 ( .A(n15723), .B(n15703), .Z(n15722) );
  OR U15940 ( .A(n15635), .B(n15638), .Z(n15703) );
  XNOR U15941 ( .A(n14558), .B(n15639), .Z(n15638) );
  IV U15942 ( .A(n15721), .Z(n15639) );
  XOR U15943 ( .A(n14611), .B(n15704), .Z(n15635) );
  IV U15944 ( .A(n15632), .Z(n15704) );
  XOR U15945 ( .A(n15700), .B(n15724), .Z(n15632) );
  XNOR U15946 ( .A(n15725), .B(n15713), .Z(n15724) );
  XOR U15947 ( .A(n15726), .B(n15727), .Z(n15713) );
  XOR U15948 ( .A(n12490), .B(n14158), .Z(n15727) );
  XOR U15949 ( .A(n12467), .B(n14124), .Z(n12490) );
  XOR U15950 ( .A(n15728), .B(n15729), .Z(n12467) );
  XOR U15951 ( .A(n15730), .B(n15731), .Z(n15729) );
  XNOR U15952 ( .A(n15732), .B(n15733), .Z(n15728) );
  XNOR U15953 ( .A(key[722]), .B(n13119), .Z(n15726) );
  IV U15954 ( .A(n14126), .Z(n13119) );
  NOR U15955 ( .A(n14611), .B(n14558), .Z(n15723) );
  XOR U15956 ( .A(n15734), .B(n15735), .Z(n15721) );
  XNOR U15957 ( .A(n15736), .B(n15737), .Z(n15735) );
  XNOR U15958 ( .A(n14558), .B(n15715), .Z(n15734) );
  XOR U15959 ( .A(n15738), .B(n15739), .Z(n15715) );
  XNOR U15960 ( .A(n14154), .B(n15740), .Z(n15739) );
  XNOR U15961 ( .A(n12480), .B(n15725), .Z(n15740) );
  IV U15962 ( .A(n15719), .Z(n15725) );
  XNOR U15963 ( .A(n15741), .B(n15742), .Z(n15719) );
  XNOR U15964 ( .A(n14163), .B(n12468), .Z(n15742) );
  XOR U15965 ( .A(n14123), .B(n14158), .Z(n12468) );
  XNOR U15966 ( .A(key[721]), .B(n13127), .Z(n15741) );
  XNOR U15967 ( .A(n13121), .B(n14165), .Z(n13127) );
  IV U15968 ( .A(n12489), .Z(n14165) );
  XOR U15969 ( .A(n15743), .B(n15744), .Z(n12489) );
  XNOR U15970 ( .A(n15745), .B(n15746), .Z(n15744) );
  IV U15971 ( .A(n12499), .Z(n13121) );
  XNOR U15972 ( .A(n15747), .B(n15748), .Z(n12499) );
  XOR U15973 ( .A(n15749), .B(n15750), .Z(n15748) );
  XOR U15974 ( .A(n12497), .B(n13108), .Z(n12480) );
  XNOR U15975 ( .A(n15751), .B(n12486), .Z(n13108) );
  IV U15976 ( .A(n14123), .Z(n12486) );
  XNOR U15977 ( .A(n15752), .B(n15730), .Z(n14123) );
  XNOR U15978 ( .A(n15753), .B(n13109), .Z(n14154) );
  XNOR U15979 ( .A(n13080), .B(n15754), .Z(n15738) );
  XOR U15980 ( .A(key[723]), .B(n14124), .Z(n15754) );
  XNOR U15981 ( .A(n15755), .B(n15756), .Z(n14124) );
  XNOR U15982 ( .A(n15757), .B(n15758), .Z(n15756) );
  XNOR U15983 ( .A(n15759), .B(n15760), .Z(n15755) );
  IV U15984 ( .A(n14153), .Z(n13080) );
  XOR U15985 ( .A(n12469), .B(n12482), .Z(n14153) );
  XOR U15986 ( .A(n15761), .B(n15762), .Z(n12482) );
  XNOR U15987 ( .A(n15763), .B(n15764), .Z(n15762) );
  XOR U15988 ( .A(n15745), .B(n15765), .Z(n15761) );
  XOR U15989 ( .A(n15766), .B(n15767), .Z(n12469) );
  XNOR U15990 ( .A(n15768), .B(n15769), .Z(n15767) );
  XNOR U15991 ( .A(n15749), .B(n15750), .Z(n15766) );
  IV U15992 ( .A(n15648), .Z(n15700) );
  XOR U15993 ( .A(n15717), .B(n15770), .Z(n15648) );
  XOR U15994 ( .A(n15716), .B(n15737), .Z(n15770) );
  XNOR U15995 ( .A(n15771), .B(n15772), .Z(n15737) );
  XNOR U15996 ( .A(n15773), .B(n14145), .Z(n15772) );
  XNOR U15997 ( .A(n14135), .B(n13104), .Z(n14145) );
  XNOR U15998 ( .A(n15774), .B(n15775), .Z(n13104) );
  XNOR U15999 ( .A(n15747), .B(n15776), .Z(n15775) );
  XOR U16000 ( .A(n15777), .B(n15750), .Z(n15774) );
  XNOR U16001 ( .A(n15779), .B(n15780), .Z(n15778) );
  OR U16002 ( .A(n15781), .B(n15782), .Z(n15780) );
  IV U16003 ( .A(n12461), .Z(n14135) );
  XOR U16004 ( .A(n15784), .B(n15785), .Z(n12461) );
  XNOR U16005 ( .A(n15763), .B(n15786), .Z(n15785) );
  XOR U16006 ( .A(n15745), .B(n15746), .Z(n15784) );
  XNOR U16007 ( .A(n15787), .B(n15765), .Z(n15746) );
  XNOR U16008 ( .A(n15789), .B(n15790), .Z(n15788) );
  NANDN U16009 ( .A(n15791), .B(n15792), .Z(n15790) );
  XOR U16010 ( .A(n15717), .B(n15794), .Z(n14611) );
  XOR U16011 ( .A(n15716), .B(n15736), .Z(n15794) );
  XNOR U16012 ( .A(n15795), .B(n14147), .Z(n15736) );
  XOR U16013 ( .A(n15796), .B(n15797), .Z(n14147) );
  XNOR U16014 ( .A(n12449), .B(n13113), .Z(n15797) );
  XOR U16015 ( .A(n15798), .B(n12487), .Z(n13113) );
  XNOR U16016 ( .A(n15749), .B(n15799), .Z(n12487) );
  IV U16017 ( .A(n15777), .Z(n15749) );
  XOR U16018 ( .A(n15800), .B(n15801), .Z(n15777) );
  XOR U16019 ( .A(n15802), .B(n15803), .Z(n15801) );
  NAND U16020 ( .A(n15804), .B(n15805), .Z(n15803) );
  XOR U16021 ( .A(n15806), .B(n12471), .Z(n12449) );
  XOR U16022 ( .A(n15787), .B(n15763), .Z(n12471) );
  IV U16023 ( .A(n15743), .Z(n15763) );
  XOR U16024 ( .A(n15807), .B(n15808), .Z(n15743) );
  XOR U16025 ( .A(n15809), .B(n15810), .Z(n15808) );
  NANDN U16026 ( .A(n15811), .B(n15812), .Z(n15810) );
  XNOR U16027 ( .A(n15753), .B(n13095), .Z(n15796) );
  XNOR U16028 ( .A(n12446), .B(n15813), .Z(n15795) );
  XNOR U16029 ( .A(key[724]), .B(n13109), .Z(n15813) );
  XOR U16030 ( .A(n15814), .B(n14158), .Z(n13109) );
  XOR U16031 ( .A(n15815), .B(n15816), .Z(n14158) );
  XOR U16032 ( .A(n12497), .B(n13094), .Z(n12446) );
  XOR U16033 ( .A(n15817), .B(n15818), .Z(n13094) );
  XNOR U16034 ( .A(n15819), .B(n15820), .Z(n15818) );
  XNOR U16035 ( .A(n15751), .B(n15821), .Z(n15817) );
  XNOR U16036 ( .A(n15822), .B(n15823), .Z(n15821) );
  ANDN U16037 ( .B(n15824), .A(n15825), .Z(n15823) );
  XOR U16038 ( .A(n15826), .B(n15827), .Z(n15716) );
  XNOR U16039 ( .A(n14558), .B(n14133), .Z(n15827) );
  XOR U16040 ( .A(n13093), .B(n15773), .Z(n14133) );
  XOR U16041 ( .A(n15753), .B(n13102), .Z(n15773) );
  XNOR U16042 ( .A(n15828), .B(n15829), .Z(n13102) );
  XOR U16043 ( .A(n15830), .B(n15831), .Z(n15829) );
  XOR U16044 ( .A(n15832), .B(n15816), .Z(n15828) );
  XNOR U16045 ( .A(n12456), .B(n12475), .Z(n13093) );
  XNOR U16046 ( .A(n15764), .B(n15833), .Z(n12475) );
  XOR U16047 ( .A(n15787), .B(n15765), .Z(n15833) );
  XOR U16048 ( .A(n15834), .B(n15835), .Z(n15765) );
  XOR U16049 ( .A(n15836), .B(n15789), .Z(n15835) );
  OR U16050 ( .A(n15837), .B(n15838), .Z(n15789) );
  AND U16051 ( .A(n15839), .B(n15840), .Z(n15836) );
  XNOR U16052 ( .A(n15793), .B(n15841), .Z(n15764) );
  XNOR U16053 ( .A(n15842), .B(n15843), .Z(n15841) );
  NANDN U16054 ( .A(n15844), .B(n15845), .Z(n15843) );
  XNOR U16055 ( .A(n15834), .B(n15846), .Z(n15793) );
  XNOR U16056 ( .A(n15847), .B(n15848), .Z(n15846) );
  NANDN U16057 ( .A(n15849), .B(n15850), .Z(n15848) );
  XNOR U16058 ( .A(n15747), .B(n15769), .Z(n12456) );
  XNOR U16059 ( .A(n15783), .B(n15851), .Z(n15769) );
  XNOR U16060 ( .A(n15852), .B(n15853), .Z(n15851) );
  ANDN U16061 ( .B(n15854), .A(n15855), .Z(n15852) );
  XNOR U16062 ( .A(n15856), .B(n15857), .Z(n15783) );
  XNOR U16063 ( .A(n15858), .B(n15859), .Z(n15857) );
  NANDN U16064 ( .A(n15860), .B(n15861), .Z(n15859) );
  XNOR U16065 ( .A(n15768), .B(n15799), .Z(n15747) );
  XNOR U16066 ( .A(n15856), .B(n15862), .Z(n15768) );
  XNOR U16067 ( .A(n15779), .B(n15863), .Z(n15862) );
  NANDN U16068 ( .A(n15864), .B(n15865), .Z(n15863) );
  OR U16069 ( .A(n15866), .B(n15867), .Z(n15779) );
  XNOR U16070 ( .A(n15868), .B(n15869), .Z(n14558) );
  XOR U16071 ( .A(n13120), .B(n12496), .Z(n15869) );
  XNOR U16072 ( .A(n15753), .B(n13105), .Z(n12496) );
  XOR U16073 ( .A(n15787), .B(n15806), .Z(n13105) );
  XNOR U16074 ( .A(n15807), .B(n15870), .Z(n15787) );
  XOR U16075 ( .A(n15871), .B(n15872), .Z(n15870) );
  ANDN U16076 ( .B(n15840), .A(n15873), .Z(n15871) );
  IV U16077 ( .A(n13126), .Z(n15753) );
  XOR U16078 ( .A(n15815), .B(n15814), .Z(n13126) );
  IV U16079 ( .A(n12485), .Z(n13120) );
  XOR U16080 ( .A(n14157), .B(n14163), .Z(n12485) );
  XNOR U16081 ( .A(n15830), .B(n15874), .Z(n14163) );
  XOR U16082 ( .A(n15832), .B(n15760), .Z(n15874) );
  IV U16083 ( .A(n15816), .Z(n15760) );
  XNOR U16084 ( .A(n15875), .B(n15876), .Z(n15816) );
  XNOR U16085 ( .A(n15877), .B(n15878), .Z(n15876) );
  NANDN U16086 ( .A(n15879), .B(n15880), .Z(n15878) );
  IV U16087 ( .A(n15757), .Z(n15830) );
  XOR U16088 ( .A(n15882), .B(n15883), .Z(n15881) );
  NOR U16089 ( .A(n15884), .B(n15885), .Z(n15882) );
  IV U16090 ( .A(n12495), .Z(n14157) );
  XOR U16091 ( .A(n15732), .B(n15888), .Z(n15887) );
  XNOR U16092 ( .A(key[720]), .B(n13103), .Z(n15868) );
  XNOR U16093 ( .A(n15800), .B(n15889), .Z(n15799) );
  XOR U16094 ( .A(n15890), .B(n15891), .Z(n15889) );
  NOR U16095 ( .A(n15892), .B(n15864), .Z(n15890) );
  XNOR U16096 ( .A(n12474), .B(n15893), .Z(n15826) );
  XNOR U16097 ( .A(key[726]), .B(n14140), .Z(n15893) );
  XOR U16098 ( .A(n12497), .B(n13101), .Z(n12474) );
  XOR U16099 ( .A(n15894), .B(n15895), .Z(n13101) );
  XNOR U16100 ( .A(n15730), .B(n15820), .Z(n15895) );
  XNOR U16101 ( .A(n15896), .B(n15897), .Z(n15820) );
  XNOR U16102 ( .A(n15898), .B(n15899), .Z(n15897) );
  NANDN U16103 ( .A(n15900), .B(n15901), .Z(n15899) );
  XNOR U16104 ( .A(n15902), .B(n15903), .Z(n15730) );
  XNOR U16105 ( .A(n15904), .B(n15905), .Z(n15903) );
  NANDN U16106 ( .A(n15906), .B(n15824), .Z(n15905) );
  XNOR U16107 ( .A(n15732), .B(n15888), .Z(n15894) );
  XNOR U16108 ( .A(n15907), .B(n15908), .Z(n15732) );
  XNOR U16109 ( .A(n15909), .B(n15910), .Z(n15908) );
  NANDN U16110 ( .A(n15911), .B(n15901), .Z(n15910) );
  XOR U16111 ( .A(n15751), .B(n15912), .Z(n12497) );
  XNOR U16112 ( .A(n15896), .B(n15913), .Z(n15751) );
  XOR U16113 ( .A(n15914), .B(n15904), .Z(n15913) );
  NANDN U16114 ( .A(n15915), .B(n15916), .Z(n15904) );
  ANDN U16115 ( .B(n15917), .A(n15918), .Z(n15914) );
  XNOR U16116 ( .A(n15902), .B(n15919), .Z(n15896) );
  XNOR U16117 ( .A(n15920), .B(n15921), .Z(n15919) );
  NAND U16118 ( .A(n15922), .B(n15923), .Z(n15921) );
  IV U16119 ( .A(n15720), .Z(n15717) );
  XOR U16120 ( .A(n15924), .B(n15925), .Z(n15720) );
  XNOR U16121 ( .A(n13095), .B(n14138), .Z(n15925) );
  XNOR U16122 ( .A(n14149), .B(n13096), .Z(n14138) );
  XNOR U16123 ( .A(n15926), .B(n15927), .Z(n13096) );
  XNOR U16124 ( .A(n15798), .B(n15776), .Z(n15927) );
  XNOR U16125 ( .A(n15928), .B(n15929), .Z(n15776) );
  XNOR U16126 ( .A(n15891), .B(n15930), .Z(n15929) );
  OR U16127 ( .A(n15781), .B(n15931), .Z(n15930) );
  OR U16128 ( .A(n15932), .B(n15866), .Z(n15891) );
  XNOR U16129 ( .A(n15781), .B(n15864), .Z(n15866) );
  XNOR U16130 ( .A(n15928), .B(n15933), .Z(n15798) );
  XNOR U16131 ( .A(n15934), .B(n15802), .Z(n15933) );
  ANDN U16132 ( .B(n15854), .A(n15937), .Z(n15934) );
  XNOR U16133 ( .A(n15800), .B(n15938), .Z(n15928) );
  XNOR U16134 ( .A(n15939), .B(n15940), .Z(n15938) );
  NANDN U16135 ( .A(n15860), .B(n15941), .Z(n15940) );
  XOR U16136 ( .A(n15942), .B(n15939), .Z(n15800) );
  OR U16137 ( .A(n15943), .B(n15944), .Z(n15939) );
  ANDN U16138 ( .B(n15945), .A(n15946), .Z(n15942) );
  XNOR U16139 ( .A(n15856), .B(n15947), .Z(n15926) );
  XOR U16140 ( .A(n15853), .B(n15948), .Z(n15947) );
  ANDN U16141 ( .B(n15805), .A(n15949), .Z(n15948) );
  ANDN U16142 ( .B(n15936), .A(n15950), .Z(n15853) );
  XOR U16143 ( .A(n15854), .B(n15805), .Z(n15936) );
  XOR U16144 ( .A(n15951), .B(n15858), .Z(n15856) );
  NANDN U16145 ( .A(n15943), .B(n15952), .Z(n15858) );
  XOR U16146 ( .A(n15945), .B(n15860), .Z(n15943) );
  XOR U16147 ( .A(n15864), .B(n15805), .Z(n15860) );
  XOR U16148 ( .A(n15953), .B(n15954), .Z(n15805) );
  NANDN U16149 ( .A(n15955), .B(n15956), .Z(n15954) );
  XNOR U16150 ( .A(n15957), .B(n15958), .Z(n15864) );
  OR U16151 ( .A(n15955), .B(n15959), .Z(n15958) );
  IV U16152 ( .A(n15960), .Z(n15945) );
  ANDN U16153 ( .B(n15961), .A(n15960), .Z(n15951) );
  XOR U16154 ( .A(n15781), .B(n15854), .Z(n15960) );
  XNOR U16155 ( .A(n15962), .B(n15953), .Z(n15854) );
  NANDN U16156 ( .A(n15963), .B(n15964), .Z(n15953) );
  ANDN U16157 ( .B(n15965), .A(n15966), .Z(n15962) );
  NANDN U16158 ( .A(n15963), .B(n15968), .Z(n15957) );
  XOR U16159 ( .A(n15969), .B(n15955), .Z(n15963) );
  XNOR U16160 ( .A(n15970), .B(n15971), .Z(n15955) );
  XOR U16161 ( .A(n15972), .B(n15965), .Z(n15971) );
  XNOR U16162 ( .A(n15973), .B(n15974), .Z(n15970) );
  XNOR U16163 ( .A(n15975), .B(n15976), .Z(n15974) );
  ANDN U16164 ( .B(n15965), .A(n15977), .Z(n15975) );
  IV U16165 ( .A(n15978), .Z(n15965) );
  ANDN U16166 ( .B(n15969), .A(n15977), .Z(n15967) );
  IV U16167 ( .A(n15973), .Z(n15977) );
  IV U16168 ( .A(n15966), .Z(n15969) );
  XNOR U16169 ( .A(n15972), .B(n15979), .Z(n15966) );
  XOR U16170 ( .A(n15980), .B(n15976), .Z(n15979) );
  NAND U16171 ( .A(n15968), .B(n15964), .Z(n15976) );
  XNOR U16172 ( .A(n15956), .B(n15978), .Z(n15964) );
  XOR U16173 ( .A(n15981), .B(n15982), .Z(n15978) );
  XOR U16174 ( .A(n15983), .B(n15984), .Z(n15982) );
  XNOR U16175 ( .A(n15865), .B(n15985), .Z(n15984) );
  XNOR U16176 ( .A(n15986), .B(n15987), .Z(n15981) );
  XNOR U16177 ( .A(n15988), .B(n15989), .Z(n15987) );
  ANDN U16178 ( .B(n15990), .A(n15931), .Z(n15988) );
  XNOR U16179 ( .A(n15973), .B(n15959), .Z(n15968) );
  XOR U16180 ( .A(n15991), .B(n15992), .Z(n15973) );
  XNOR U16181 ( .A(n15993), .B(n15985), .Z(n15992) );
  XOR U16182 ( .A(n15994), .B(n15995), .Z(n15985) );
  XNOR U16183 ( .A(n15996), .B(n15997), .Z(n15995) );
  NAND U16184 ( .A(n15941), .B(n15861), .Z(n15997) );
  XNOR U16185 ( .A(n15998), .B(n15999), .Z(n15991) );
  ANDN U16186 ( .B(n16000), .A(n15937), .Z(n15998) );
  ANDN U16187 ( .B(n15956), .A(n15959), .Z(n15980) );
  XOR U16188 ( .A(n15959), .B(n15956), .Z(n15972) );
  XNOR U16189 ( .A(n16001), .B(n16002), .Z(n15956) );
  XNOR U16190 ( .A(n15994), .B(n16003), .Z(n16002) );
  XOR U16191 ( .A(n15993), .B(n15782), .Z(n16003) );
  XOR U16192 ( .A(n15931), .B(n16004), .Z(n16001) );
  XNOR U16193 ( .A(n16005), .B(n15989), .Z(n16004) );
  OR U16194 ( .A(n15867), .B(n15932), .Z(n15989) );
  XNOR U16195 ( .A(n15931), .B(n15892), .Z(n15932) );
  XOR U16196 ( .A(n15782), .B(n15865), .Z(n15867) );
  ANDN U16197 ( .B(n15865), .A(n15892), .Z(n16005) );
  XOR U16198 ( .A(n16006), .B(n16007), .Z(n15959) );
  XOR U16199 ( .A(n15994), .B(n15983), .Z(n16007) );
  XOR U16200 ( .A(n15804), .B(n15949), .Z(n15983) );
  XOR U16201 ( .A(n16008), .B(n15996), .Z(n15994) );
  NANDN U16202 ( .A(n15944), .B(n15952), .Z(n15996) );
  XOR U16203 ( .A(n15961), .B(n15861), .Z(n15952) );
  XNOR U16204 ( .A(n16000), .B(n16009), .Z(n15865) );
  XNOR U16205 ( .A(n16010), .B(n16011), .Z(n16009) );
  XOR U16206 ( .A(n15946), .B(n15941), .Z(n15944) );
  XNOR U16207 ( .A(n15892), .B(n15804), .Z(n15941) );
  IV U16208 ( .A(n15986), .Z(n15892) );
  XOR U16209 ( .A(n16012), .B(n16013), .Z(n15986) );
  XOR U16210 ( .A(n16014), .B(n16015), .Z(n16013) );
  XNOR U16211 ( .A(n15931), .B(n16016), .Z(n16012) );
  ANDN U16212 ( .B(n15961), .A(n15946), .Z(n16008) );
  XNOR U16213 ( .A(n15931), .B(n15937), .Z(n15946) );
  XOR U16214 ( .A(n15993), .B(n16017), .Z(n16006) );
  XNOR U16215 ( .A(n16018), .B(n15999), .Z(n16017) );
  OR U16216 ( .A(n15950), .B(n15935), .Z(n15999) );
  XNOR U16217 ( .A(n16019), .B(n15804), .Z(n15935) );
  XNOR U16218 ( .A(n15855), .B(n15949), .Z(n15950) );
  ANDN U16219 ( .B(n15804), .A(n15949), .Z(n16018) );
  XOR U16220 ( .A(n16020), .B(n16021), .Z(n15949) );
  XOR U16221 ( .A(n16010), .B(n16022), .Z(n16021) );
  XOR U16222 ( .A(n16023), .B(n16020), .Z(n15804) );
  XNOR U16223 ( .A(n15937), .B(n15855), .Z(n15993) );
  IV U16224 ( .A(n16019), .Z(n15937) );
  XNOR U16225 ( .A(n16011), .B(n16024), .Z(n16019) );
  XOR U16226 ( .A(n16016), .B(n16022), .Z(n16024) );
  IV U16227 ( .A(n16023), .Z(n16022) );
  XOR U16228 ( .A(n16025), .B(n16026), .Z(n16016) );
  XNOR U16229 ( .A(n16010), .B(n16027), .Z(n16026) );
  XNOR U16230 ( .A(n16028), .B(n16029), .Z(n16027) );
  XOR U16231 ( .A(n16030), .B(n16031), .Z(n16010) );
  XNOR U16232 ( .A(n15346), .B(n16032), .Z(n16031) );
  XNOR U16233 ( .A(n15309), .B(n16033), .Z(n16030) );
  XOR U16234 ( .A(key[601]), .B(n16034), .Z(n16033) );
  XOR U16235 ( .A(n15343), .B(n16035), .Z(n16025) );
  XNOR U16236 ( .A(key[603]), .B(n15351), .Z(n16035) );
  XOR U16237 ( .A(n16036), .B(n15338), .Z(n15351) );
  XOR U16238 ( .A(n16037), .B(n16038), .Z(n16011) );
  XNOR U16239 ( .A(n16039), .B(n15307), .Z(n16038) );
  XOR U16240 ( .A(n16040), .B(n16041), .Z(n16037) );
  XNOR U16241 ( .A(key[602]), .B(n16042), .Z(n16041) );
  XOR U16242 ( .A(n16000), .B(n15990), .Z(n15961) );
  IV U16243 ( .A(n15782), .Z(n15990) );
  XOR U16244 ( .A(n16020), .B(n16043), .Z(n15782) );
  XOR U16245 ( .A(n16023), .B(n16015), .Z(n16043) );
  XNOR U16246 ( .A(n16044), .B(n16045), .Z(n16015) );
  XNOR U16247 ( .A(n15334), .B(n16046), .Z(n16045) );
  XNOR U16248 ( .A(n16047), .B(n16048), .Z(n15334) );
  XNOR U16249 ( .A(n15336), .B(n16049), .Z(n16044) );
  XNOR U16250 ( .A(key[604]), .B(n16050), .Z(n16049) );
  XOR U16251 ( .A(n16036), .B(n15324), .Z(n15336) );
  IV U16252 ( .A(n15855), .Z(n16000) );
  XOR U16253 ( .A(n16020), .B(n16051), .Z(n15855) );
  XNOR U16254 ( .A(n16023), .B(n16014), .Z(n16051) );
  XOR U16255 ( .A(n16052), .B(n16053), .Z(n16014) );
  XOR U16256 ( .A(n16054), .B(n15330), .Z(n16053) );
  XOR U16257 ( .A(n16055), .B(n16056), .Z(n15330) );
  XNOR U16258 ( .A(key[607]), .B(n16057), .Z(n16052) );
  XOR U16259 ( .A(n16058), .B(n16059), .Z(n16023) );
  XOR U16260 ( .A(n15931), .B(n16060), .Z(n16059) );
  XNOR U16261 ( .A(n16061), .B(n16062), .Z(n15931) );
  XNOR U16262 ( .A(n16063), .B(n16064), .Z(n16062) );
  XNOR U16263 ( .A(n16065), .B(n16066), .Z(n16061) );
  XOR U16264 ( .A(key[600]), .B(n16067), .Z(n16066) );
  XOR U16265 ( .A(n16068), .B(n16069), .Z(n16058) );
  XNOR U16266 ( .A(key[606]), .B(n15316), .Z(n16069) );
  XNOR U16267 ( .A(n16070), .B(n15329), .Z(n15316) );
  XOR U16268 ( .A(n16036), .B(n16071), .Z(n15329) );
  XNOR U16269 ( .A(n16072), .B(n16073), .Z(n16020) );
  XOR U16270 ( .A(n16074), .B(n15322), .Z(n16073) );
  XNOR U16271 ( .A(n16075), .B(n16076), .Z(n15322) );
  XOR U16272 ( .A(n16077), .B(n16078), .Z(n16072) );
  XNOR U16273 ( .A(key[605]), .B(n16079), .Z(n16078) );
  IV U16274 ( .A(n12454), .Z(n14149) );
  XOR U16275 ( .A(n16080), .B(n16081), .Z(n12454) );
  XNOR U16276 ( .A(n15806), .B(n15786), .Z(n16081) );
  XNOR U16277 ( .A(n16082), .B(n16083), .Z(n15786) );
  XNOR U16278 ( .A(n15872), .B(n16084), .Z(n16083) );
  NANDN U16279 ( .A(n15791), .B(n16085), .Z(n16084) );
  OR U16280 ( .A(n16086), .B(n15837), .Z(n15872) );
  XOR U16281 ( .A(n15791), .B(n15840), .Z(n15837) );
  XNOR U16282 ( .A(n16082), .B(n16087), .Z(n15806) );
  XNOR U16283 ( .A(n16088), .B(n15809), .Z(n16087) );
  ANDN U16284 ( .B(n16089), .A(n16090), .Z(n15809) );
  AND U16285 ( .A(n16091), .B(n15845), .Z(n16088) );
  XNOR U16286 ( .A(n15807), .B(n16092), .Z(n16082) );
  XNOR U16287 ( .A(n16093), .B(n16094), .Z(n16092) );
  NANDN U16288 ( .A(n15849), .B(n16095), .Z(n16094) );
  XOR U16289 ( .A(n16096), .B(n16093), .Z(n15807) );
  OR U16290 ( .A(n16097), .B(n16098), .Z(n16093) );
  AND U16291 ( .A(n16099), .B(n16100), .Z(n16096) );
  XNOR U16292 ( .A(n15834), .B(n16101), .Z(n16080) );
  XNOR U16293 ( .A(n16102), .B(n15842), .Z(n16101) );
  NAND U16294 ( .A(n16089), .B(n16103), .Z(n15842) );
  XOR U16295 ( .A(n15845), .B(n15812), .Z(n16089) );
  ANDN U16296 ( .B(n15812), .A(n16104), .Z(n16102) );
  XOR U16297 ( .A(n16105), .B(n15847), .Z(n15834) );
  OR U16298 ( .A(n16097), .B(n16106), .Z(n15847) );
  XOR U16299 ( .A(n16100), .B(n15849), .Z(n16097) );
  XNOR U16300 ( .A(n15840), .B(n15812), .Z(n15849) );
  XOR U16301 ( .A(n16107), .B(n16108), .Z(n15812) );
  NANDN U16302 ( .A(n16109), .B(n16110), .Z(n16108) );
  XOR U16303 ( .A(n16111), .B(n16112), .Z(n15840) );
  OR U16304 ( .A(n16109), .B(n16113), .Z(n16112) );
  ANDN U16305 ( .B(n16100), .A(n16114), .Z(n16105) );
  XNOR U16306 ( .A(n15791), .B(n15845), .Z(n16100) );
  XNOR U16307 ( .A(n16115), .B(n16107), .Z(n15845) );
  NANDN U16308 ( .A(n16116), .B(n16117), .Z(n16107) );
  ANDN U16309 ( .B(n16118), .A(n16119), .Z(n16115) );
  NANDN U16310 ( .A(n16116), .B(n16121), .Z(n16111) );
  XOR U16311 ( .A(n16122), .B(n16109), .Z(n16116) );
  XNOR U16312 ( .A(n16123), .B(n16124), .Z(n16109) );
  XOR U16313 ( .A(n16125), .B(n16118), .Z(n16124) );
  XNOR U16314 ( .A(n16126), .B(n16127), .Z(n16123) );
  XNOR U16315 ( .A(n16128), .B(n16129), .Z(n16127) );
  ANDN U16316 ( .B(n16118), .A(n16130), .Z(n16128) );
  IV U16317 ( .A(n16131), .Z(n16118) );
  ANDN U16318 ( .B(n16122), .A(n16130), .Z(n16120) );
  IV U16319 ( .A(n16126), .Z(n16130) );
  IV U16320 ( .A(n16119), .Z(n16122) );
  XNOR U16321 ( .A(n16125), .B(n16132), .Z(n16119) );
  XOR U16322 ( .A(n16133), .B(n16129), .Z(n16132) );
  NAND U16323 ( .A(n16121), .B(n16117), .Z(n16129) );
  XNOR U16324 ( .A(n16110), .B(n16131), .Z(n16117) );
  XOR U16325 ( .A(n16134), .B(n16135), .Z(n16131) );
  XOR U16326 ( .A(n16136), .B(n16137), .Z(n16135) );
  XOR U16327 ( .A(n16138), .B(n16139), .Z(n16137) );
  XOR U16328 ( .A(n15839), .B(n16140), .Z(n16134) );
  XNOR U16329 ( .A(n16141), .B(n16142), .Z(n16140) );
  AND U16330 ( .A(n15792), .B(n16085), .Z(n16141) );
  XNOR U16331 ( .A(n16126), .B(n16113), .Z(n16121) );
  XOR U16332 ( .A(n16143), .B(n16144), .Z(n16126) );
  XNOR U16333 ( .A(n16145), .B(n16139), .Z(n16144) );
  XOR U16334 ( .A(n16146), .B(n16147), .Z(n16139) );
  XNOR U16335 ( .A(n16148), .B(n16149), .Z(n16147) );
  NAND U16336 ( .A(n16095), .B(n15850), .Z(n16149) );
  XNOR U16337 ( .A(n16150), .B(n16151), .Z(n16143) );
  ANDN U16338 ( .B(n16091), .A(n15844), .Z(n16150) );
  ANDN U16339 ( .B(n16110), .A(n16113), .Z(n16133) );
  XOR U16340 ( .A(n16113), .B(n16110), .Z(n16125) );
  XNOR U16341 ( .A(n16152), .B(n16153), .Z(n16110) );
  XNOR U16342 ( .A(n16146), .B(n16154), .Z(n16153) );
  XNOR U16343 ( .A(n15792), .B(n16145), .Z(n16154) );
  XNOR U16344 ( .A(n16085), .B(n16155), .Z(n16152) );
  XNOR U16345 ( .A(n16156), .B(n16142), .Z(n16155) );
  OR U16346 ( .A(n15838), .B(n16086), .Z(n16142) );
  XNOR U16347 ( .A(n16085), .B(n16138), .Z(n16086) );
  XNOR U16348 ( .A(n15792), .B(n15839), .Z(n15838) );
  ANDN U16349 ( .B(n15839), .A(n15873), .Z(n16156) );
  IV U16350 ( .A(n16138), .Z(n15873) );
  XOR U16351 ( .A(n16157), .B(n16158), .Z(n16113) );
  XOR U16352 ( .A(n16146), .B(n16136), .Z(n16158) );
  XOR U16353 ( .A(n16159), .B(n15811), .Z(n16136) );
  XOR U16354 ( .A(n16160), .B(n16148), .Z(n16146) );
  OR U16355 ( .A(n16098), .B(n16106), .Z(n16148) );
  XOR U16356 ( .A(n16114), .B(n15850), .Z(n16106) );
  XOR U16357 ( .A(n16159), .B(n15839), .Z(n15850) );
  XOR U16358 ( .A(n16161), .B(n16162), .Z(n15839) );
  XNOR U16359 ( .A(n15844), .B(n16163), .Z(n16162) );
  XNOR U16360 ( .A(n16099), .B(n16095), .Z(n16098) );
  XNOR U16361 ( .A(n15811), .B(n16138), .Z(n16095) );
  XOR U16362 ( .A(n16164), .B(n16165), .Z(n16138) );
  XNOR U16363 ( .A(n16166), .B(n16167), .Z(n16165) );
  XOR U16364 ( .A(n16168), .B(n16085), .Z(n16164) );
  ANDN U16365 ( .B(n16099), .A(n16114), .Z(n16160) );
  XNOR U16366 ( .A(n16169), .B(n15792), .Z(n16114) );
  XOR U16367 ( .A(n16166), .B(n16170), .Z(n15792) );
  XOR U16368 ( .A(n16171), .B(n16172), .Z(n16170) );
  XOR U16369 ( .A(n16173), .B(n16174), .Z(n16166) );
  XNOR U16370 ( .A(n16175), .B(n16176), .Z(n16173) );
  XNOR U16371 ( .A(key[612]), .B(n15170), .Z(n16176) );
  XOR U16372 ( .A(n15183), .B(n16177), .Z(n15170) );
  XOR U16373 ( .A(n16085), .B(n16091), .Z(n16099) );
  XOR U16374 ( .A(n16145), .B(n16178), .Z(n16157) );
  XNOR U16375 ( .A(n16179), .B(n16151), .Z(n16178) );
  NANDN U16376 ( .A(n16090), .B(n16103), .Z(n16151) );
  XOR U16377 ( .A(n15844), .B(n16104), .Z(n16103) );
  XNOR U16378 ( .A(n16091), .B(n16180), .Z(n16090) );
  ANDN U16379 ( .B(n16159), .A(n15811), .Z(n16179) );
  IV U16380 ( .A(n16180), .Z(n15811) );
  IV U16381 ( .A(n16104), .Z(n16159) );
  XNOR U16382 ( .A(n16163), .B(n16180), .Z(n16104) );
  XNOR U16383 ( .A(n16181), .B(n16172), .Z(n16180) );
  XNOR U16384 ( .A(n16169), .B(n16091), .Z(n16145) );
  XNOR U16385 ( .A(n16167), .B(n16182), .Z(n16091) );
  XNOR U16386 ( .A(n16172), .B(n16161), .Z(n16182) );
  XOR U16387 ( .A(n16183), .B(n16184), .Z(n16161) );
  XOR U16388 ( .A(n16185), .B(n16186), .Z(n16184) );
  XOR U16389 ( .A(key[610]), .B(n15148), .Z(n16183) );
  XOR U16390 ( .A(n16187), .B(n16188), .Z(n16167) );
  XNOR U16391 ( .A(n16189), .B(n16190), .Z(n16188) );
  XNOR U16392 ( .A(n16191), .B(n16163), .Z(n16190) );
  XOR U16393 ( .A(n16192), .B(n16193), .Z(n16163) );
  XNOR U16394 ( .A(n16194), .B(n16195), .Z(n16193) );
  XOR U16395 ( .A(key[609]), .B(n16196), .Z(n16192) );
  XOR U16396 ( .A(n16197), .B(n16198), .Z(n16187) );
  XNOR U16397 ( .A(key[611]), .B(n15156), .Z(n16198) );
  XOR U16398 ( .A(n15183), .B(n16199), .Z(n15156) );
  IV U16399 ( .A(n15844), .Z(n16169) );
  XNOR U16400 ( .A(n16181), .B(n16168), .Z(n16200) );
  XOR U16401 ( .A(n16201), .B(n16202), .Z(n16168) );
  XNOR U16402 ( .A(n16203), .B(n16204), .Z(n16202) );
  XNOR U16403 ( .A(key[615]), .B(n15183), .Z(n16201) );
  IV U16404 ( .A(n16171), .Z(n16181) );
  XNOR U16405 ( .A(n16205), .B(n16206), .Z(n16171) );
  XNOR U16406 ( .A(n16207), .B(n16208), .Z(n16206) );
  XOR U16407 ( .A(key[613]), .B(n16209), .Z(n16205) );
  XOR U16408 ( .A(n16210), .B(n16211), .Z(n16172) );
  XNOR U16409 ( .A(n16085), .B(n16212), .Z(n16211) );
  XOR U16410 ( .A(n16213), .B(n16214), .Z(n16085) );
  XNOR U16411 ( .A(n16215), .B(n16216), .Z(n16214) );
  XOR U16412 ( .A(key[608]), .B(n15181), .Z(n16213) );
  XOR U16413 ( .A(n16217), .B(n16218), .Z(n16210) );
  XNOR U16414 ( .A(key[614]), .B(n15175), .Z(n16218) );
  XOR U16415 ( .A(n15183), .B(n16219), .Z(n15175) );
  XOR U16416 ( .A(n16220), .B(n16221), .Z(n13095) );
  XNOR U16417 ( .A(n16222), .B(n15831), .Z(n16221) );
  XNOR U16418 ( .A(n16223), .B(n16224), .Z(n15831) );
  XNOR U16419 ( .A(n16225), .B(n16226), .Z(n16224) );
  OR U16420 ( .A(n15885), .B(n16227), .Z(n16226) );
  XNOR U16421 ( .A(n15814), .B(n16228), .Z(n16220) );
  XOR U16422 ( .A(n16229), .B(n16230), .Z(n16228) );
  ANDN U16423 ( .B(n16231), .A(n15879), .Z(n16230) );
  XNOR U16424 ( .A(n16223), .B(n16232), .Z(n15814) );
  XNOR U16425 ( .A(n15877), .B(n16233), .Z(n16232) );
  OR U16426 ( .A(n16234), .B(n16235), .Z(n16233) );
  OR U16427 ( .A(n16236), .B(n16237), .Z(n15877) );
  XNOR U16428 ( .A(n15875), .B(n16238), .Z(n16223) );
  XNOR U16429 ( .A(n16239), .B(n16240), .Z(n16238) );
  NAND U16430 ( .A(n16241), .B(n16242), .Z(n16240) );
  XNOR U16431 ( .A(key[725]), .B(n13087), .Z(n15924) );
  XNOR U16432 ( .A(n12458), .B(n14140), .Z(n13087) );
  XNOR U16433 ( .A(n15758), .B(n15832), .Z(n14140) );
  XNOR U16434 ( .A(n15815), .B(n15759), .Z(n15832) );
  XNOR U16435 ( .A(n16222), .B(n16243), .Z(n15759) );
  XNOR U16436 ( .A(n15883), .B(n16244), .Z(n16243) );
  NANDN U16437 ( .A(n16245), .B(n16246), .Z(n16244) );
  OR U16438 ( .A(n16247), .B(n16248), .Z(n15883) );
  XNOR U16439 ( .A(n15875), .B(n16249), .Z(n15815) );
  XOR U16440 ( .A(n16250), .B(n16225), .Z(n16249) );
  OR U16441 ( .A(n16248), .B(n16251), .Z(n16225) );
  XNOR U16442 ( .A(n15885), .B(n16245), .Z(n16248) );
  NOR U16443 ( .A(n16252), .B(n16245), .Z(n16250) );
  XOR U16444 ( .A(n16253), .B(n16239), .Z(n15875) );
  OR U16445 ( .A(n16254), .B(n16255), .Z(n16239) );
  ANDN U16446 ( .B(n16256), .A(n16257), .Z(n16253) );
  XNOR U16447 ( .A(n15886), .B(n16258), .Z(n15758) );
  XNOR U16448 ( .A(n16259), .B(n16229), .Z(n16258) );
  NOR U16449 ( .A(n16237), .B(n16260), .Z(n16229) );
  XOR U16450 ( .A(n16234), .B(n16261), .Z(n16237) );
  NOR U16451 ( .A(n16262), .B(n16234), .Z(n16259) );
  XNOR U16452 ( .A(n16222), .B(n16263), .Z(n15886) );
  XNOR U16453 ( .A(n16264), .B(n16265), .Z(n16263) );
  NAND U16454 ( .A(n16266), .B(n16241), .Z(n16265) );
  XOR U16455 ( .A(n16267), .B(n16264), .Z(n16222) );
  NANDN U16456 ( .A(n16254), .B(n16268), .Z(n16264) );
  XOR U16457 ( .A(n16269), .B(n16241), .Z(n16254) );
  XOR U16458 ( .A(n16245), .B(n15879), .Z(n16241) );
  IV U16459 ( .A(n16261), .Z(n15879) );
  XOR U16460 ( .A(n16270), .B(n16271), .Z(n16261) );
  NANDN U16461 ( .A(n16272), .B(n16273), .Z(n16271) );
  XNOR U16462 ( .A(n16274), .B(n16275), .Z(n16245) );
  OR U16463 ( .A(n16272), .B(n16276), .Z(n16275) );
  ANDN U16464 ( .B(n16277), .A(n16269), .Z(n16267) );
  IV U16465 ( .A(n16256), .Z(n16269) );
  XOR U16466 ( .A(n15885), .B(n16234), .Z(n16256) );
  XNOR U16467 ( .A(n16270), .B(n16278), .Z(n16234) );
  NANDN U16468 ( .A(n16279), .B(n16280), .Z(n16278) );
  NANDN U16469 ( .A(n16281), .B(n16282), .Z(n16270) );
  OR U16470 ( .A(n16284), .B(n16281), .Z(n16274) );
  XOR U16471 ( .A(n16285), .B(n16272), .Z(n16281) );
  XNOR U16472 ( .A(n16286), .B(n16287), .Z(n16272) );
  XOR U16473 ( .A(n16288), .B(n16280), .Z(n16287) );
  XNOR U16474 ( .A(n16289), .B(n16290), .Z(n16286) );
  XNOR U16475 ( .A(n16291), .B(n16292), .Z(n16290) );
  ANDN U16476 ( .B(n16280), .A(n16293), .Z(n16291) );
  IV U16477 ( .A(n16294), .Z(n16280) );
  ANDN U16478 ( .B(n16285), .A(n16293), .Z(n16283) );
  IV U16479 ( .A(n16279), .Z(n16285) );
  XNOR U16480 ( .A(n16288), .B(n16295), .Z(n16279) );
  XNOR U16481 ( .A(n16292), .B(n16296), .Z(n16295) );
  NANDN U16482 ( .A(n16276), .B(n16273), .Z(n16296) );
  NANDN U16483 ( .A(n16284), .B(n16282), .Z(n16292) );
  XNOR U16484 ( .A(n16273), .B(n16294), .Z(n16282) );
  XOR U16485 ( .A(n16297), .B(n16298), .Z(n16294) );
  XOR U16486 ( .A(n16299), .B(n16300), .Z(n16298) );
  XNOR U16487 ( .A(n16246), .B(n16301), .Z(n16300) );
  XNOR U16488 ( .A(n16302), .B(n16303), .Z(n16297) );
  XNOR U16489 ( .A(n16304), .B(n16305), .Z(n16303) );
  ANDN U16490 ( .B(n16306), .A(n16227), .Z(n16304) );
  XNOR U16491 ( .A(n16293), .B(n16276), .Z(n16284) );
  IV U16492 ( .A(n16289), .Z(n16293) );
  XOR U16493 ( .A(n16307), .B(n16308), .Z(n16289) );
  XNOR U16494 ( .A(n16309), .B(n16301), .Z(n16308) );
  XOR U16495 ( .A(n16310), .B(n16311), .Z(n16301) );
  XNOR U16496 ( .A(n16312), .B(n16313), .Z(n16311) );
  NAND U16497 ( .A(n16242), .B(n16266), .Z(n16313) );
  XNOR U16498 ( .A(n16314), .B(n16315), .Z(n16307) );
  ANDN U16499 ( .B(n16316), .A(n16235), .Z(n16314) );
  XOR U16500 ( .A(n16276), .B(n16273), .Z(n16288) );
  XNOR U16501 ( .A(n16317), .B(n16318), .Z(n16273) );
  XNOR U16502 ( .A(n16310), .B(n16319), .Z(n16318) );
  XOR U16503 ( .A(n16309), .B(n15884), .Z(n16319) );
  XOR U16504 ( .A(n16227), .B(n16320), .Z(n16317) );
  XNOR U16505 ( .A(n16321), .B(n16305), .Z(n16320) );
  OR U16506 ( .A(n16247), .B(n16251), .Z(n16305) );
  XNOR U16507 ( .A(n16227), .B(n16252), .Z(n16251) );
  XOR U16508 ( .A(n15884), .B(n16246), .Z(n16247) );
  ANDN U16509 ( .B(n16246), .A(n16252), .Z(n16321) );
  XOR U16510 ( .A(n16322), .B(n16323), .Z(n16276) );
  XOR U16511 ( .A(n16310), .B(n16299), .Z(n16323) );
  XNOR U16512 ( .A(n15880), .B(n16231), .Z(n16299) );
  XOR U16513 ( .A(n16324), .B(n16312), .Z(n16310) );
  NANDN U16514 ( .A(n16255), .B(n16268), .Z(n16312) );
  XOR U16515 ( .A(n16277), .B(n16266), .Z(n16268) );
  XOR U16516 ( .A(n16231), .B(n16246), .Z(n16266) );
  XNOR U16517 ( .A(n16316), .B(n16325), .Z(n16246) );
  XOR U16518 ( .A(n16326), .B(n16327), .Z(n16325) );
  XOR U16519 ( .A(n16257), .B(n16242), .Z(n16255) );
  XNOR U16520 ( .A(n16252), .B(n15880), .Z(n16242) );
  IV U16521 ( .A(n16302), .Z(n16252) );
  XOR U16522 ( .A(n16328), .B(n16329), .Z(n16302) );
  XOR U16523 ( .A(n16330), .B(n16331), .Z(n16329) );
  XNOR U16524 ( .A(n16227), .B(n16332), .Z(n16328) );
  ANDN U16525 ( .B(n16277), .A(n16257), .Z(n16324) );
  XNOR U16526 ( .A(n16227), .B(n16235), .Z(n16257) );
  XOR U16527 ( .A(n16309), .B(n16333), .Z(n16322) );
  XNOR U16528 ( .A(n16334), .B(n16315), .Z(n16333) );
  OR U16529 ( .A(n16260), .B(n16236), .Z(n16315) );
  XNOR U16530 ( .A(n16335), .B(n15880), .Z(n16236) );
  XNOR U16531 ( .A(n16316), .B(n16231), .Z(n16260) );
  AND U16532 ( .A(n16231), .B(n15880), .Z(n16334) );
  XOR U16533 ( .A(n16336), .B(n16337), .Z(n15880) );
  XNOR U16534 ( .A(n16337), .B(n16338), .Z(n16231) );
  XNOR U16535 ( .A(n16339), .B(n16336), .Z(n16338) );
  XNOR U16536 ( .A(n16235), .B(n16262), .Z(n16309) );
  IV U16537 ( .A(n16335), .Z(n16235) );
  XNOR U16538 ( .A(n16326), .B(n16332), .Z(n16340) );
  XOR U16539 ( .A(n16341), .B(n16342), .Z(n16332) );
  XNOR U16540 ( .A(n16343), .B(n16344), .Z(n16342) );
  XNOR U16541 ( .A(n16345), .B(n16327), .Z(n16344) );
  IV U16542 ( .A(n16339), .Z(n16327) );
  XOR U16543 ( .A(n16346), .B(n16347), .Z(n16339) );
  XNOR U16544 ( .A(n15619), .B(n16348), .Z(n16347) );
  XNOR U16545 ( .A(n15584), .B(n16349), .Z(n16346) );
  XOR U16546 ( .A(key[521]), .B(n16350), .Z(n16349) );
  XNOR U16547 ( .A(n15622), .B(n16351), .Z(n16341) );
  XOR U16548 ( .A(key[523]), .B(n15624), .Z(n16351) );
  XOR U16549 ( .A(n16352), .B(n15611), .Z(n15622) );
  XOR U16550 ( .A(n16353), .B(n16354), .Z(n16326) );
  XNOR U16551 ( .A(n16355), .B(n15582), .Z(n16354) );
  XOR U16552 ( .A(n16356), .B(n16357), .Z(n16353) );
  XNOR U16553 ( .A(key[522]), .B(n16358), .Z(n16357) );
  XOR U16554 ( .A(n16316), .B(n16306), .Z(n16277) );
  IV U16555 ( .A(n15884), .Z(n16306) );
  XOR U16556 ( .A(n16337), .B(n16359), .Z(n15884) );
  XOR U16557 ( .A(n16336), .B(n16331), .Z(n16359) );
  XNOR U16558 ( .A(n16360), .B(n16361), .Z(n16331) );
  XOR U16559 ( .A(n15609), .B(n16362), .Z(n16361) );
  XOR U16560 ( .A(n16363), .B(n16364), .Z(n15609) );
  XNOR U16561 ( .A(n16365), .B(n16366), .Z(n16364) );
  XNOR U16562 ( .A(n16367), .B(n15599), .Z(n16363) );
  XNOR U16563 ( .A(key[524]), .B(n16368), .Z(n16360) );
  IV U16564 ( .A(n16262), .Z(n16316) );
  XOR U16565 ( .A(n16337), .B(n16369), .Z(n16262) );
  XNOR U16566 ( .A(n16336), .B(n16330), .Z(n16369) );
  XOR U16567 ( .A(n16370), .B(n16371), .Z(n16330) );
  XOR U16568 ( .A(n16372), .B(n15605), .Z(n16371) );
  XOR U16569 ( .A(n16373), .B(n16374), .Z(n15605) );
  XOR U16570 ( .A(key[527]), .B(n15629), .Z(n16370) );
  XOR U16571 ( .A(n16375), .B(n16376), .Z(n16336) );
  XOR U16572 ( .A(n16227), .B(n16377), .Z(n16376) );
  XNOR U16573 ( .A(n16378), .B(n16379), .Z(n16227) );
  XNOR U16574 ( .A(n16380), .B(n16381), .Z(n16379) );
  XNOR U16575 ( .A(n16382), .B(n16383), .Z(n16378) );
  XNOR U16576 ( .A(key[520]), .B(n16384), .Z(n16383) );
  XNOR U16577 ( .A(n16385), .B(n16386), .Z(n16375) );
  XNOR U16578 ( .A(key[526]), .B(n15591), .Z(n16386) );
  XNOR U16579 ( .A(n15604), .B(n16387), .Z(n15591) );
  XOR U16580 ( .A(n16352), .B(n16388), .Z(n15604) );
  XNOR U16581 ( .A(n16389), .B(n16390), .Z(n16337) );
  XOR U16582 ( .A(n16391), .B(n15597), .Z(n16390) );
  XNOR U16583 ( .A(n16392), .B(n16393), .Z(n15597) );
  XNOR U16584 ( .A(n16394), .B(n16395), .Z(n16389) );
  XOR U16585 ( .A(key[525]), .B(n15593), .Z(n16395) );
  XOR U16586 ( .A(n15888), .B(n15731), .Z(n12458) );
  XNOR U16587 ( .A(n15907), .B(n16396), .Z(n15731) );
  XOR U16588 ( .A(n16397), .B(n15822), .Z(n16396) );
  NANDN U16589 ( .A(n16398), .B(n15916), .Z(n15822) );
  XNOR U16590 ( .A(n15918), .B(n15824), .Z(n15916) );
  NOR U16591 ( .A(n16399), .B(n15918), .Z(n16397) );
  XOR U16592 ( .A(n15819), .B(n16400), .Z(n15907) );
  XNOR U16593 ( .A(n16401), .B(n16402), .Z(n16400) );
  NAND U16594 ( .A(n16403), .B(n15922), .Z(n16402) );
  XOR U16595 ( .A(n15752), .B(n15733), .Z(n15888) );
  XNOR U16596 ( .A(n15819), .B(n16404), .Z(n15733) );
  XNOR U16597 ( .A(n15909), .B(n16405), .Z(n16404) );
  NANDN U16598 ( .A(n16406), .B(n16407), .Z(n16405) );
  OR U16599 ( .A(n16408), .B(n16409), .Z(n15909) );
  XOR U16600 ( .A(n16410), .B(n16401), .Z(n15819) );
  NANDN U16601 ( .A(n16411), .B(n16412), .Z(n16401) );
  ANDN U16602 ( .B(n16413), .A(n16414), .Z(n16410) );
  IV U16603 ( .A(n15912), .Z(n15752) );
  XNOR U16604 ( .A(n15902), .B(n16415), .Z(n15912) );
  XOR U16605 ( .A(n16416), .B(n15898), .Z(n16415) );
  OR U16606 ( .A(n16408), .B(n16417), .Z(n15898) );
  XNOR U16607 ( .A(n15901), .B(n16407), .Z(n16408) );
  ANDN U16608 ( .B(n16407), .A(n16418), .Z(n16416) );
  XOR U16609 ( .A(n16419), .B(n15920), .Z(n15902) );
  OR U16610 ( .A(n16411), .B(n16420), .Z(n15920) );
  XNOR U16611 ( .A(n16421), .B(n15922), .Z(n16411) );
  XOR U16612 ( .A(n16407), .B(n15824), .Z(n15922) );
  XOR U16613 ( .A(n16422), .B(n16423), .Z(n15824) );
  NANDN U16614 ( .A(n16424), .B(n16425), .Z(n16423) );
  XOR U16615 ( .A(n16426), .B(n16427), .Z(n16407) );
  NANDN U16616 ( .A(n16424), .B(n16428), .Z(n16427) );
  ANDN U16617 ( .B(n16421), .A(n16429), .Z(n16419) );
  IV U16618 ( .A(n16414), .Z(n16421) );
  XOR U16619 ( .A(n15918), .B(n15901), .Z(n16414) );
  XNOR U16620 ( .A(n16430), .B(n16426), .Z(n15901) );
  NANDN U16621 ( .A(n16431), .B(n16432), .Z(n16426) );
  XOR U16622 ( .A(n16428), .B(n16433), .Z(n16432) );
  ANDN U16623 ( .B(n16433), .A(n16434), .Z(n16430) );
  XOR U16624 ( .A(n16435), .B(n16422), .Z(n15918) );
  NANDN U16625 ( .A(n16431), .B(n16436), .Z(n16422) );
  XOR U16626 ( .A(n16437), .B(n16425), .Z(n16436) );
  XNOR U16627 ( .A(n16438), .B(n16439), .Z(n16424) );
  XOR U16628 ( .A(n16440), .B(n16441), .Z(n16439) );
  XNOR U16629 ( .A(n16442), .B(n16443), .Z(n16438) );
  XNOR U16630 ( .A(n16444), .B(n16445), .Z(n16443) );
  ANDN U16631 ( .B(n16437), .A(n16441), .Z(n16444) );
  ANDN U16632 ( .B(n16437), .A(n16434), .Z(n16435) );
  XNOR U16633 ( .A(n16440), .B(n16446), .Z(n16434) );
  XOR U16634 ( .A(n16447), .B(n16445), .Z(n16446) );
  NAND U16635 ( .A(n16448), .B(n16449), .Z(n16445) );
  XNOR U16636 ( .A(n16442), .B(n16425), .Z(n16449) );
  IV U16637 ( .A(n16437), .Z(n16442) );
  XNOR U16638 ( .A(n16428), .B(n16441), .Z(n16448) );
  IV U16639 ( .A(n16433), .Z(n16441) );
  XOR U16640 ( .A(n16450), .B(n16451), .Z(n16433) );
  XNOR U16641 ( .A(n16452), .B(n16453), .Z(n16451) );
  XNOR U16642 ( .A(n16454), .B(n16455), .Z(n16450) );
  ANDN U16643 ( .B(n15917), .A(n16399), .Z(n16454) );
  AND U16644 ( .A(n16425), .B(n16428), .Z(n16447) );
  XNOR U16645 ( .A(n16425), .B(n16428), .Z(n16440) );
  XNOR U16646 ( .A(n16456), .B(n16457), .Z(n16428) );
  XNOR U16647 ( .A(n16458), .B(n16453), .Z(n16457) );
  XOR U16648 ( .A(n16459), .B(n16460), .Z(n16456) );
  XNOR U16649 ( .A(n16461), .B(n16455), .Z(n16460) );
  OR U16650 ( .A(n16398), .B(n15915), .Z(n16455) );
  XNOR U16651 ( .A(n15917), .B(n16462), .Z(n15915) );
  XNOR U16652 ( .A(n16399), .B(n15825), .Z(n16398) );
  ANDN U16653 ( .B(n16463), .A(n15906), .Z(n16461) );
  XNOR U16654 ( .A(n16464), .B(n16465), .Z(n16425) );
  XNOR U16655 ( .A(n16453), .B(n16466), .Z(n16465) );
  XOR U16656 ( .A(n15911), .B(n16459), .Z(n16466) );
  XNOR U16657 ( .A(n15917), .B(n16399), .Z(n16453) );
  XOR U16658 ( .A(n15900), .B(n16467), .Z(n16464) );
  XNOR U16659 ( .A(n16468), .B(n16469), .Z(n16467) );
  ANDN U16660 ( .B(n16470), .A(n16418), .Z(n16468) );
  XNOR U16661 ( .A(n16471), .B(n16472), .Z(n16437) );
  XNOR U16662 ( .A(n16458), .B(n16473), .Z(n16472) );
  XNOR U16663 ( .A(n16406), .B(n16452), .Z(n16473) );
  XOR U16664 ( .A(n16459), .B(n16474), .Z(n16452) );
  XNOR U16665 ( .A(n16475), .B(n16476), .Z(n16474) );
  NAND U16666 ( .A(n15923), .B(n16403), .Z(n16476) );
  XNOR U16667 ( .A(n16477), .B(n16475), .Z(n16459) );
  NANDN U16668 ( .A(n16420), .B(n16412), .Z(n16475) );
  XOR U16669 ( .A(n16413), .B(n16403), .Z(n16412) );
  XNOR U16670 ( .A(n16470), .B(n15825), .Z(n16403) );
  XOR U16671 ( .A(n16429), .B(n15923), .Z(n16420) );
  XNOR U16672 ( .A(n16418), .B(n16462), .Z(n15923) );
  ANDN U16673 ( .B(n16413), .A(n16429), .Z(n16477) );
  XOR U16674 ( .A(n15900), .B(n15917), .Z(n16429) );
  XNOR U16675 ( .A(n16478), .B(n16479), .Z(n15917) );
  XNOR U16676 ( .A(n16480), .B(n16481), .Z(n16479) );
  XOR U16677 ( .A(n16462), .B(n16463), .Z(n16458) );
  IV U16678 ( .A(n15825), .Z(n16463) );
  XOR U16679 ( .A(n16482), .B(n16483), .Z(n15825) );
  XOR U16680 ( .A(n16484), .B(n16481), .Z(n16483) );
  IV U16681 ( .A(n15906), .Z(n16462) );
  XOR U16682 ( .A(n16481), .B(n16485), .Z(n15906) );
  XNOR U16683 ( .A(n16486), .B(n16487), .Z(n16471) );
  XNOR U16684 ( .A(n16488), .B(n16469), .Z(n16487) );
  OR U16685 ( .A(n16409), .B(n16417), .Z(n16469) );
  XNOR U16686 ( .A(n15900), .B(n16418), .Z(n16417) );
  IV U16687 ( .A(n16486), .Z(n16418) );
  XOR U16688 ( .A(n15911), .B(n16470), .Z(n16409) );
  IV U16689 ( .A(n16406), .Z(n16470) );
  XNOR U16690 ( .A(n16490), .B(n16478), .Z(n16489) );
  XOR U16691 ( .A(n16491), .B(n16492), .Z(n16478) );
  XNOR U16692 ( .A(n16493), .B(n16494), .Z(n16492) );
  XNOR U16693 ( .A(key[562]), .B(n16495), .Z(n16491) );
  IV U16694 ( .A(n16484), .Z(n16490) );
  XOR U16695 ( .A(n16482), .B(n16496), .Z(n16399) );
  XOR U16696 ( .A(n16481), .B(n16497), .Z(n16496) );
  NOR U16697 ( .A(n15911), .B(n15900), .Z(n16488) );
  XOR U16698 ( .A(n16482), .B(n16498), .Z(n15911) );
  XOR U16699 ( .A(n16481), .B(n16499), .Z(n16498) );
  XOR U16700 ( .A(n16500), .B(n16501), .Z(n16481) );
  XNOR U16701 ( .A(n15900), .B(n16502), .Z(n16501) );
  XNOR U16702 ( .A(n16503), .B(n16504), .Z(n16500) );
  XNOR U16703 ( .A(key[566]), .B(n15473), .Z(n16504) );
  XOR U16704 ( .A(n16505), .B(n16506), .Z(n15473) );
  IV U16705 ( .A(n16485), .Z(n16482) );
  XOR U16706 ( .A(n16507), .B(n16508), .Z(n16485) );
  XOR U16707 ( .A(n16509), .B(n16510), .Z(n16508) );
  XNOR U16708 ( .A(key[565]), .B(n16511), .Z(n16507) );
  XOR U16709 ( .A(n16512), .B(n16513), .Z(n16486) );
  XNOR U16710 ( .A(n16499), .B(n16497), .Z(n16513) );
  XNOR U16711 ( .A(n16514), .B(n16515), .Z(n16497) );
  XNOR U16712 ( .A(n16516), .B(n16517), .Z(n16515) );
  XNOR U16713 ( .A(key[567]), .B(n15495), .Z(n16514) );
  XNOR U16714 ( .A(n16518), .B(n16519), .Z(n16499) );
  XOR U16715 ( .A(n16520), .B(n16521), .Z(n16518) );
  XNOR U16716 ( .A(key[564]), .B(n15443), .Z(n16521) );
  XNOR U16717 ( .A(n16522), .B(n16505), .Z(n15443) );
  XNOR U16718 ( .A(n15900), .B(n16480), .Z(n16512) );
  XOR U16719 ( .A(n16523), .B(n16524), .Z(n16480) );
  XNOR U16720 ( .A(n16525), .B(n16526), .Z(n16524) );
  XOR U16721 ( .A(n16527), .B(n16484), .Z(n16526) );
  XNOR U16722 ( .A(n16528), .B(n16529), .Z(n16484) );
  XNOR U16723 ( .A(n15464), .B(n16530), .Z(n16529) );
  XNOR U16724 ( .A(key[561]), .B(n16531), .Z(n16528) );
  XNOR U16725 ( .A(n15479), .B(n16532), .Z(n16523) );
  XOR U16726 ( .A(key[563]), .B(n16533), .Z(n16532) );
  XNOR U16727 ( .A(n15495), .B(n16534), .Z(n15479) );
  XNOR U16728 ( .A(n16535), .B(n16536), .Z(n15900) );
  XOR U16729 ( .A(n15493), .B(n16537), .Z(n16536) );
  XNOR U16730 ( .A(key[560]), .B(n16538), .Z(n16535) );
  XNOR U16731 ( .A(n9605), .B(n16539), .Z(n14653) );
  XNOR U16732 ( .A(key[870]), .B(n10493), .Z(n16539) );
  XNOR U16733 ( .A(n14657), .B(n14652), .Z(n10493) );
  XNOR U16734 ( .A(n14691), .B(n16540), .Z(n14652) );
  XNOR U16735 ( .A(n16541), .B(n14585), .Z(n16540) );
  ANDN U16736 ( .B(n14704), .A(n16542), .Z(n14585) );
  XOR U16737 ( .A(n14705), .B(n14587), .Z(n14704) );
  ANDN U16738 ( .B(n14705), .A(n16543), .Z(n16541) );
  XNOR U16739 ( .A(n14581), .B(n16544), .Z(n14691) );
  XNOR U16740 ( .A(n16545), .B(n16546), .Z(n16544) );
  NANDN U16741 ( .A(n14710), .B(n16547), .Z(n16546) );
  XNOR U16742 ( .A(n14635), .B(n14651), .Z(n14657) );
  XOR U16743 ( .A(n14581), .B(n16548), .Z(n14651) );
  XNOR U16744 ( .A(n14693), .B(n16549), .Z(n16548) );
  NANDN U16745 ( .A(n16550), .B(n16551), .Z(n16549) );
  OR U16746 ( .A(n16552), .B(n16553), .Z(n14693) );
  XOR U16747 ( .A(n16554), .B(n16545), .Z(n14581) );
  NANDN U16748 ( .A(n16555), .B(n16556), .Z(n16545) );
  ANDN U16749 ( .B(n16557), .A(n16558), .Z(n16554) );
  XOR U16750 ( .A(n14696), .B(n16559), .Z(n14635) );
  XOR U16751 ( .A(n16560), .B(n14687), .Z(n16559) );
  OR U16752 ( .A(n16561), .B(n16552), .Z(n14687) );
  XNOR U16753 ( .A(n14689), .B(n16550), .Z(n16552) );
  NOR U16754 ( .A(n16562), .B(n16550), .Z(n16560) );
  XOR U16755 ( .A(n16563), .B(n14708), .Z(n14696) );
  OR U16756 ( .A(n16555), .B(n16564), .Z(n14708) );
  XOR U16757 ( .A(n16565), .B(n14710), .Z(n16555) );
  XOR U16758 ( .A(n16550), .B(n14587), .Z(n14710) );
  XOR U16759 ( .A(n16566), .B(n16567), .Z(n14587) );
  NANDN U16760 ( .A(n16568), .B(n16569), .Z(n16567) );
  XNOR U16761 ( .A(n16570), .B(n16571), .Z(n16550) );
  OR U16762 ( .A(n16568), .B(n16572), .Z(n16571) );
  ANDN U16763 ( .B(n16565), .A(n16573), .Z(n16563) );
  IV U16764 ( .A(n16558), .Z(n16565) );
  XOR U16765 ( .A(n14689), .B(n14705), .Z(n16558) );
  XNOR U16766 ( .A(n16574), .B(n16566), .Z(n14705) );
  NANDN U16767 ( .A(n16575), .B(n16576), .Z(n16566) );
  ANDN U16768 ( .B(n16577), .A(n16578), .Z(n16574) );
  NANDN U16769 ( .A(n16575), .B(n16580), .Z(n16570) );
  XOR U16770 ( .A(n16581), .B(n16568), .Z(n16575) );
  XNOR U16771 ( .A(n16582), .B(n16583), .Z(n16568) );
  XOR U16772 ( .A(n16584), .B(n16577), .Z(n16583) );
  XNOR U16773 ( .A(n16585), .B(n16586), .Z(n16582) );
  XNOR U16774 ( .A(n16587), .B(n16588), .Z(n16586) );
  ANDN U16775 ( .B(n16577), .A(n16589), .Z(n16587) );
  IV U16776 ( .A(n16590), .Z(n16577) );
  ANDN U16777 ( .B(n16581), .A(n16589), .Z(n16579) );
  IV U16778 ( .A(n16585), .Z(n16589) );
  IV U16779 ( .A(n16578), .Z(n16581) );
  XNOR U16780 ( .A(n16584), .B(n16591), .Z(n16578) );
  XOR U16781 ( .A(n16592), .B(n16588), .Z(n16591) );
  NAND U16782 ( .A(n16580), .B(n16576), .Z(n16588) );
  XNOR U16783 ( .A(n16569), .B(n16590), .Z(n16576) );
  XOR U16784 ( .A(n16593), .B(n16594), .Z(n16590) );
  XOR U16785 ( .A(n16595), .B(n16596), .Z(n16594) );
  XNOR U16786 ( .A(n16551), .B(n16597), .Z(n16596) );
  XNOR U16787 ( .A(n16598), .B(n16599), .Z(n16593) );
  XNOR U16788 ( .A(n16600), .B(n16601), .Z(n16599) );
  ANDN U16789 ( .B(n16602), .A(n14690), .Z(n16600) );
  XNOR U16790 ( .A(n16585), .B(n16572), .Z(n16580) );
  XOR U16791 ( .A(n16603), .B(n16604), .Z(n16585) );
  XNOR U16792 ( .A(n16605), .B(n16597), .Z(n16604) );
  XOR U16793 ( .A(n16606), .B(n16607), .Z(n16597) );
  XNOR U16794 ( .A(n16608), .B(n16609), .Z(n16607) );
  NAND U16795 ( .A(n14711), .B(n16547), .Z(n16609) );
  XNOR U16796 ( .A(n16610), .B(n16611), .Z(n16603) );
  ANDN U16797 ( .B(n16612), .A(n14706), .Z(n16610) );
  ANDN U16798 ( .B(n16569), .A(n16572), .Z(n16592) );
  XOR U16799 ( .A(n16572), .B(n16569), .Z(n16584) );
  XNOR U16800 ( .A(n16613), .B(n16614), .Z(n16569) );
  XNOR U16801 ( .A(n16606), .B(n16615), .Z(n16614) );
  XOR U16802 ( .A(n16605), .B(n14695), .Z(n16615) );
  XOR U16803 ( .A(n14690), .B(n16616), .Z(n16613) );
  XNOR U16804 ( .A(n16617), .B(n16601), .Z(n16616) );
  OR U16805 ( .A(n16553), .B(n16561), .Z(n16601) );
  XNOR U16806 ( .A(n14690), .B(n16562), .Z(n16561) );
  XOR U16807 ( .A(n14695), .B(n16551), .Z(n16553) );
  ANDN U16808 ( .B(n16551), .A(n16562), .Z(n16617) );
  XOR U16809 ( .A(n16618), .B(n16619), .Z(n16572) );
  XOR U16810 ( .A(n16606), .B(n16595), .Z(n16619) );
  XOR U16811 ( .A(n14700), .B(n14588), .Z(n16595) );
  XOR U16812 ( .A(n16620), .B(n16608), .Z(n16606) );
  NANDN U16813 ( .A(n16564), .B(n16556), .Z(n16608) );
  XOR U16814 ( .A(n16557), .B(n16547), .Z(n16556) );
  XNOR U16815 ( .A(n16612), .B(n16621), .Z(n16551) );
  XOR U16816 ( .A(n16622), .B(n16623), .Z(n16621) );
  XOR U16817 ( .A(n16573), .B(n14711), .Z(n16564) );
  XNOR U16818 ( .A(n16562), .B(n14700), .Z(n14711) );
  IV U16819 ( .A(n16598), .Z(n16562) );
  XOR U16820 ( .A(n16624), .B(n16625), .Z(n16598) );
  XOR U16821 ( .A(n16626), .B(n16627), .Z(n16625) );
  XNOR U16822 ( .A(n14690), .B(n16628), .Z(n16624) );
  ANDN U16823 ( .B(n16557), .A(n16573), .Z(n16620) );
  XNOR U16824 ( .A(n14690), .B(n14706), .Z(n16573) );
  XOR U16825 ( .A(n16612), .B(n16602), .Z(n16557) );
  IV U16826 ( .A(n14695), .Z(n16602) );
  XOR U16827 ( .A(n16629), .B(n16630), .Z(n14695) );
  XOR U16828 ( .A(n16631), .B(n16627), .Z(n16630) );
  XNOR U16829 ( .A(n16632), .B(n16633), .Z(n16627) );
  XOR U16830 ( .A(n12124), .B(n13987), .Z(n16633) );
  XOR U16831 ( .A(n13984), .B(n13537), .Z(n13987) );
  XNOR U16832 ( .A(n13990), .B(n13518), .Z(n12124) );
  XOR U16833 ( .A(n16634), .B(n13563), .Z(n13990) );
  XNOR U16834 ( .A(n12123), .B(n16635), .Z(n16632) );
  XNOR U16835 ( .A(key[764]), .B(n13564), .Z(n16635) );
  IV U16836 ( .A(n13988), .Z(n13564) );
  XOR U16837 ( .A(n16636), .B(n13561), .Z(n13988) );
  XNOR U16838 ( .A(n14002), .B(n13975), .Z(n12123) );
  IV U16839 ( .A(n12141), .Z(n13975) );
  XOR U16840 ( .A(n16637), .B(n16638), .Z(n12141) );
  XNOR U16841 ( .A(n16639), .B(n16640), .Z(n16638) );
  XNOR U16842 ( .A(n16641), .B(n16642), .Z(n16637) );
  XOR U16843 ( .A(n16643), .B(n16644), .Z(n16642) );
  ANDN U16844 ( .B(n16645), .A(n16646), .Z(n16644) );
  IV U16845 ( .A(n16543), .Z(n16612) );
  XOR U16846 ( .A(n16605), .B(n16647), .Z(n16618) );
  XNOR U16847 ( .A(n16648), .B(n16611), .Z(n16647) );
  OR U16848 ( .A(n16542), .B(n14703), .Z(n16611) );
  XNOR U16849 ( .A(n16649), .B(n14700), .Z(n14703) );
  XNOR U16850 ( .A(n16543), .B(n14588), .Z(n16542) );
  ANDN U16851 ( .B(n14700), .A(n14588), .Z(n16648) );
  XOR U16852 ( .A(n16629), .B(n16650), .Z(n14588) );
  XNOR U16853 ( .A(n16651), .B(n16631), .Z(n16650) );
  XOR U16854 ( .A(n16631), .B(n16629), .Z(n14700) );
  XNOR U16855 ( .A(n14706), .B(n16543), .Z(n16605) );
  XOR U16856 ( .A(n16629), .B(n16652), .Z(n16543) );
  XNOR U16857 ( .A(n16631), .B(n16626), .Z(n16652) );
  XOR U16858 ( .A(n16653), .B(n16654), .Z(n16626) );
  XNOR U16859 ( .A(n13553), .B(n12137), .Z(n16654) );
  XNOR U16860 ( .A(n13983), .B(n13532), .Z(n12137) );
  XNOR U16861 ( .A(n16655), .B(n16656), .Z(n13983) );
  XNOR U16862 ( .A(n16657), .B(n16658), .Z(n16656) );
  XOR U16863 ( .A(n16659), .B(n16660), .Z(n16655) );
  XOR U16864 ( .A(n16661), .B(n16662), .Z(n13553) );
  XNOR U16865 ( .A(n16663), .B(n16664), .Z(n16662) );
  XOR U16866 ( .A(n16665), .B(n16666), .Z(n16661) );
  XOR U16867 ( .A(n13984), .B(n14002), .Z(n12170) );
  XNOR U16868 ( .A(n16667), .B(n16668), .Z(n16629) );
  XNOR U16869 ( .A(n13522), .B(n12142), .Z(n16668) );
  XNOR U16870 ( .A(n16669), .B(n16670), .Z(n13537) );
  XNOR U16871 ( .A(n16671), .B(n16672), .Z(n16670) );
  XNOR U16872 ( .A(n16673), .B(n16674), .Z(n16669) );
  XOR U16873 ( .A(n16675), .B(n16676), .Z(n16674) );
  ANDN U16874 ( .B(n16677), .A(n16678), .Z(n16676) );
  XOR U16875 ( .A(n16679), .B(n16680), .Z(n13976) );
  XNOR U16876 ( .A(n16634), .B(n16658), .Z(n16680) );
  XNOR U16877 ( .A(n16681), .B(n16682), .Z(n16658) );
  XNOR U16878 ( .A(n16683), .B(n16684), .Z(n16682) );
  OR U16879 ( .A(n16685), .B(n16686), .Z(n16684) );
  XNOR U16880 ( .A(n16687), .B(n16688), .Z(n16679) );
  XOR U16881 ( .A(n16689), .B(n16690), .Z(n16688) );
  ANDN U16882 ( .B(n16691), .A(n16692), .Z(n16690) );
  XNOR U16883 ( .A(n16693), .B(n16694), .Z(n13522) );
  XNOR U16884 ( .A(n16636), .B(n16664), .Z(n16694) );
  XNOR U16885 ( .A(n16695), .B(n16696), .Z(n16664) );
  XNOR U16886 ( .A(n16697), .B(n16698), .Z(n16696) );
  OR U16887 ( .A(n16699), .B(n16700), .Z(n16698) );
  XNOR U16888 ( .A(n16701), .B(n16702), .Z(n16693) );
  XOR U16889 ( .A(n16703), .B(n16704), .Z(n16702) );
  ANDN U16890 ( .B(n16705), .A(n16706), .Z(n16704) );
  XNOR U16891 ( .A(n12171), .B(n16707), .Z(n16667) );
  XNOR U16892 ( .A(key[765]), .B(n13544), .Z(n16707) );
  IV U16893 ( .A(n13971), .Z(n12171) );
  XNOR U16894 ( .A(n16708), .B(n16709), .Z(n13971) );
  IV U16895 ( .A(n16649), .Z(n14706) );
  XNOR U16896 ( .A(n16623), .B(n16710), .Z(n16649) );
  XOR U16897 ( .A(n16711), .B(n16712), .Z(n16631) );
  XNOR U16898 ( .A(n14690), .B(n13967), .Z(n16712) );
  XOR U16899 ( .A(n13984), .B(n13532), .Z(n13967) );
  XNOR U16900 ( .A(n16713), .B(n16714), .Z(n13532) );
  XOR U16901 ( .A(n16715), .B(n16672), .Z(n16714) );
  XNOR U16902 ( .A(n16716), .B(n16717), .Z(n16672) );
  XNOR U16903 ( .A(n16718), .B(n16719), .Z(n16717) );
  NANDN U16904 ( .A(n16720), .B(n16721), .Z(n16719) );
  XOR U16905 ( .A(n16722), .B(n16723), .Z(n16713) );
  XNOR U16906 ( .A(n16724), .B(n16725), .Z(n14690) );
  XOR U16907 ( .A(n13560), .B(n13531), .Z(n16725) );
  XNOR U16908 ( .A(n13550), .B(n13982), .Z(n13531) );
  XNOR U16909 ( .A(n16726), .B(n16634), .Z(n13982) );
  XNOR U16910 ( .A(n16681), .B(n16727), .Z(n16634) );
  XOR U16911 ( .A(n16728), .B(n16729), .Z(n16727) );
  NOR U16912 ( .A(n16730), .B(n16731), .Z(n16728) );
  XNOR U16913 ( .A(n16732), .B(n16733), .Z(n16681) );
  XNOR U16914 ( .A(n16734), .B(n16735), .Z(n16733) );
  NAND U16915 ( .A(n16736), .B(n16737), .Z(n16735) );
  XNOR U16916 ( .A(n16738), .B(n16636), .Z(n13550) );
  XNOR U16917 ( .A(n16695), .B(n16739), .Z(n16636) );
  XOR U16918 ( .A(n16740), .B(n16741), .Z(n16739) );
  NOR U16919 ( .A(n16742), .B(n16743), .Z(n16740) );
  XNOR U16920 ( .A(n16744), .B(n16745), .Z(n16695) );
  XNOR U16921 ( .A(n16746), .B(n16747), .Z(n16745) );
  NAND U16922 ( .A(n16748), .B(n16749), .Z(n16747) );
  XOR U16923 ( .A(n12154), .B(n16750), .Z(n16724) );
  XNOR U16924 ( .A(key[760]), .B(n16751), .Z(n16750) );
  XOR U16925 ( .A(n16709), .B(n16752), .Z(n12154) );
  XNOR U16926 ( .A(n12165), .B(n16753), .Z(n16711) );
  XOR U16927 ( .A(key[766]), .B(n13540), .Z(n16753) );
  XOR U16928 ( .A(n16663), .B(n16754), .Z(n13540) );
  XNOR U16929 ( .A(n13974), .B(n12136), .Z(n12165) );
  XNOR U16930 ( .A(n14002), .B(n13981), .Z(n12136) );
  XNOR U16931 ( .A(n16755), .B(n16756), .Z(n13981) );
  XNOR U16932 ( .A(n16709), .B(n16640), .Z(n16756) );
  XNOR U16933 ( .A(n16757), .B(n16758), .Z(n16640) );
  XNOR U16934 ( .A(n16759), .B(n16760), .Z(n16758) );
  NANDN U16935 ( .A(n16761), .B(n16762), .Z(n16760) );
  XOR U16936 ( .A(n16763), .B(n16764), .Z(n16709) );
  XNOR U16937 ( .A(n16765), .B(n16766), .Z(n16755) );
  XOR U16938 ( .A(n13544), .B(n13968), .Z(n13974) );
  IV U16939 ( .A(n13536), .Z(n13968) );
  XNOR U16940 ( .A(n16657), .B(n16767), .Z(n13536) );
  XOR U16941 ( .A(n16723), .B(n16768), .Z(n13544) );
  XOR U16942 ( .A(n16769), .B(n16770), .Z(n16628) );
  XNOR U16943 ( .A(n13994), .B(n16771), .Z(n16770) );
  XNOR U16944 ( .A(n12147), .B(n16651), .Z(n16771) );
  IV U16945 ( .A(n16622), .Z(n16651) );
  XNOR U16946 ( .A(n16772), .B(n16773), .Z(n16622) );
  XNOR U16947 ( .A(n13570), .B(n12153), .Z(n16773) );
  XOR U16948 ( .A(n13998), .B(n13560), .Z(n12153) );
  XNOR U16949 ( .A(n16715), .B(n16774), .Z(n13560) );
  XOR U16950 ( .A(n16775), .B(n16776), .Z(n16723) );
  IV U16951 ( .A(n13552), .Z(n13998) );
  XNOR U16952 ( .A(n16657), .B(n16777), .Z(n13552) );
  XOR U16953 ( .A(n16778), .B(n16660), .Z(n16777) );
  XOR U16954 ( .A(n16779), .B(n16726), .Z(n16657) );
  XOR U16955 ( .A(n12160), .B(n16780), .Z(n16772) );
  XNOR U16956 ( .A(key[761]), .B(n13549), .Z(n16780) );
  XNOR U16957 ( .A(n16663), .B(n16781), .Z(n13549) );
  XOR U16958 ( .A(n16782), .B(n16666), .Z(n16781) );
  XOR U16959 ( .A(n16783), .B(n16738), .Z(n16663) );
  XNOR U16960 ( .A(n14002), .B(n12125), .Z(n12147) );
  XNOR U16961 ( .A(n16641), .B(n12160), .Z(n12125) );
  XNOR U16962 ( .A(n16763), .B(n16765), .Z(n12160) );
  XOR U16963 ( .A(n16641), .B(n16763), .Z(n14002) );
  XNOR U16964 ( .A(n16784), .B(n16785), .Z(n16763) );
  XOR U16965 ( .A(n16786), .B(n16759), .Z(n16785) );
  OR U16966 ( .A(n16787), .B(n16788), .Z(n16759) );
  ANDN U16967 ( .B(n16789), .A(n16790), .Z(n16786) );
  XNOR U16968 ( .A(n16757), .B(n16791), .Z(n16641) );
  XOR U16969 ( .A(n16792), .B(n16793), .Z(n16791) );
  NOR U16970 ( .A(n16794), .B(n16795), .Z(n16792) );
  XNOR U16971 ( .A(n16784), .B(n16796), .Z(n16757) );
  XNOR U16972 ( .A(n16797), .B(n16798), .Z(n16796) );
  NAND U16973 ( .A(n16799), .B(n16800), .Z(n16798) );
  XNOR U16974 ( .A(n16751), .B(n13518), .Z(n13994) );
  XOR U16975 ( .A(n16673), .B(n13570), .Z(n13518) );
  IV U16976 ( .A(n13984), .Z(n16751) );
  XOR U16977 ( .A(n16673), .B(n16801), .Z(n13984) );
  XNOR U16978 ( .A(n16716), .B(n16802), .Z(n16673) );
  XOR U16979 ( .A(n16803), .B(n16804), .Z(n16802) );
  NOR U16980 ( .A(n16805), .B(n16806), .Z(n16803) );
  XNOR U16981 ( .A(n16807), .B(n16808), .Z(n16716) );
  XNOR U16982 ( .A(n16809), .B(n16810), .Z(n16808) );
  NAND U16983 ( .A(n16811), .B(n16812), .Z(n16810) );
  XNOR U16984 ( .A(n12149), .B(n16813), .Z(n16769) );
  XNOR U16985 ( .A(key[763]), .B(n13572), .Z(n16813) );
  XOR U16986 ( .A(n16814), .B(n16815), .Z(n13572) );
  XNOR U16987 ( .A(n16783), .B(n16754), .Z(n16815) );
  XNOR U16988 ( .A(n16816), .B(n16817), .Z(n16754) );
  XNOR U16989 ( .A(n16818), .B(n16703), .Z(n16817) );
  ANDN U16990 ( .B(n16819), .A(n16820), .Z(n16703) );
  NOR U16991 ( .A(n16821), .B(n16743), .Z(n16818) );
  XNOR U16992 ( .A(n16701), .B(n16822), .Z(n16783) );
  XNOR U16993 ( .A(n16823), .B(n16824), .Z(n16822) );
  NANDN U16994 ( .A(n16825), .B(n16826), .Z(n16824) );
  XNOR U16995 ( .A(n16782), .B(n16666), .Z(n16814) );
  XNOR U16996 ( .A(n16823), .B(n16828), .Z(n16827) );
  NANDN U16997 ( .A(n16699), .B(n16829), .Z(n16828) );
  OR U16998 ( .A(n16830), .B(n16831), .Z(n16823) );
  XNOR U16999 ( .A(n16701), .B(n16832), .Z(n16816) );
  XNOR U17000 ( .A(n16833), .B(n16834), .Z(n16832) );
  NAND U17001 ( .A(n16835), .B(n16748), .Z(n16834) );
  XOR U17002 ( .A(n16836), .B(n16833), .Z(n16701) );
  NANDN U17003 ( .A(n16837), .B(n16838), .Z(n16833) );
  AND U17004 ( .A(n16839), .B(n16840), .Z(n16836) );
  XNOR U17005 ( .A(n13557), .B(n13569), .Z(n12149) );
  XOR U17006 ( .A(n16841), .B(n16842), .Z(n13569) );
  XNOR U17007 ( .A(n16779), .B(n16767), .Z(n16842) );
  XNOR U17008 ( .A(n16843), .B(n16844), .Z(n16767) );
  XNOR U17009 ( .A(n16845), .B(n16689), .Z(n16844) );
  ANDN U17010 ( .B(n16846), .A(n16847), .Z(n16689) );
  NOR U17011 ( .A(n16848), .B(n16731), .Z(n16845) );
  XNOR U17012 ( .A(n16687), .B(n16849), .Z(n16779) );
  XNOR U17013 ( .A(n16850), .B(n16851), .Z(n16849) );
  NANDN U17014 ( .A(n16852), .B(n16853), .Z(n16851) );
  XNOR U17015 ( .A(n16778), .B(n16660), .Z(n16841) );
  XNOR U17016 ( .A(n16850), .B(n16855), .Z(n16854) );
  NANDN U17017 ( .A(n16685), .B(n16856), .Z(n16855) );
  OR U17018 ( .A(n16857), .B(n16858), .Z(n16850) );
  XNOR U17019 ( .A(n16687), .B(n16859), .Z(n16843) );
  XNOR U17020 ( .A(n16860), .B(n16861), .Z(n16859) );
  NAND U17021 ( .A(n16862), .B(n16736), .Z(n16861) );
  XOR U17022 ( .A(n16863), .B(n16860), .Z(n16687) );
  NANDN U17023 ( .A(n16864), .B(n16865), .Z(n16860) );
  AND U17024 ( .A(n16866), .B(n16867), .Z(n16863) );
  XOR U17025 ( .A(n16868), .B(n16869), .Z(n16623) );
  XNOR U17026 ( .A(n13557), .B(n13997), .Z(n16869) );
  IV U17027 ( .A(n12161), .Z(n13997) );
  XOR U17028 ( .A(n13563), .B(n13570), .Z(n12161) );
  XOR U17029 ( .A(n16775), .B(n16715), .Z(n13570) );
  IV U17030 ( .A(n16801), .Z(n16775) );
  XNOR U17031 ( .A(n16807), .B(n16870), .Z(n16801) );
  XOR U17032 ( .A(n16871), .B(n16718), .Z(n16870) );
  OR U17033 ( .A(n16872), .B(n16873), .Z(n16718) );
  ANDN U17034 ( .B(n16874), .A(n16875), .Z(n16871) );
  XOR U17035 ( .A(n16659), .B(n16726), .Z(n13563) );
  XOR U17036 ( .A(n16732), .B(n16876), .Z(n16726) );
  XOR U17037 ( .A(n16877), .B(n16683), .Z(n16876) );
  OR U17038 ( .A(n16878), .B(n16857), .Z(n16683) );
  XNOR U17039 ( .A(n16685), .B(n16852), .Z(n16857) );
  NOR U17040 ( .A(n16879), .B(n16852), .Z(n16877) );
  IV U17041 ( .A(n16778), .Z(n16659) );
  XNOR U17042 ( .A(n16732), .B(n16880), .Z(n16778) );
  XNOR U17043 ( .A(n16729), .B(n16881), .Z(n16880) );
  NAND U17044 ( .A(n16882), .B(n16691), .Z(n16881) );
  XNOR U17045 ( .A(n16731), .B(n16691), .Z(n16846) );
  XOR U17046 ( .A(n16884), .B(n16734), .Z(n16732) );
  OR U17047 ( .A(n16864), .B(n16885), .Z(n16734) );
  XNOR U17048 ( .A(n16866), .B(n16736), .Z(n16864) );
  XNOR U17049 ( .A(n16852), .B(n16691), .Z(n16736) );
  XOR U17050 ( .A(n16886), .B(n16887), .Z(n16691) );
  NANDN U17051 ( .A(n16888), .B(n16889), .Z(n16887) );
  XNOR U17052 ( .A(n16890), .B(n16891), .Z(n16852) );
  OR U17053 ( .A(n16888), .B(n16892), .Z(n16891) );
  ANDN U17054 ( .B(n16866), .A(n16893), .Z(n16884) );
  XOR U17055 ( .A(n16685), .B(n16731), .Z(n16866) );
  XOR U17056 ( .A(n16894), .B(n16886), .Z(n16731) );
  NANDN U17057 ( .A(n16895), .B(n16896), .Z(n16886) );
  ANDN U17058 ( .B(n16897), .A(n16898), .Z(n16894) );
  NANDN U17059 ( .A(n16895), .B(n16900), .Z(n16890) );
  XOR U17060 ( .A(n16901), .B(n16888), .Z(n16895) );
  XNOR U17061 ( .A(n16902), .B(n16903), .Z(n16888) );
  XOR U17062 ( .A(n16904), .B(n16897), .Z(n16903) );
  XNOR U17063 ( .A(n16905), .B(n16906), .Z(n16902) );
  XNOR U17064 ( .A(n16907), .B(n16908), .Z(n16906) );
  ANDN U17065 ( .B(n16897), .A(n16909), .Z(n16907) );
  IV U17066 ( .A(n16910), .Z(n16897) );
  ANDN U17067 ( .B(n16901), .A(n16909), .Z(n16899) );
  IV U17068 ( .A(n16905), .Z(n16909) );
  IV U17069 ( .A(n16898), .Z(n16901) );
  XNOR U17070 ( .A(n16904), .B(n16911), .Z(n16898) );
  XOR U17071 ( .A(n16912), .B(n16908), .Z(n16911) );
  NAND U17072 ( .A(n16900), .B(n16896), .Z(n16908) );
  XNOR U17073 ( .A(n16889), .B(n16910), .Z(n16896) );
  XOR U17074 ( .A(n16913), .B(n16914), .Z(n16910) );
  XOR U17075 ( .A(n16915), .B(n16916), .Z(n16914) );
  XNOR U17076 ( .A(n16853), .B(n16917), .Z(n16916) );
  XNOR U17077 ( .A(n16918), .B(n16919), .Z(n16913) );
  XNOR U17078 ( .A(n16920), .B(n16921), .Z(n16919) );
  ANDN U17079 ( .B(n16856), .A(n16686), .Z(n16920) );
  XNOR U17080 ( .A(n16905), .B(n16892), .Z(n16900) );
  XOR U17081 ( .A(n16922), .B(n16923), .Z(n16905) );
  XNOR U17082 ( .A(n16924), .B(n16917), .Z(n16923) );
  XOR U17083 ( .A(n16925), .B(n16926), .Z(n16917) );
  XNOR U17084 ( .A(n16927), .B(n16928), .Z(n16926) );
  NAND U17085 ( .A(n16737), .B(n16862), .Z(n16928) );
  XNOR U17086 ( .A(n16929), .B(n16930), .Z(n16922) );
  ANDN U17087 ( .B(n16931), .A(n16730), .Z(n16929) );
  ANDN U17088 ( .B(n16889), .A(n16892), .Z(n16912) );
  XOR U17089 ( .A(n16892), .B(n16889), .Z(n16904) );
  XNOR U17090 ( .A(n16932), .B(n16933), .Z(n16889) );
  XNOR U17091 ( .A(n16925), .B(n16934), .Z(n16933) );
  XNOR U17092 ( .A(n16924), .B(n16856), .Z(n16934) );
  XNOR U17093 ( .A(n16935), .B(n16936), .Z(n16932) );
  XNOR U17094 ( .A(n16937), .B(n16921), .Z(n16936) );
  OR U17095 ( .A(n16858), .B(n16878), .Z(n16921) );
  XNOR U17096 ( .A(n16935), .B(n16918), .Z(n16878) );
  XNOR U17097 ( .A(n16856), .B(n16853), .Z(n16858) );
  ANDN U17098 ( .B(n16853), .A(n16879), .Z(n16937) );
  XOR U17099 ( .A(n16938), .B(n16939), .Z(n16892) );
  XOR U17100 ( .A(n16925), .B(n16915), .Z(n16939) );
  XOR U17101 ( .A(n16882), .B(n16692), .Z(n16915) );
  XOR U17102 ( .A(n16940), .B(n16927), .Z(n16925) );
  NANDN U17103 ( .A(n16885), .B(n16865), .Z(n16927) );
  XOR U17104 ( .A(n16867), .B(n16862), .Z(n16865) );
  XNOR U17105 ( .A(n16931), .B(n16941), .Z(n16853) );
  XNOR U17106 ( .A(n16942), .B(n16943), .Z(n16941) );
  XOR U17107 ( .A(n16893), .B(n16737), .Z(n16885) );
  XNOR U17108 ( .A(n16879), .B(n16882), .Z(n16737) );
  IV U17109 ( .A(n16918), .Z(n16879) );
  XOR U17110 ( .A(n16944), .B(n16945), .Z(n16918) );
  XOR U17111 ( .A(n16946), .B(n16947), .Z(n16945) );
  XOR U17112 ( .A(n16935), .B(n16948), .Z(n16944) );
  ANDN U17113 ( .B(n16867), .A(n16893), .Z(n16940) );
  XNOR U17114 ( .A(n16935), .B(n16949), .Z(n16893) );
  XOR U17115 ( .A(n16931), .B(n16856), .Z(n16867) );
  XNOR U17116 ( .A(n16950), .B(n16951), .Z(n16856) );
  XOR U17117 ( .A(n16952), .B(n16947), .Z(n16951) );
  XNOR U17118 ( .A(n16953), .B(n16519), .Z(n16947) );
  XOR U17119 ( .A(n16954), .B(n16955), .Z(n16519) );
  XOR U17120 ( .A(n15441), .B(n16956), .Z(n16955) );
  XNOR U17121 ( .A(n16958), .B(n16959), .Z(n16953) );
  XNOR U17122 ( .A(key[556]), .B(n16534), .Z(n16959) );
  IV U17123 ( .A(n16960), .Z(n16534) );
  IV U17124 ( .A(n16848), .Z(n16931) );
  XOR U17125 ( .A(n16924), .B(n16961), .Z(n16938) );
  XNOR U17126 ( .A(n16962), .B(n16930), .Z(n16961) );
  OR U17127 ( .A(n16847), .B(n16883), .Z(n16930) );
  XNOR U17128 ( .A(n16949), .B(n16882), .Z(n16883) );
  XNOR U17129 ( .A(n16848), .B(n16692), .Z(n16847) );
  ANDN U17130 ( .B(n16882), .A(n16692), .Z(n16962) );
  XOR U17131 ( .A(n16950), .B(n16963), .Z(n16692) );
  XOR U17132 ( .A(n16942), .B(n16964), .Z(n16963) );
  XOR U17133 ( .A(n16952), .B(n16950), .Z(n16882) );
  XNOR U17134 ( .A(n16730), .B(n16848), .Z(n16924) );
  XOR U17135 ( .A(n16950), .B(n16965), .Z(n16848) );
  XNOR U17136 ( .A(n16952), .B(n16946), .Z(n16965) );
  XOR U17137 ( .A(n16966), .B(n16967), .Z(n16946) );
  XOR U17138 ( .A(n15493), .B(n16517), .Z(n16967) );
  XOR U17139 ( .A(n16968), .B(n15459), .Z(n16517) );
  XNOR U17140 ( .A(n16969), .B(n16957), .Z(n15493) );
  XNOR U17141 ( .A(key[559]), .B(n16506), .Z(n16966) );
  XNOR U17142 ( .A(n16970), .B(n16971), .Z(n16950) );
  XNOR U17143 ( .A(n16503), .B(n16510), .Z(n16971) );
  XOR U17144 ( .A(n15454), .B(n16972), .Z(n16510) );
  XNOR U17145 ( .A(n15471), .B(n16973), .Z(n16970) );
  XOR U17146 ( .A(key[557]), .B(n16522), .Z(n16973) );
  IV U17147 ( .A(n16949), .Z(n16730) );
  XNOR U17148 ( .A(n16943), .B(n16974), .Z(n16949) );
  XOR U17149 ( .A(n16948), .B(n16964), .Z(n16974) );
  IV U17150 ( .A(n16952), .Z(n16964) );
  XOR U17151 ( .A(n16975), .B(n16976), .Z(n16952) );
  XNOR U17152 ( .A(n16502), .B(n16686), .Z(n16976) );
  IV U17153 ( .A(n16935), .Z(n16686) );
  XOR U17154 ( .A(n16977), .B(n16978), .Z(n16935) );
  XOR U17155 ( .A(n16531), .B(n15485), .Z(n16978) );
  XOR U17156 ( .A(n15457), .B(n16979), .Z(n16977) );
  XNOR U17157 ( .A(key[552]), .B(n16980), .Z(n16979) );
  XOR U17158 ( .A(n16981), .B(n16516), .Z(n16502) );
  XOR U17159 ( .A(n16957), .B(n16982), .Z(n16516) );
  XNOR U17160 ( .A(n16983), .B(n16984), .Z(n16975) );
  XNOR U17161 ( .A(key[558]), .B(n15450), .Z(n16984) );
  XOR U17162 ( .A(n16985), .B(n16986), .Z(n16948) );
  XNOR U17163 ( .A(n16942), .B(n16987), .Z(n16986) );
  XNOR U17164 ( .A(n16527), .B(n16525), .Z(n16987) );
  XOR U17165 ( .A(n16957), .B(n16520), .Z(n16525) );
  XOR U17166 ( .A(n16988), .B(n16989), .Z(n16942) );
  XNOR U17167 ( .A(n16495), .B(n16530), .Z(n16989) );
  XNOR U17168 ( .A(n15467), .B(n16990), .Z(n16988) );
  XOR U17169 ( .A(key[553]), .B(n15491), .Z(n16990) );
  XNOR U17170 ( .A(n16991), .B(n16992), .Z(n16985) );
  XNOR U17171 ( .A(key[555]), .B(n15465), .Z(n16992) );
  XOR U17172 ( .A(n16993), .B(n16994), .Z(n16943) );
  XOR U17173 ( .A(n16533), .B(n16494), .Z(n16994) );
  IV U17174 ( .A(n16995), .Z(n16494) );
  XNOR U17175 ( .A(n15480), .B(n16996), .Z(n16993) );
  XNOR U17176 ( .A(key[554]), .B(n15488), .Z(n16996) );
  XOR U17177 ( .A(n16997), .B(n16998), .Z(n13557) );
  XOR U17178 ( .A(n16715), .B(n16768), .Z(n16998) );
  XNOR U17179 ( .A(n16999), .B(n17000), .Z(n16768) );
  XNOR U17180 ( .A(n17001), .B(n16675), .Z(n17000) );
  ANDN U17181 ( .B(n17002), .A(n17003), .Z(n16675) );
  NOR U17182 ( .A(n17004), .B(n16806), .Z(n17001) );
  XOR U17183 ( .A(n16807), .B(n17005), .Z(n16715) );
  XNOR U17184 ( .A(n16804), .B(n17006), .Z(n17005) );
  NANDN U17185 ( .A(n17007), .B(n16677), .Z(n17006) );
  XNOR U17186 ( .A(n16806), .B(n16677), .Z(n17002) );
  XOR U17187 ( .A(n17009), .B(n16809), .Z(n16807) );
  OR U17188 ( .A(n17010), .B(n17011), .Z(n16809) );
  ANDN U17189 ( .B(n17012), .A(n17013), .Z(n17009) );
  XOR U17190 ( .A(n16722), .B(n16776), .Z(n16997) );
  XOR U17191 ( .A(n16671), .B(n17014), .Z(n16776) );
  XNOR U17192 ( .A(n17015), .B(n17016), .Z(n17014) );
  NANDN U17193 ( .A(n17017), .B(n17018), .Z(n17016) );
  XNOR U17194 ( .A(n17015), .B(n17020), .Z(n17019) );
  NANDN U17195 ( .A(n17021), .B(n16721), .Z(n17020) );
  OR U17196 ( .A(n16872), .B(n17022), .Z(n17015) );
  XNOR U17197 ( .A(n16721), .B(n17018), .Z(n16872) );
  XNOR U17198 ( .A(n16671), .B(n17023), .Z(n16999) );
  XNOR U17199 ( .A(n17024), .B(n17025), .Z(n17023) );
  NAND U17200 ( .A(n17026), .B(n16811), .Z(n17025) );
  XOR U17201 ( .A(n17027), .B(n17024), .Z(n16671) );
  NANDN U17202 ( .A(n17010), .B(n17028), .Z(n17024) );
  XOR U17203 ( .A(n17013), .B(n16811), .Z(n17010) );
  XOR U17204 ( .A(n17018), .B(n16677), .Z(n16811) );
  XOR U17205 ( .A(n17029), .B(n17030), .Z(n16677) );
  NANDN U17206 ( .A(n17031), .B(n17032), .Z(n17030) );
  IV U17207 ( .A(n16875), .Z(n17018) );
  XNOR U17208 ( .A(n17033), .B(n17034), .Z(n16875) );
  NANDN U17209 ( .A(n17031), .B(n17035), .Z(n17034) );
  ANDN U17210 ( .B(n17036), .A(n17013), .Z(n17027) );
  XOR U17211 ( .A(n16806), .B(n16721), .Z(n17013) );
  XNOR U17212 ( .A(n17037), .B(n17033), .Z(n16721) );
  NANDN U17213 ( .A(n17038), .B(n17039), .Z(n17033) );
  XOR U17214 ( .A(n17035), .B(n17040), .Z(n17039) );
  ANDN U17215 ( .B(n17040), .A(n17041), .Z(n17037) );
  XOR U17216 ( .A(n17042), .B(n17029), .Z(n16806) );
  NANDN U17217 ( .A(n17038), .B(n17043), .Z(n17029) );
  XOR U17218 ( .A(n17044), .B(n17032), .Z(n17043) );
  XNOR U17219 ( .A(n17045), .B(n17046), .Z(n17031) );
  XOR U17220 ( .A(n17047), .B(n17048), .Z(n17046) );
  XNOR U17221 ( .A(n17049), .B(n17050), .Z(n17045) );
  XNOR U17222 ( .A(n17051), .B(n17052), .Z(n17050) );
  ANDN U17223 ( .B(n17044), .A(n17048), .Z(n17051) );
  ANDN U17224 ( .B(n17044), .A(n17041), .Z(n17042) );
  XNOR U17225 ( .A(n17047), .B(n17053), .Z(n17041) );
  XOR U17226 ( .A(n17054), .B(n17052), .Z(n17053) );
  NAND U17227 ( .A(n17055), .B(n17056), .Z(n17052) );
  XNOR U17228 ( .A(n17049), .B(n17032), .Z(n17056) );
  IV U17229 ( .A(n17044), .Z(n17049) );
  XNOR U17230 ( .A(n17035), .B(n17048), .Z(n17055) );
  IV U17231 ( .A(n17040), .Z(n17048) );
  XOR U17232 ( .A(n17057), .B(n17058), .Z(n17040) );
  XNOR U17233 ( .A(n17059), .B(n17060), .Z(n17058) );
  XNOR U17234 ( .A(n17061), .B(n17062), .Z(n17057) );
  NOR U17235 ( .A(n17004), .B(n16805), .Z(n17061) );
  AND U17236 ( .A(n17032), .B(n17035), .Z(n17054) );
  XNOR U17237 ( .A(n17032), .B(n17035), .Z(n17047) );
  XNOR U17238 ( .A(n17063), .B(n17064), .Z(n17035) );
  XNOR U17239 ( .A(n17065), .B(n17060), .Z(n17064) );
  XOR U17240 ( .A(n17066), .B(n17067), .Z(n17063) );
  XNOR U17241 ( .A(n17068), .B(n17062), .Z(n17067) );
  OR U17242 ( .A(n17003), .B(n17008), .Z(n17062) );
  XNOR U17243 ( .A(n16805), .B(n17007), .Z(n17008) );
  XNOR U17244 ( .A(n17004), .B(n16678), .Z(n17003) );
  ANDN U17245 ( .B(n17069), .A(n17007), .Z(n17068) );
  XNOR U17246 ( .A(n17070), .B(n17071), .Z(n17032) );
  XNOR U17247 ( .A(n17060), .B(n17072), .Z(n17071) );
  XOR U17248 ( .A(n17021), .B(n17066), .Z(n17072) );
  XNOR U17249 ( .A(n16805), .B(n17073), .Z(n17060) );
  XNOR U17250 ( .A(n17074), .B(n17075), .Z(n17070) );
  XNOR U17251 ( .A(n17076), .B(n17077), .Z(n17075) );
  ANDN U17252 ( .B(n16874), .A(n17017), .Z(n17076) );
  XNOR U17253 ( .A(n17078), .B(n17079), .Z(n17044) );
  XNOR U17254 ( .A(n17065), .B(n17080), .Z(n17079) );
  XNOR U17255 ( .A(n17017), .B(n17059), .Z(n17080) );
  XOR U17256 ( .A(n17066), .B(n17081), .Z(n17059) );
  XNOR U17257 ( .A(n17082), .B(n17083), .Z(n17081) );
  NAND U17258 ( .A(n16812), .B(n17026), .Z(n17083) );
  XNOR U17259 ( .A(n17084), .B(n17082), .Z(n17066) );
  NANDN U17260 ( .A(n17011), .B(n17028), .Z(n17082) );
  XOR U17261 ( .A(n17036), .B(n17026), .Z(n17028) );
  XNOR U17262 ( .A(n17085), .B(n16678), .Z(n17026) );
  XOR U17263 ( .A(n17086), .B(n16812), .Z(n17011) );
  XOR U17264 ( .A(n16874), .B(n17087), .Z(n16812) );
  ANDN U17265 ( .B(n17036), .A(n17086), .Z(n17084) );
  IV U17266 ( .A(n17012), .Z(n17086) );
  XOR U17267 ( .A(n16720), .B(n16805), .Z(n17012) );
  XOR U17268 ( .A(n17088), .B(n17089), .Z(n16805) );
  XNOR U17269 ( .A(n17090), .B(n17091), .Z(n17089) );
  XOR U17270 ( .A(n17087), .B(n17069), .Z(n17065) );
  IV U17271 ( .A(n16678), .Z(n17069) );
  XOR U17272 ( .A(n17092), .B(n17093), .Z(n16678) );
  XNOR U17273 ( .A(n17094), .B(n17091), .Z(n17093) );
  IV U17274 ( .A(n17007), .Z(n17087) );
  XOR U17275 ( .A(n17091), .B(n17095), .Z(n17007) );
  XNOR U17276 ( .A(n16874), .B(n17096), .Z(n17078) );
  XNOR U17277 ( .A(n17097), .B(n17077), .Z(n17096) );
  OR U17278 ( .A(n17022), .B(n16873), .Z(n17077) );
  XNOR U17279 ( .A(n17074), .B(n16874), .Z(n16873) );
  XOR U17280 ( .A(n17021), .B(n17085), .Z(n17022) );
  IV U17281 ( .A(n17017), .Z(n17085) );
  XOR U17282 ( .A(n17073), .B(n17098), .Z(n17017) );
  XNOR U17283 ( .A(n17094), .B(n17088), .Z(n17098) );
  XOR U17284 ( .A(n17099), .B(n17100), .Z(n17088) );
  XNOR U17285 ( .A(n15343), .B(n17101), .Z(n17100) );
  XOR U17286 ( .A(n16039), .B(n17102), .Z(n15343) );
  IV U17287 ( .A(n17103), .Z(n16039) );
  XOR U17288 ( .A(key[594]), .B(n15347), .Z(n17099) );
  ANDN U17289 ( .B(n17104), .A(n16720), .Z(n17097) );
  XOR U17290 ( .A(n17105), .B(n17106), .Z(n16874) );
  XNOR U17291 ( .A(n17107), .B(n17108), .Z(n17106) );
  XOR U17292 ( .A(n17074), .B(n17090), .Z(n17105) );
  XOR U17293 ( .A(n17109), .B(n17110), .Z(n17090) );
  XNOR U17294 ( .A(n17094), .B(n17111), .Z(n17110) );
  XOR U17295 ( .A(n17112), .B(n16029), .Z(n17111) );
  XNOR U17296 ( .A(n16067), .B(n16047), .Z(n16029) );
  IV U17297 ( .A(n17113), .Z(n16047) );
  XOR U17298 ( .A(n17114), .B(n17115), .Z(n17094) );
  XNOR U17299 ( .A(n17116), .B(n15307), .Z(n17115) );
  XOR U17300 ( .A(key[593]), .B(n15355), .Z(n17114) );
  XNOR U17301 ( .A(n15308), .B(n17117), .Z(n17109) );
  XNOR U17302 ( .A(key[595]), .B(n17102), .Z(n17117) );
  XOR U17303 ( .A(n17104), .B(n17073), .Z(n17036) );
  IV U17304 ( .A(n17004), .Z(n17073) );
  XOR U17305 ( .A(n17092), .B(n17118), .Z(n17004) );
  XOR U17306 ( .A(n17091), .B(n17108), .Z(n17118) );
  XNOR U17307 ( .A(n17119), .B(n17120), .Z(n17108) );
  XNOR U17308 ( .A(n17121), .B(n17122), .Z(n17120) );
  XOR U17309 ( .A(key[599]), .B(n16067), .Z(n17119) );
  IV U17310 ( .A(n17021), .Z(n17104) );
  XOR U17311 ( .A(n17092), .B(n17123), .Z(n17021) );
  XOR U17312 ( .A(n17091), .B(n17107), .Z(n17123) );
  XNOR U17313 ( .A(n17124), .B(n17125), .Z(n17107) );
  XOR U17314 ( .A(n17126), .B(n16046), .Z(n17125) );
  XNOR U17315 ( .A(n16067), .B(n16075), .Z(n16046) );
  XOR U17316 ( .A(n17127), .B(n17128), .Z(n17124) );
  XNOR U17317 ( .A(key[596]), .B(n16048), .Z(n17128) );
  XOR U17318 ( .A(n17129), .B(n17130), .Z(n17091) );
  XOR U17319 ( .A(n16060), .B(n16720), .Z(n17130) );
  IV U17320 ( .A(n17074), .Z(n16720) );
  XOR U17321 ( .A(n17131), .B(n17132), .Z(n17074) );
  XOR U17322 ( .A(n17133), .B(n17116), .Z(n15346) );
  XNOR U17323 ( .A(key[592]), .B(n17134), .Z(n17131) );
  XOR U17324 ( .A(n16067), .B(n16055), .Z(n16060) );
  XOR U17325 ( .A(n17135), .B(n17136), .Z(n17129) );
  XNOR U17326 ( .A(key[598]), .B(n17137), .Z(n17136) );
  IV U17327 ( .A(n17095), .Z(n17092) );
  XOR U17328 ( .A(n17138), .B(n17139), .Z(n17095) );
  XNOR U17329 ( .A(n16076), .B(n17140), .Z(n17139) );
  XNOR U17330 ( .A(key[597]), .B(n16070), .Z(n17138) );
  XOR U17331 ( .A(n16077), .B(n17137), .Z(n16070) );
  XNOR U17332 ( .A(n13561), .B(n17141), .Z(n16868) );
  XOR U17333 ( .A(key[762]), .B(n12157), .Z(n17141) );
  XNOR U17334 ( .A(n17142), .B(n16752), .Z(n12157) );
  XOR U17335 ( .A(n16765), .B(n16766), .Z(n16752) );
  XNOR U17336 ( .A(n17143), .B(n17144), .Z(n16766) );
  XNOR U17337 ( .A(n17145), .B(n17146), .Z(n17144) );
  NANDN U17338 ( .A(n17147), .B(n16762), .Z(n17146) );
  XOR U17339 ( .A(n16784), .B(n17148), .Z(n16765) );
  XNOR U17340 ( .A(n16793), .B(n17149), .Z(n17148) );
  NANDN U17341 ( .A(n17150), .B(n16645), .Z(n17149) );
  NANDN U17342 ( .A(n17151), .B(n17152), .Z(n16793) );
  XOR U17343 ( .A(n17153), .B(n16797), .Z(n16784) );
  OR U17344 ( .A(n17154), .B(n17155), .Z(n16797) );
  ANDN U17345 ( .B(n17156), .A(n17157), .Z(n17153) );
  XOR U17346 ( .A(n16708), .B(n16764), .Z(n17142) );
  XOR U17347 ( .A(n16639), .B(n17158), .Z(n16764) );
  XNOR U17348 ( .A(n17145), .B(n17159), .Z(n17158) );
  NANDN U17349 ( .A(n17160), .B(n17161), .Z(n17159) );
  OR U17350 ( .A(n16787), .B(n17162), .Z(n17145) );
  XNOR U17351 ( .A(n16762), .B(n17161), .Z(n16787) );
  XNOR U17352 ( .A(n17164), .B(n16643), .Z(n17163) );
  ANDN U17353 ( .B(n17152), .A(n17165), .Z(n16643) );
  XNOR U17354 ( .A(n16795), .B(n16645), .Z(n17152) );
  NOR U17355 ( .A(n17166), .B(n16795), .Z(n17164) );
  XNOR U17356 ( .A(n16639), .B(n17167), .Z(n17143) );
  XNOR U17357 ( .A(n17168), .B(n17169), .Z(n17167) );
  NAND U17358 ( .A(n17170), .B(n16799), .Z(n17169) );
  XOR U17359 ( .A(n17171), .B(n17168), .Z(n16639) );
  NANDN U17360 ( .A(n17154), .B(n17172), .Z(n17168) );
  XOR U17361 ( .A(n17157), .B(n16799), .Z(n17154) );
  XOR U17362 ( .A(n17161), .B(n16645), .Z(n16799) );
  XOR U17363 ( .A(n17173), .B(n17174), .Z(n16645) );
  NANDN U17364 ( .A(n17175), .B(n17176), .Z(n17174) );
  IV U17365 ( .A(n16790), .Z(n17161) );
  XNOR U17366 ( .A(n17177), .B(n17178), .Z(n16790) );
  NANDN U17367 ( .A(n17175), .B(n17179), .Z(n17178) );
  ANDN U17368 ( .B(n17180), .A(n17157), .Z(n17171) );
  XOR U17369 ( .A(n16795), .B(n16762), .Z(n17157) );
  XNOR U17370 ( .A(n17181), .B(n17177), .Z(n16762) );
  NANDN U17371 ( .A(n17182), .B(n17183), .Z(n17177) );
  XOR U17372 ( .A(n17179), .B(n17184), .Z(n17183) );
  ANDN U17373 ( .B(n17184), .A(n17185), .Z(n17181) );
  XOR U17374 ( .A(n17186), .B(n17173), .Z(n16795) );
  NANDN U17375 ( .A(n17182), .B(n17187), .Z(n17173) );
  XOR U17376 ( .A(n17188), .B(n17176), .Z(n17187) );
  XNOR U17377 ( .A(n17189), .B(n17190), .Z(n17175) );
  XOR U17378 ( .A(n17191), .B(n17192), .Z(n17190) );
  XNOR U17379 ( .A(n17193), .B(n17194), .Z(n17189) );
  XNOR U17380 ( .A(n17195), .B(n17196), .Z(n17194) );
  ANDN U17381 ( .B(n17188), .A(n17192), .Z(n17195) );
  ANDN U17382 ( .B(n17188), .A(n17185), .Z(n17186) );
  XNOR U17383 ( .A(n17191), .B(n17197), .Z(n17185) );
  XOR U17384 ( .A(n17198), .B(n17196), .Z(n17197) );
  NAND U17385 ( .A(n17199), .B(n17200), .Z(n17196) );
  XNOR U17386 ( .A(n17193), .B(n17176), .Z(n17200) );
  IV U17387 ( .A(n17188), .Z(n17193) );
  XNOR U17388 ( .A(n17179), .B(n17192), .Z(n17199) );
  IV U17389 ( .A(n17184), .Z(n17192) );
  XOR U17390 ( .A(n17201), .B(n17202), .Z(n17184) );
  XNOR U17391 ( .A(n17203), .B(n17204), .Z(n17202) );
  XNOR U17392 ( .A(n17205), .B(n17206), .Z(n17201) );
  NOR U17393 ( .A(n17166), .B(n16794), .Z(n17205) );
  AND U17394 ( .A(n17176), .B(n17179), .Z(n17198) );
  XNOR U17395 ( .A(n17176), .B(n17179), .Z(n17191) );
  XNOR U17396 ( .A(n17207), .B(n17208), .Z(n17179) );
  XNOR U17397 ( .A(n17209), .B(n17204), .Z(n17208) );
  XOR U17398 ( .A(n17210), .B(n17211), .Z(n17207) );
  XNOR U17399 ( .A(n17212), .B(n17206), .Z(n17211) );
  OR U17400 ( .A(n17165), .B(n17151), .Z(n17206) );
  XNOR U17401 ( .A(n16794), .B(n17150), .Z(n17151) );
  XNOR U17402 ( .A(n17166), .B(n16646), .Z(n17165) );
  ANDN U17403 ( .B(n17213), .A(n17150), .Z(n17212) );
  XNOR U17404 ( .A(n17214), .B(n17215), .Z(n17176) );
  XNOR U17405 ( .A(n17204), .B(n17216), .Z(n17215) );
  XOR U17406 ( .A(n17147), .B(n17210), .Z(n17216) );
  XNOR U17407 ( .A(n16794), .B(n17217), .Z(n17204) );
  XNOR U17408 ( .A(n17218), .B(n17219), .Z(n17214) );
  XNOR U17409 ( .A(n17220), .B(n17221), .Z(n17219) );
  ANDN U17410 ( .B(n16789), .A(n17160), .Z(n17220) );
  XNOR U17411 ( .A(n17222), .B(n17223), .Z(n17188) );
  XNOR U17412 ( .A(n17209), .B(n17224), .Z(n17223) );
  XNOR U17413 ( .A(n17160), .B(n17203), .Z(n17224) );
  XOR U17414 ( .A(n17210), .B(n17225), .Z(n17203) );
  XNOR U17415 ( .A(n17226), .B(n17227), .Z(n17225) );
  NAND U17416 ( .A(n16800), .B(n17170), .Z(n17227) );
  XNOR U17417 ( .A(n17228), .B(n17226), .Z(n17210) );
  NANDN U17418 ( .A(n17155), .B(n17172), .Z(n17226) );
  XOR U17419 ( .A(n17180), .B(n17170), .Z(n17172) );
  XNOR U17420 ( .A(n17229), .B(n16646), .Z(n17170) );
  XOR U17421 ( .A(n17230), .B(n16800), .Z(n17155) );
  XOR U17422 ( .A(n16789), .B(n17231), .Z(n16800) );
  ANDN U17423 ( .B(n17180), .A(n17230), .Z(n17228) );
  IV U17424 ( .A(n17156), .Z(n17230) );
  XOR U17425 ( .A(n16761), .B(n16794), .Z(n17156) );
  XOR U17426 ( .A(n17232), .B(n17233), .Z(n16794) );
  XNOR U17427 ( .A(n17234), .B(n17235), .Z(n17233) );
  XOR U17428 ( .A(n17231), .B(n17213), .Z(n17209) );
  IV U17429 ( .A(n16646), .Z(n17213) );
  XOR U17430 ( .A(n17236), .B(n17237), .Z(n16646) );
  XNOR U17431 ( .A(n17238), .B(n17235), .Z(n17237) );
  IV U17432 ( .A(n17150), .Z(n17231) );
  XOR U17433 ( .A(n17235), .B(n17239), .Z(n17150) );
  XNOR U17434 ( .A(n16789), .B(n17240), .Z(n17222) );
  XNOR U17435 ( .A(n17241), .B(n17221), .Z(n17240) );
  OR U17436 ( .A(n17162), .B(n16788), .Z(n17221) );
  XNOR U17437 ( .A(n17218), .B(n16789), .Z(n16788) );
  XOR U17438 ( .A(n17147), .B(n17229), .Z(n17162) );
  IV U17439 ( .A(n17160), .Z(n17229) );
  XOR U17440 ( .A(n17217), .B(n17242), .Z(n17160) );
  XNOR U17441 ( .A(n17238), .B(n17232), .Z(n17242) );
  XOR U17442 ( .A(n17243), .B(n17244), .Z(n17232) );
  XOR U17443 ( .A(n16197), .B(n16186), .Z(n17244) );
  XOR U17444 ( .A(n15155), .B(n17245), .Z(n17243) );
  XNOR U17445 ( .A(key[634]), .B(n15158), .Z(n17245) );
  ANDN U17446 ( .B(n17246), .A(n16761), .Z(n17241) );
  XOR U17447 ( .A(n17247), .B(n17248), .Z(n16789) );
  XNOR U17448 ( .A(n17249), .B(n17250), .Z(n17248) );
  XOR U17449 ( .A(n17218), .B(n17234), .Z(n17247) );
  XOR U17450 ( .A(n17251), .B(n17252), .Z(n17234) );
  XNOR U17451 ( .A(n17238), .B(n17253), .Z(n17252) );
  XNOR U17452 ( .A(n16191), .B(n16189), .Z(n17253) );
  XNOR U17453 ( .A(n17254), .B(n16175), .Z(n16189) );
  XOR U17454 ( .A(n17255), .B(n17256), .Z(n17238) );
  XOR U17455 ( .A(n16185), .B(n16195), .Z(n17256) );
  XOR U17456 ( .A(n15135), .B(n17257), .Z(n17255) );
  XOR U17457 ( .A(key[633]), .B(n15185), .Z(n17257) );
  XOR U17458 ( .A(n17258), .B(n17259), .Z(n17251) );
  XNOR U17459 ( .A(key[635]), .B(n15139), .Z(n17259) );
  XOR U17460 ( .A(n17246), .B(n17217), .Z(n17180) );
  IV U17461 ( .A(n17166), .Z(n17217) );
  XOR U17462 ( .A(n17236), .B(n17260), .Z(n17166) );
  XOR U17463 ( .A(n17235), .B(n17250), .Z(n17260) );
  XNOR U17464 ( .A(n17261), .B(n17262), .Z(n17250) );
  XOR U17465 ( .A(n16219), .B(n16204), .Z(n17262) );
  XNOR U17466 ( .A(n17263), .B(n15164), .Z(n16204) );
  XOR U17467 ( .A(key[639]), .B(n15181), .Z(n17261) );
  XNOR U17468 ( .A(n17254), .B(n17264), .Z(n15181) );
  IV U17469 ( .A(n17147), .Z(n17246) );
  XOR U17470 ( .A(n17236), .B(n17265), .Z(n17147) );
  XOR U17471 ( .A(n17235), .B(n17249), .Z(n17265) );
  XNOR U17472 ( .A(n17266), .B(n16174), .Z(n17249) );
  XNOR U17473 ( .A(n17267), .B(n17268), .Z(n16174) );
  XNOR U17474 ( .A(n17254), .B(n16207), .Z(n17267) );
  XNOR U17475 ( .A(n17270), .B(n17271), .Z(n17266) );
  XOR U17476 ( .A(key[636]), .B(n16199), .Z(n17271) );
  IV U17477 ( .A(n17272), .Z(n16199) );
  XOR U17478 ( .A(n17273), .B(n17274), .Z(n17235) );
  XOR U17479 ( .A(n16212), .B(n16761), .Z(n17274) );
  IV U17480 ( .A(n17218), .Z(n16761) );
  XOR U17481 ( .A(n17275), .B(n17276), .Z(n17218) );
  XNOR U17482 ( .A(n15152), .B(n15162), .Z(n17276) );
  XOR U17483 ( .A(n16196), .B(n17277), .Z(n17275) );
  XOR U17484 ( .A(key[632]), .B(n17264), .Z(n17277) );
  XNOR U17485 ( .A(n17278), .B(n16203), .Z(n16212) );
  XOR U17486 ( .A(n17254), .B(n17279), .Z(n16203) );
  XNOR U17487 ( .A(n17280), .B(n17281), .Z(n17273) );
  XOR U17488 ( .A(key[638]), .B(n15192), .Z(n17281) );
  IV U17489 ( .A(n17239), .Z(n17236) );
  XOR U17490 ( .A(n17282), .B(n17283), .Z(n17239) );
  XOR U17491 ( .A(n16177), .B(n16208), .Z(n17283) );
  XOR U17492 ( .A(n16217), .B(n17285), .Z(n17282) );
  XNOR U17493 ( .A(key[637]), .B(n15177), .Z(n17285) );
  IV U17494 ( .A(n13960), .Z(n13561) );
  XOR U17495 ( .A(n16665), .B(n16738), .Z(n13960) );
  XOR U17496 ( .A(n16744), .B(n17286), .Z(n16738) );
  XOR U17497 ( .A(n17287), .B(n16697), .Z(n17286) );
  OR U17498 ( .A(n17288), .B(n16830), .Z(n16697) );
  XNOR U17499 ( .A(n16699), .B(n16825), .Z(n16830) );
  NOR U17500 ( .A(n17289), .B(n16825), .Z(n17287) );
  IV U17501 ( .A(n16782), .Z(n16665) );
  XNOR U17502 ( .A(n16744), .B(n17290), .Z(n16782) );
  XNOR U17503 ( .A(n16741), .B(n17291), .Z(n17290) );
  NAND U17504 ( .A(n17292), .B(n16705), .Z(n17291) );
  XNOR U17505 ( .A(n16743), .B(n16705), .Z(n16819) );
  XOR U17506 ( .A(n17294), .B(n16746), .Z(n16744) );
  OR U17507 ( .A(n16837), .B(n17295), .Z(n16746) );
  XNOR U17508 ( .A(n16839), .B(n16748), .Z(n16837) );
  XNOR U17509 ( .A(n16825), .B(n16705), .Z(n16748) );
  XOR U17510 ( .A(n17296), .B(n17297), .Z(n16705) );
  NANDN U17511 ( .A(n17298), .B(n17299), .Z(n17297) );
  XNOR U17512 ( .A(n17300), .B(n17301), .Z(n16825) );
  OR U17513 ( .A(n17298), .B(n17302), .Z(n17301) );
  ANDN U17514 ( .B(n16839), .A(n17303), .Z(n17294) );
  XOR U17515 ( .A(n16699), .B(n16743), .Z(n16839) );
  XOR U17516 ( .A(n17304), .B(n17296), .Z(n16743) );
  NANDN U17517 ( .A(n17305), .B(n17306), .Z(n17296) );
  ANDN U17518 ( .B(n17307), .A(n17308), .Z(n17304) );
  NANDN U17519 ( .A(n17305), .B(n17310), .Z(n17300) );
  XOR U17520 ( .A(n17311), .B(n17298), .Z(n17305) );
  XNOR U17521 ( .A(n17312), .B(n17313), .Z(n17298) );
  XOR U17522 ( .A(n17314), .B(n17307), .Z(n17313) );
  XNOR U17523 ( .A(n17315), .B(n17316), .Z(n17312) );
  XNOR U17524 ( .A(n17317), .B(n17318), .Z(n17316) );
  ANDN U17525 ( .B(n17307), .A(n17319), .Z(n17317) );
  IV U17526 ( .A(n17320), .Z(n17307) );
  ANDN U17527 ( .B(n17311), .A(n17319), .Z(n17309) );
  IV U17528 ( .A(n17315), .Z(n17319) );
  IV U17529 ( .A(n17308), .Z(n17311) );
  XNOR U17530 ( .A(n17314), .B(n17321), .Z(n17308) );
  XOR U17531 ( .A(n17322), .B(n17318), .Z(n17321) );
  NAND U17532 ( .A(n17310), .B(n17306), .Z(n17318) );
  XNOR U17533 ( .A(n17299), .B(n17320), .Z(n17306) );
  XOR U17534 ( .A(n17323), .B(n17324), .Z(n17320) );
  XOR U17535 ( .A(n17325), .B(n17326), .Z(n17324) );
  XNOR U17536 ( .A(n16826), .B(n17327), .Z(n17326) );
  XNOR U17537 ( .A(n17328), .B(n17329), .Z(n17323) );
  XNOR U17538 ( .A(n17330), .B(n17331), .Z(n17329) );
  ANDN U17539 ( .B(n16829), .A(n16700), .Z(n17330) );
  XNOR U17540 ( .A(n17315), .B(n17302), .Z(n17310) );
  XOR U17541 ( .A(n17332), .B(n17333), .Z(n17315) );
  XNOR U17542 ( .A(n17334), .B(n17327), .Z(n17333) );
  XOR U17543 ( .A(n17335), .B(n17336), .Z(n17327) );
  XNOR U17544 ( .A(n17337), .B(n17338), .Z(n17336) );
  NAND U17545 ( .A(n16749), .B(n16835), .Z(n17338) );
  XNOR U17546 ( .A(n17339), .B(n17340), .Z(n17332) );
  ANDN U17547 ( .B(n17341), .A(n16742), .Z(n17339) );
  ANDN U17548 ( .B(n17299), .A(n17302), .Z(n17322) );
  XOR U17549 ( .A(n17302), .B(n17299), .Z(n17314) );
  XNOR U17550 ( .A(n17342), .B(n17343), .Z(n17299) );
  XNOR U17551 ( .A(n17335), .B(n17344), .Z(n17343) );
  XNOR U17552 ( .A(n17334), .B(n16829), .Z(n17344) );
  XNOR U17553 ( .A(n17345), .B(n17346), .Z(n17342) );
  XNOR U17554 ( .A(n17347), .B(n17331), .Z(n17346) );
  OR U17555 ( .A(n16831), .B(n17288), .Z(n17331) );
  XNOR U17556 ( .A(n17345), .B(n17328), .Z(n17288) );
  XNOR U17557 ( .A(n16829), .B(n16826), .Z(n16831) );
  ANDN U17558 ( .B(n16826), .A(n17289), .Z(n17347) );
  XOR U17559 ( .A(n17348), .B(n17349), .Z(n17302) );
  XOR U17560 ( .A(n17335), .B(n17325), .Z(n17349) );
  XOR U17561 ( .A(n17292), .B(n16706), .Z(n17325) );
  XOR U17562 ( .A(n17350), .B(n17337), .Z(n17335) );
  NANDN U17563 ( .A(n17295), .B(n16838), .Z(n17337) );
  XOR U17564 ( .A(n16840), .B(n16835), .Z(n16838) );
  XNOR U17565 ( .A(n17341), .B(n17351), .Z(n16826) );
  XNOR U17566 ( .A(n17352), .B(n17353), .Z(n17351) );
  XOR U17567 ( .A(n17303), .B(n16749), .Z(n17295) );
  XNOR U17568 ( .A(n17289), .B(n17292), .Z(n16749) );
  IV U17569 ( .A(n17328), .Z(n17289) );
  XOR U17570 ( .A(n17354), .B(n17355), .Z(n17328) );
  XOR U17571 ( .A(n17356), .B(n17357), .Z(n17355) );
  XOR U17572 ( .A(n17345), .B(n17358), .Z(n17354) );
  ANDN U17573 ( .B(n16840), .A(n17303), .Z(n17350) );
  XNOR U17574 ( .A(n17345), .B(n17359), .Z(n17303) );
  XOR U17575 ( .A(n17341), .B(n16829), .Z(n16840) );
  XNOR U17576 ( .A(n17360), .B(n17361), .Z(n16829) );
  XOR U17577 ( .A(n17362), .B(n17357), .Z(n17361) );
  XNOR U17578 ( .A(n17363), .B(n17364), .Z(n17357) );
  XNOR U17579 ( .A(n17365), .B(n16362), .Z(n17364) );
  XOR U17580 ( .A(n17366), .B(n16392), .Z(n16362) );
  XNOR U17581 ( .A(n17367), .B(n17368), .Z(n17363) );
  XNOR U17582 ( .A(key[516]), .B(n16366), .Z(n17368) );
  IV U17583 ( .A(n16821), .Z(n17341) );
  XOR U17584 ( .A(n17334), .B(n17369), .Z(n17348) );
  XNOR U17585 ( .A(n17370), .B(n17340), .Z(n17369) );
  OR U17586 ( .A(n16820), .B(n17293), .Z(n17340) );
  XNOR U17587 ( .A(n17359), .B(n17292), .Z(n17293) );
  XNOR U17588 ( .A(n16821), .B(n16706), .Z(n16820) );
  ANDN U17589 ( .B(n17292), .A(n16706), .Z(n17370) );
  XOR U17590 ( .A(n17360), .B(n17371), .Z(n16706) );
  XOR U17591 ( .A(n17352), .B(n17372), .Z(n17371) );
  XOR U17592 ( .A(n17362), .B(n17360), .Z(n17292) );
  XNOR U17593 ( .A(n16742), .B(n16821), .Z(n17334) );
  XOR U17594 ( .A(n17360), .B(n17373), .Z(n16821) );
  XNOR U17595 ( .A(n17362), .B(n17356), .Z(n17373) );
  XOR U17596 ( .A(n17374), .B(n17375), .Z(n17356) );
  XNOR U17597 ( .A(n17376), .B(n17377), .Z(n17375) );
  XNOR U17598 ( .A(key[519]), .B(n16384), .Z(n17374) );
  XNOR U17599 ( .A(n17378), .B(n17379), .Z(n17360) );
  XOR U17600 ( .A(n16393), .B(n17380), .Z(n17379) );
  XNOR U17601 ( .A(key[517]), .B(n16387), .Z(n17378) );
  XNOR U17602 ( .A(n16394), .B(n17381), .Z(n16387) );
  IV U17603 ( .A(n17359), .Z(n16742) );
  XNOR U17604 ( .A(n17353), .B(n17382), .Z(n17359) );
  XOR U17605 ( .A(n17358), .B(n17372), .Z(n17382) );
  IV U17606 ( .A(n17362), .Z(n17372) );
  XOR U17607 ( .A(n17383), .B(n17384), .Z(n17362) );
  XOR U17608 ( .A(n16377), .B(n16700), .Z(n17384) );
  IV U17609 ( .A(n17345), .Z(n16700) );
  XOR U17610 ( .A(n17385), .B(n17386), .Z(n17345) );
  XOR U17611 ( .A(n15619), .B(n16381), .Z(n17386) );
  XOR U17612 ( .A(n17387), .B(n17388), .Z(n15619) );
  XOR U17613 ( .A(key[512]), .B(n16352), .Z(n17385) );
  XOR U17614 ( .A(n17366), .B(n16373), .Z(n16377) );
  XOR U17615 ( .A(n17389), .B(n17390), .Z(n17383) );
  XNOR U17616 ( .A(key[518]), .B(n17381), .Z(n17390) );
  XOR U17617 ( .A(n17391), .B(n17392), .Z(n17358) );
  XNOR U17618 ( .A(n17352), .B(n17393), .Z(n17392) );
  XNOR U17619 ( .A(n17394), .B(n16343), .Z(n17393) );
  XOR U17620 ( .A(n17366), .B(n16365), .Z(n16343) );
  XOR U17621 ( .A(n17395), .B(n17396), .Z(n17352) );
  XOR U17622 ( .A(n17388), .B(n15582), .Z(n17396) );
  XNOR U17623 ( .A(n16348), .B(n17397), .Z(n15582) );
  XOR U17624 ( .A(key[513]), .B(n15628), .Z(n17395) );
  XOR U17625 ( .A(n15583), .B(n17398), .Z(n17391) );
  XNOR U17626 ( .A(key[515]), .B(n17399), .Z(n17398) );
  XOR U17627 ( .A(n17400), .B(n17401), .Z(n17353) );
  XNOR U17628 ( .A(n15620), .B(n17397), .Z(n17401) );
  XOR U17629 ( .A(key[514]), .B(n15624), .Z(n17400) );
  XOR U17630 ( .A(n16358), .B(n17399), .Z(n15624) );
  IV U17631 ( .A(n17402), .Z(n16358) );
  XOR U17632 ( .A(n9612), .B(n10484), .Z(n9605) );
  XOR U17633 ( .A(n17403), .B(n17404), .Z(n10484) );
  XNOR U17634 ( .A(n14639), .B(n14522), .Z(n17404) );
  XNOR U17635 ( .A(n17405), .B(n17406), .Z(n14522) );
  XNOR U17636 ( .A(n17407), .B(n17408), .Z(n17406) );
  NANDN U17637 ( .A(n17409), .B(n17410), .Z(n17408) );
  XOR U17638 ( .A(n17411), .B(n17412), .Z(n14639) );
  XNOR U17639 ( .A(n17413), .B(n17414), .Z(n17412) );
  NANDN U17640 ( .A(n17415), .B(n14527), .Z(n17414) );
  XOR U17641 ( .A(n14647), .B(n14589), .Z(n17403) );
  XOR U17642 ( .A(n14619), .B(n14648), .Z(n14589) );
  XOR U17643 ( .A(n14521), .B(n17416), .Z(n14648) );
  XNOR U17644 ( .A(n17417), .B(n17418), .Z(n17416) );
  NANDN U17645 ( .A(n17419), .B(n17420), .Z(n17418) );
  XNOR U17646 ( .A(n17417), .B(n17422), .Z(n17421) );
  NANDN U17647 ( .A(n17423), .B(n17410), .Z(n17422) );
  OR U17648 ( .A(n17424), .B(n17425), .Z(n17417) );
  XNOR U17649 ( .A(n14521), .B(n17426), .Z(n14640) );
  XNOR U17650 ( .A(n17427), .B(n17428), .Z(n17426) );
  NANDN U17651 ( .A(n17429), .B(n17430), .Z(n17428) );
  XOR U17652 ( .A(n17431), .B(n17427), .Z(n14521) );
  NANDN U17653 ( .A(n17432), .B(n17433), .Z(n17427) );
  ANDN U17654 ( .B(n17434), .A(n17435), .Z(n17431) );
  XOR U17655 ( .A(n17437), .B(n17407), .Z(n17436) );
  OR U17656 ( .A(n17424), .B(n17438), .Z(n17407) );
  XNOR U17657 ( .A(n17410), .B(n17420), .Z(n17424) );
  ANDN U17658 ( .B(n17420), .A(n17439), .Z(n17437) );
  XNOR U17659 ( .A(n17405), .B(n17440), .Z(n14523) );
  XOR U17660 ( .A(n17441), .B(n17413), .Z(n17440) );
  XOR U17661 ( .A(n14645), .B(n14527), .Z(n14643) );
  XOR U17662 ( .A(n17411), .B(n17444), .Z(n17405) );
  XNOR U17663 ( .A(n17445), .B(n17446), .Z(n17444) );
  NANDN U17664 ( .A(n17429), .B(n17447), .Z(n17446) );
  XNOR U17665 ( .A(n17448), .B(n17445), .Z(n17411) );
  OR U17666 ( .A(n17432), .B(n17449), .Z(n17445) );
  XNOR U17667 ( .A(n17435), .B(n17429), .Z(n17432) );
  XNOR U17668 ( .A(n17420), .B(n14527), .Z(n17429) );
  XOR U17669 ( .A(n17450), .B(n17451), .Z(n14527) );
  NANDN U17670 ( .A(n17452), .B(n17453), .Z(n17451) );
  XOR U17671 ( .A(n17454), .B(n17455), .Z(n17420) );
  NANDN U17672 ( .A(n17452), .B(n17456), .Z(n17455) );
  NOR U17673 ( .A(n17435), .B(n17457), .Z(n17448) );
  XNOR U17674 ( .A(n14645), .B(n17410), .Z(n17435) );
  XNOR U17675 ( .A(n17458), .B(n17454), .Z(n17410) );
  NANDN U17676 ( .A(n17459), .B(n17460), .Z(n17454) );
  XOR U17677 ( .A(n17456), .B(n17461), .Z(n17460) );
  ANDN U17678 ( .B(n17461), .A(n17462), .Z(n17458) );
  XNOR U17679 ( .A(n17463), .B(n17450), .Z(n14645) );
  NANDN U17680 ( .A(n17459), .B(n17464), .Z(n17450) );
  XOR U17681 ( .A(n17465), .B(n17453), .Z(n17464) );
  XNOR U17682 ( .A(n17466), .B(n17467), .Z(n17452) );
  XOR U17683 ( .A(n17468), .B(n17469), .Z(n17467) );
  XNOR U17684 ( .A(n17470), .B(n17471), .Z(n17466) );
  XNOR U17685 ( .A(n17472), .B(n17473), .Z(n17471) );
  ANDN U17686 ( .B(n17465), .A(n17469), .Z(n17472) );
  ANDN U17687 ( .B(n17465), .A(n17462), .Z(n17463) );
  XNOR U17688 ( .A(n17468), .B(n17474), .Z(n17462) );
  XOR U17689 ( .A(n17475), .B(n17473), .Z(n17474) );
  NAND U17690 ( .A(n17476), .B(n17477), .Z(n17473) );
  XNOR U17691 ( .A(n17470), .B(n17453), .Z(n17477) );
  IV U17692 ( .A(n17465), .Z(n17470) );
  XNOR U17693 ( .A(n17456), .B(n17469), .Z(n17476) );
  IV U17694 ( .A(n17461), .Z(n17469) );
  XOR U17695 ( .A(n17478), .B(n17479), .Z(n17461) );
  XNOR U17696 ( .A(n17480), .B(n17481), .Z(n17479) );
  XNOR U17697 ( .A(n17482), .B(n17483), .Z(n17478) );
  NOR U17698 ( .A(n14646), .B(n17443), .Z(n17482) );
  AND U17699 ( .A(n17453), .B(n17456), .Z(n17475) );
  XNOR U17700 ( .A(n17453), .B(n17456), .Z(n17468) );
  XNOR U17701 ( .A(n17484), .B(n17485), .Z(n17456) );
  XNOR U17702 ( .A(n17486), .B(n17481), .Z(n17485) );
  XOR U17703 ( .A(n17487), .B(n17488), .Z(n17484) );
  XNOR U17704 ( .A(n17489), .B(n17483), .Z(n17488) );
  OR U17705 ( .A(n14644), .B(n17442), .Z(n17483) );
  XNOR U17706 ( .A(n17443), .B(n17415), .Z(n17442) );
  XNOR U17707 ( .A(n14646), .B(n14528), .Z(n14644) );
  ANDN U17708 ( .B(n17490), .A(n17415), .Z(n17489) );
  XNOR U17709 ( .A(n17491), .B(n17492), .Z(n17453) );
  XNOR U17710 ( .A(n17481), .B(n17493), .Z(n17492) );
  XOR U17711 ( .A(n17423), .B(n17487), .Z(n17493) );
  XNOR U17712 ( .A(n17443), .B(n17494), .Z(n17481) );
  XOR U17713 ( .A(n17409), .B(n17495), .Z(n17491) );
  XNOR U17714 ( .A(n17496), .B(n17497), .Z(n17495) );
  ANDN U17715 ( .B(n17498), .A(n17439), .Z(n17496) );
  XNOR U17716 ( .A(n17499), .B(n17500), .Z(n17465) );
  XNOR U17717 ( .A(n17486), .B(n17501), .Z(n17500) );
  XNOR U17718 ( .A(n17419), .B(n17480), .Z(n17501) );
  XOR U17719 ( .A(n17487), .B(n17502), .Z(n17480) );
  XNOR U17720 ( .A(n17503), .B(n17504), .Z(n17502) );
  NAND U17721 ( .A(n17447), .B(n17430), .Z(n17504) );
  XNOR U17722 ( .A(n17505), .B(n17503), .Z(n17487) );
  NANDN U17723 ( .A(n17449), .B(n17433), .Z(n17503) );
  XOR U17724 ( .A(n17434), .B(n17430), .Z(n17433) );
  XNOR U17725 ( .A(n17498), .B(n14528), .Z(n17430) );
  XOR U17726 ( .A(n17457), .B(n17447), .Z(n17449) );
  XNOR U17727 ( .A(n17439), .B(n17506), .Z(n17447) );
  ANDN U17728 ( .B(n17434), .A(n17457), .Z(n17505) );
  XNOR U17729 ( .A(n17409), .B(n17443), .Z(n17457) );
  XOR U17730 ( .A(n17507), .B(n17508), .Z(n17443) );
  XNOR U17731 ( .A(n17509), .B(n17510), .Z(n17508) );
  XOR U17732 ( .A(n17506), .B(n17490), .Z(n17486) );
  IV U17733 ( .A(n14528), .Z(n17490) );
  XOR U17734 ( .A(n17511), .B(n17512), .Z(n14528) );
  XOR U17735 ( .A(n17513), .B(n17510), .Z(n17512) );
  IV U17736 ( .A(n17415), .Z(n17506) );
  XOR U17737 ( .A(n17510), .B(n17514), .Z(n17415) );
  XNOR U17738 ( .A(n17515), .B(n17516), .Z(n17499) );
  XNOR U17739 ( .A(n17517), .B(n17497), .Z(n17516) );
  OR U17740 ( .A(n17425), .B(n17438), .Z(n17497) );
  XNOR U17741 ( .A(n17409), .B(n17439), .Z(n17438) );
  IV U17742 ( .A(n17515), .Z(n17439) );
  XOR U17743 ( .A(n17423), .B(n17498), .Z(n17425) );
  IV U17744 ( .A(n17419), .Z(n17498) );
  XOR U17745 ( .A(n17494), .B(n17518), .Z(n17419) );
  XNOR U17746 ( .A(n17519), .B(n17507), .Z(n17518) );
  XOR U17747 ( .A(n17520), .B(n17521), .Z(n17507) );
  XOR U17748 ( .A(n12291), .B(n14423), .Z(n17521) );
  XOR U17749 ( .A(n12296), .B(n14410), .Z(n12291) );
  XOR U17750 ( .A(n17522), .B(n17523), .Z(n12296) );
  XOR U17751 ( .A(n17524), .B(n17525), .Z(n17523) );
  XNOR U17752 ( .A(n17526), .B(n17527), .Z(n17522) );
  XOR U17753 ( .A(n12288), .B(n12298), .Z(n13382) );
  IV U17754 ( .A(n14646), .Z(n17494) );
  XOR U17755 ( .A(n17511), .B(n17528), .Z(n14646) );
  XOR U17756 ( .A(n17510), .B(n17529), .Z(n17528) );
  NOR U17757 ( .A(n17423), .B(n17409), .Z(n17517) );
  XOR U17758 ( .A(n17511), .B(n17530), .Z(n17423) );
  XOR U17759 ( .A(n17510), .B(n17531), .Z(n17530) );
  XOR U17760 ( .A(n17532), .B(n17533), .Z(n17510) );
  XNOR U17761 ( .A(n17409), .B(n14414), .Z(n17533) );
  XNOR U17762 ( .A(n13416), .B(n17534), .Z(n14414) );
  XOR U17763 ( .A(n12277), .B(n14400), .Z(n13416) );
  IV U17764 ( .A(n12304), .Z(n14400) );
  XNOR U17765 ( .A(n17535), .B(n17536), .Z(n12304) );
  XOR U17766 ( .A(n17537), .B(n17538), .Z(n12277) );
  XNOR U17767 ( .A(n12303), .B(n17539), .Z(n17532) );
  XNOR U17768 ( .A(key[646]), .B(n17540), .Z(n17539) );
  XOR U17769 ( .A(n12311), .B(n13391), .Z(n12303) );
  XOR U17770 ( .A(n17541), .B(n17542), .Z(n13391) );
  XNOR U17771 ( .A(n17524), .B(n17543), .Z(n17542) );
  XNOR U17772 ( .A(n17526), .B(n17544), .Z(n17541) );
  IV U17773 ( .A(n17514), .Z(n17511) );
  XOR U17774 ( .A(n17545), .B(n17546), .Z(n17514) );
  XOR U17775 ( .A(n13418), .B(n14401), .Z(n17546) );
  XNOR U17776 ( .A(n13403), .B(n12273), .Z(n14401) );
  XNOR U17777 ( .A(n17547), .B(n17548), .Z(n12273) );
  XOR U17778 ( .A(n17549), .B(n17550), .Z(n17548) );
  XNOR U17779 ( .A(n17551), .B(n17552), .Z(n17547) );
  XOR U17780 ( .A(n17553), .B(n17554), .Z(n17552) );
  ANDN U17781 ( .B(n17555), .A(n17556), .Z(n17554) );
  XOR U17782 ( .A(n17557), .B(n17558), .Z(n13403) );
  XNOR U17783 ( .A(n17559), .B(n17560), .Z(n17558) );
  XNOR U17784 ( .A(n17561), .B(n17562), .Z(n17557) );
  XOR U17785 ( .A(n17563), .B(n17564), .Z(n17562) );
  ANDN U17786 ( .B(n17565), .A(n17566), .Z(n17564) );
  XNOR U17787 ( .A(key[645]), .B(n13407), .Z(n17545) );
  XOR U17788 ( .A(n12275), .B(n14403), .Z(n13407) );
  IV U17789 ( .A(n17540), .Z(n14403) );
  XOR U17790 ( .A(n17567), .B(n17568), .Z(n17540) );
  XOR U17791 ( .A(n17544), .B(n17525), .Z(n12275) );
  XNOR U17792 ( .A(n17569), .B(n17570), .Z(n17525) );
  XOR U17793 ( .A(n17571), .B(n17572), .Z(n17570) );
  NOR U17794 ( .A(n17573), .B(n17574), .Z(n17571) );
  XOR U17795 ( .A(n17575), .B(n17576), .Z(n17515) );
  XNOR U17796 ( .A(n17531), .B(n17529), .Z(n17576) );
  XNOR U17797 ( .A(n17577), .B(n17578), .Z(n17529) );
  XOR U17798 ( .A(n17534), .B(n14406), .Z(n17578) );
  XNOR U17799 ( .A(n17579), .B(n17580), .Z(n13408) );
  XOR U17800 ( .A(n17537), .B(n17560), .Z(n17580) );
  XNOR U17801 ( .A(n17581), .B(n17582), .Z(n17560) );
  XNOR U17802 ( .A(n17583), .B(n17584), .Z(n17582) );
  OR U17803 ( .A(n17585), .B(n17586), .Z(n17584) );
  XOR U17804 ( .A(n17587), .B(n17588), .Z(n17579) );
  XOR U17805 ( .A(n17589), .B(n17590), .Z(n12268) );
  XNOR U17806 ( .A(n17535), .B(n17550), .Z(n17590) );
  XNOR U17807 ( .A(n17591), .B(n17592), .Z(n17550) );
  XNOR U17808 ( .A(n17593), .B(n17594), .Z(n17592) );
  OR U17809 ( .A(n17595), .B(n17596), .Z(n17594) );
  XOR U17810 ( .A(n17597), .B(n17598), .Z(n17589) );
  XNOR U17811 ( .A(n17599), .B(n13392), .Z(n17534) );
  XNOR U17812 ( .A(n17600), .B(n17601), .Z(n13392) );
  XNOR U17813 ( .A(n17602), .B(n17603), .Z(n17601) );
  XOR U17814 ( .A(n17604), .B(n17567), .Z(n17600) );
  XNOR U17815 ( .A(n17605), .B(n14391), .Z(n17531) );
  XOR U17816 ( .A(n17606), .B(n17607), .Z(n14391) );
  XNOR U17817 ( .A(n13386), .B(n12259), .Z(n17607) );
  XNOR U17818 ( .A(n12298), .B(n17549), .Z(n12259) );
  XNOR U17819 ( .A(n17608), .B(n17609), .Z(n12298) );
  XNOR U17820 ( .A(n17559), .B(n12288), .Z(n13386) );
  XOR U17821 ( .A(n17610), .B(n17611), .Z(n12288) );
  XNOR U17822 ( .A(n17599), .B(n13418), .Z(n17606) );
  XOR U17823 ( .A(n17612), .B(n17613), .Z(n13418) );
  XNOR U17824 ( .A(n17614), .B(n17603), .Z(n17613) );
  XNOR U17825 ( .A(n17615), .B(n17616), .Z(n17603) );
  XNOR U17826 ( .A(n17617), .B(n17618), .Z(n17616) );
  NANDN U17827 ( .A(n17619), .B(n17620), .Z(n17618) );
  XNOR U17828 ( .A(n17621), .B(n17622), .Z(n17612) );
  XOR U17829 ( .A(n17623), .B(n17624), .Z(n17622) );
  ANDN U17830 ( .B(n17625), .A(n17626), .Z(n17624) );
  XNOR U17831 ( .A(n12258), .B(n17627), .Z(n17605) );
  XNOR U17832 ( .A(key[644]), .B(n13401), .Z(n17627) );
  XOR U17833 ( .A(n12311), .B(n13417), .Z(n12258) );
  XOR U17834 ( .A(n17628), .B(n17629), .Z(n13417) );
  XNOR U17835 ( .A(n17630), .B(n17543), .Z(n17629) );
  XNOR U17836 ( .A(n17631), .B(n17632), .Z(n17543) );
  XNOR U17837 ( .A(n17633), .B(n17634), .Z(n17632) );
  NANDN U17838 ( .A(n17635), .B(n17636), .Z(n17634) );
  XNOR U17839 ( .A(n17637), .B(n17638), .Z(n17628) );
  XNOR U17840 ( .A(n17572), .B(n17639), .Z(n17638) );
  ANDN U17841 ( .B(n17640), .A(n17641), .Z(n17639) );
  NANDN U17842 ( .A(n17642), .B(n17643), .Z(n17572) );
  XNOR U17843 ( .A(n17409), .B(n17509), .Z(n17575) );
  XOR U17844 ( .A(n17644), .B(n17645), .Z(n17509) );
  XNOR U17845 ( .A(n14419), .B(n17646), .Z(n17645) );
  XNOR U17846 ( .A(n12281), .B(n17519), .Z(n17646) );
  IV U17847 ( .A(n17513), .Z(n17519) );
  XNOR U17848 ( .A(n17647), .B(n17648), .Z(n17513) );
  XOR U17849 ( .A(n17649), .B(n12297), .Z(n17648) );
  XOR U17850 ( .A(n17650), .B(n14423), .Z(n12297) );
  XNOR U17851 ( .A(key[641]), .B(n13412), .Z(n17647) );
  XNOR U17852 ( .A(n13383), .B(n14430), .Z(n13412) );
  IV U17853 ( .A(n12290), .Z(n14430) );
  XNOR U17854 ( .A(n17535), .B(n17651), .Z(n12290) );
  XOR U17855 ( .A(n17608), .B(n17598), .Z(n17651) );
  XNOR U17856 ( .A(n17652), .B(n17609), .Z(n17535) );
  IV U17857 ( .A(n12313), .Z(n13383) );
  XOR U17858 ( .A(n17537), .B(n17653), .Z(n12313) );
  XOR U17859 ( .A(n17610), .B(n17588), .Z(n17653) );
  XOR U17860 ( .A(n17611), .B(n17654), .Z(n17537) );
  XOR U17861 ( .A(n12311), .B(n13400), .Z(n12281) );
  XNOR U17862 ( .A(n17637), .B(n12287), .Z(n13400) );
  IV U17863 ( .A(n17650), .Z(n12287) );
  XNOR U17864 ( .A(n17655), .B(n17524), .Z(n17650) );
  XOR U17865 ( .A(n17637), .B(n17656), .Z(n12311) );
  XNOR U17866 ( .A(n17631), .B(n17657), .Z(n17637) );
  XOR U17867 ( .A(n17658), .B(n17659), .Z(n17657) );
  ANDN U17868 ( .B(n17660), .A(n17574), .Z(n17658) );
  XNOR U17869 ( .A(n17661), .B(n17662), .Z(n17631) );
  XNOR U17870 ( .A(n17663), .B(n17664), .Z(n17662) );
  NAND U17871 ( .A(n17665), .B(n17666), .Z(n17664) );
  XNOR U17872 ( .A(n17599), .B(n13401), .Z(n14419) );
  XOR U17873 ( .A(n17621), .B(n14423), .Z(n13401) );
  XOR U17874 ( .A(n17667), .B(n17602), .Z(n14423) );
  IV U17875 ( .A(n13413), .Z(n17599) );
  XOR U17876 ( .A(n13371), .B(n17668), .Z(n17644) );
  XOR U17877 ( .A(key[643]), .B(n14410), .Z(n17668) );
  XNOR U17878 ( .A(n17669), .B(n17670), .Z(n14410) );
  XNOR U17879 ( .A(n17602), .B(n17568), .Z(n17670) );
  XNOR U17880 ( .A(n17671), .B(n17672), .Z(n17568) );
  XNOR U17881 ( .A(n17673), .B(n17623), .Z(n17672) );
  ANDN U17882 ( .B(n17674), .A(n17675), .Z(n17623) );
  NOR U17883 ( .A(n17676), .B(n17677), .Z(n17673) );
  XNOR U17884 ( .A(n17604), .B(n17678), .Z(n17669) );
  XNOR U17885 ( .A(n12300), .B(n12283), .Z(n13371) );
  XNOR U17886 ( .A(n17679), .B(n17680), .Z(n12283) );
  XNOR U17887 ( .A(n17652), .B(n17536), .Z(n17680) );
  XNOR U17888 ( .A(n17681), .B(n17682), .Z(n17536) );
  XNOR U17889 ( .A(n17683), .B(n17553), .Z(n17682) );
  ANDN U17890 ( .B(n17684), .A(n17685), .Z(n17553) );
  ANDN U17891 ( .B(n17686), .A(n17687), .Z(n17683) );
  XNOR U17892 ( .A(n17551), .B(n17688), .Z(n17652) );
  XNOR U17893 ( .A(n17689), .B(n17690), .Z(n17688) );
  NANDN U17894 ( .A(n17691), .B(n17692), .Z(n17690) );
  XNOR U17895 ( .A(n17608), .B(n17598), .Z(n17679) );
  XNOR U17896 ( .A(n17689), .B(n17694), .Z(n17693) );
  OR U17897 ( .A(n17595), .B(n17695), .Z(n17694) );
  OR U17898 ( .A(n17696), .B(n17697), .Z(n17689) );
  XNOR U17899 ( .A(n17551), .B(n17698), .Z(n17681) );
  XNOR U17900 ( .A(n17699), .B(n17700), .Z(n17698) );
  NANDN U17901 ( .A(n17701), .B(n17702), .Z(n17700) );
  XOR U17902 ( .A(n17703), .B(n17699), .Z(n17551) );
  NANDN U17903 ( .A(n17704), .B(n17705), .Z(n17699) );
  ANDN U17904 ( .B(n17706), .A(n17707), .Z(n17703) );
  IV U17905 ( .A(n17597), .Z(n17608) );
  XOR U17906 ( .A(n17708), .B(n17709), .Z(n17597) );
  XOR U17907 ( .A(n17710), .B(n17711), .Z(n17709) );
  NAND U17908 ( .A(n17712), .B(n17555), .Z(n17711) );
  XOR U17909 ( .A(n17713), .B(n17714), .Z(n12300) );
  XOR U17910 ( .A(n17654), .B(n17538), .Z(n17714) );
  XNOR U17911 ( .A(n17715), .B(n17716), .Z(n17538) );
  XNOR U17912 ( .A(n17717), .B(n17563), .Z(n17716) );
  ANDN U17913 ( .B(n17718), .A(n17719), .Z(n17563) );
  ANDN U17914 ( .B(n17720), .A(n17721), .Z(n17717) );
  XOR U17915 ( .A(n17561), .B(n17722), .Z(n17654) );
  XNOR U17916 ( .A(n17723), .B(n17724), .Z(n17722) );
  NANDN U17917 ( .A(n17725), .B(n17726), .Z(n17724) );
  XNOR U17918 ( .A(n17610), .B(n17588), .Z(n17713) );
  XNOR U17919 ( .A(n17723), .B(n17728), .Z(n17727) );
  OR U17920 ( .A(n17585), .B(n17729), .Z(n17728) );
  OR U17921 ( .A(n17730), .B(n17731), .Z(n17723) );
  XNOR U17922 ( .A(n17561), .B(n17732), .Z(n17715) );
  XNOR U17923 ( .A(n17733), .B(n17734), .Z(n17732) );
  NANDN U17924 ( .A(n17735), .B(n17736), .Z(n17734) );
  XOR U17925 ( .A(n17737), .B(n17733), .Z(n17561) );
  NANDN U17926 ( .A(n17738), .B(n17739), .Z(n17733) );
  ANDN U17927 ( .B(n17740), .A(n17741), .Z(n17737) );
  IV U17928 ( .A(n17587), .Z(n17610) );
  XOR U17929 ( .A(n17742), .B(n17743), .Z(n17587) );
  XOR U17930 ( .A(n17744), .B(n17745), .Z(n17743) );
  NAND U17931 ( .A(n17746), .B(n17565), .Z(n17745) );
  XNOR U17932 ( .A(n17747), .B(n17748), .Z(n17409) );
  XOR U17933 ( .A(n12286), .B(n12310), .Z(n17748) );
  XOR U17934 ( .A(n13413), .B(n14393), .Z(n12310) );
  XOR U17935 ( .A(n17591), .B(n17749), .Z(n17549) );
  XNOR U17936 ( .A(n17750), .B(n17710), .Z(n17749) );
  XOR U17937 ( .A(n17686), .B(n17555), .Z(n17684) );
  ANDN U17938 ( .B(n17686), .A(n17752), .Z(n17750) );
  XNOR U17939 ( .A(n17708), .B(n17753), .Z(n17591) );
  XNOR U17940 ( .A(n17754), .B(n17755), .Z(n17753) );
  NANDN U17941 ( .A(n17701), .B(n17756), .Z(n17755) );
  XNOR U17942 ( .A(n17708), .B(n17757), .Z(n17609) );
  XOR U17943 ( .A(n17758), .B(n17593), .Z(n17757) );
  OR U17944 ( .A(n17759), .B(n17696), .Z(n17593) );
  XNOR U17945 ( .A(n17595), .B(n17691), .Z(n17696) );
  NOR U17946 ( .A(n17760), .B(n17691), .Z(n17758) );
  XOR U17947 ( .A(n17761), .B(n17754), .Z(n17708) );
  OR U17948 ( .A(n17704), .B(n17762), .Z(n17754) );
  XOR U17949 ( .A(n17763), .B(n17701), .Z(n17704) );
  XOR U17950 ( .A(n17691), .B(n17555), .Z(n17701) );
  XOR U17951 ( .A(n17764), .B(n17765), .Z(n17555) );
  NANDN U17952 ( .A(n17766), .B(n17767), .Z(n17765) );
  XNOR U17953 ( .A(n17768), .B(n17769), .Z(n17691) );
  OR U17954 ( .A(n17766), .B(n17770), .Z(n17769) );
  ANDN U17955 ( .B(n17763), .A(n17771), .Z(n17761) );
  IV U17956 ( .A(n17707), .Z(n17763) );
  XOR U17957 ( .A(n17595), .B(n17686), .Z(n17707) );
  XNOR U17958 ( .A(n17772), .B(n17764), .Z(n17686) );
  NANDN U17959 ( .A(n17773), .B(n17774), .Z(n17764) );
  ANDN U17960 ( .B(n17775), .A(n17776), .Z(n17772) );
  NANDN U17961 ( .A(n17773), .B(n17778), .Z(n17768) );
  XOR U17962 ( .A(n17779), .B(n17766), .Z(n17773) );
  XNOR U17963 ( .A(n17780), .B(n17781), .Z(n17766) );
  XOR U17964 ( .A(n17782), .B(n17775), .Z(n17781) );
  XNOR U17965 ( .A(n17783), .B(n17784), .Z(n17780) );
  XNOR U17966 ( .A(n17785), .B(n17786), .Z(n17784) );
  ANDN U17967 ( .B(n17775), .A(n17787), .Z(n17785) );
  IV U17968 ( .A(n17788), .Z(n17775) );
  ANDN U17969 ( .B(n17779), .A(n17787), .Z(n17777) );
  IV U17970 ( .A(n17783), .Z(n17787) );
  IV U17971 ( .A(n17776), .Z(n17779) );
  XNOR U17972 ( .A(n17782), .B(n17789), .Z(n17776) );
  XOR U17973 ( .A(n17790), .B(n17786), .Z(n17789) );
  NAND U17974 ( .A(n17778), .B(n17774), .Z(n17786) );
  XNOR U17975 ( .A(n17767), .B(n17788), .Z(n17774) );
  XOR U17976 ( .A(n17791), .B(n17792), .Z(n17788) );
  XOR U17977 ( .A(n17793), .B(n17794), .Z(n17792) );
  XNOR U17978 ( .A(n17692), .B(n17795), .Z(n17794) );
  XNOR U17979 ( .A(n17796), .B(n17797), .Z(n17791) );
  XNOR U17980 ( .A(n17798), .B(n17799), .Z(n17797) );
  ANDN U17981 ( .B(n17800), .A(n17596), .Z(n17798) );
  XNOR U17982 ( .A(n17783), .B(n17770), .Z(n17778) );
  XOR U17983 ( .A(n17801), .B(n17802), .Z(n17783) );
  XNOR U17984 ( .A(n17803), .B(n17795), .Z(n17802) );
  XOR U17985 ( .A(n17804), .B(n17805), .Z(n17795) );
  XNOR U17986 ( .A(n17806), .B(n17807), .Z(n17805) );
  NAND U17987 ( .A(n17756), .B(n17702), .Z(n17807) );
  XNOR U17988 ( .A(n17808), .B(n17809), .Z(n17801) );
  ANDN U17989 ( .B(n17810), .A(n17752), .Z(n17808) );
  ANDN U17990 ( .B(n17767), .A(n17770), .Z(n17790) );
  XOR U17991 ( .A(n17770), .B(n17767), .Z(n17782) );
  XNOR U17992 ( .A(n17811), .B(n17812), .Z(n17767) );
  XNOR U17993 ( .A(n17804), .B(n17813), .Z(n17812) );
  XOR U17994 ( .A(n17803), .B(n17695), .Z(n17813) );
  XOR U17995 ( .A(n17596), .B(n17814), .Z(n17811) );
  XNOR U17996 ( .A(n17815), .B(n17799), .Z(n17814) );
  OR U17997 ( .A(n17697), .B(n17759), .Z(n17799) );
  XNOR U17998 ( .A(n17596), .B(n17760), .Z(n17759) );
  XOR U17999 ( .A(n17695), .B(n17692), .Z(n17697) );
  ANDN U18000 ( .B(n17692), .A(n17760), .Z(n17815) );
  XOR U18001 ( .A(n17816), .B(n17817), .Z(n17770) );
  XOR U18002 ( .A(n17804), .B(n17793), .Z(n17817) );
  XOR U18003 ( .A(n17712), .B(n17556), .Z(n17793) );
  XOR U18004 ( .A(n17818), .B(n17806), .Z(n17804) );
  NANDN U18005 ( .A(n17762), .B(n17705), .Z(n17806) );
  XOR U18006 ( .A(n17706), .B(n17702), .Z(n17705) );
  XNOR U18007 ( .A(n17810), .B(n17819), .Z(n17692) );
  XOR U18008 ( .A(n17820), .B(n17821), .Z(n17819) );
  XOR U18009 ( .A(n17771), .B(n17756), .Z(n17762) );
  XNOR U18010 ( .A(n17760), .B(n17712), .Z(n17756) );
  IV U18011 ( .A(n17796), .Z(n17760) );
  XOR U18012 ( .A(n17822), .B(n17823), .Z(n17796) );
  XOR U18013 ( .A(n17824), .B(n17825), .Z(n17823) );
  XNOR U18014 ( .A(n17596), .B(n17826), .Z(n17822) );
  ANDN U18015 ( .B(n17706), .A(n17771), .Z(n17818) );
  XNOR U18016 ( .A(n17596), .B(n17752), .Z(n17771) );
  XOR U18017 ( .A(n17810), .B(n17800), .Z(n17706) );
  IV U18018 ( .A(n17695), .Z(n17800) );
  XOR U18019 ( .A(n17827), .B(n17828), .Z(n17695) );
  XOR U18020 ( .A(n17829), .B(n17825), .Z(n17828) );
  XNOR U18021 ( .A(n17830), .B(n17831), .Z(n17825) );
  XNOR U18022 ( .A(n15169), .B(n17270), .Z(n17831) );
  XNOR U18023 ( .A(n17264), .B(n15190), .Z(n17270) );
  XNOR U18024 ( .A(n17832), .B(n17833), .Z(n15190) );
  XOR U18025 ( .A(n17834), .B(n17835), .Z(n17833) );
  XNOR U18026 ( .A(n17836), .B(n17837), .Z(n17832) );
  XOR U18027 ( .A(n17838), .B(n17839), .Z(n17837) );
  ANDN U18028 ( .B(n17840), .A(n17841), .Z(n17839) );
  XNOR U18029 ( .A(n17272), .B(n16175), .Z(n15169) );
  XOR U18030 ( .A(n17842), .B(n16185), .Z(n16175) );
  XOR U18031 ( .A(n17843), .B(n15155), .Z(n17272) );
  XNOR U18032 ( .A(n15168), .B(n17844), .Z(n17830) );
  XNOR U18033 ( .A(key[628]), .B(n17269), .Z(n17844) );
  XNOR U18034 ( .A(n16216), .B(n17284), .Z(n15168) );
  IV U18035 ( .A(n17687), .Z(n17810) );
  XOR U18036 ( .A(n17803), .B(n17845), .Z(n17816) );
  XNOR U18037 ( .A(n17846), .B(n17809), .Z(n17845) );
  OR U18038 ( .A(n17685), .B(n17751), .Z(n17809) );
  XNOR U18039 ( .A(n17847), .B(n17712), .Z(n17751) );
  XNOR U18040 ( .A(n17687), .B(n17556), .Z(n17685) );
  ANDN U18041 ( .B(n17712), .A(n17556), .Z(n17846) );
  XOR U18042 ( .A(n17827), .B(n17848), .Z(n17556) );
  XNOR U18043 ( .A(n17849), .B(n17829), .Z(n17848) );
  XOR U18044 ( .A(n17829), .B(n17827), .Z(n17712) );
  XNOR U18045 ( .A(n17752), .B(n17687), .Z(n17803) );
  XOR U18046 ( .A(n17827), .B(n17850), .Z(n17687) );
  XNOR U18047 ( .A(n17829), .B(n17824), .Z(n17850) );
  XOR U18048 ( .A(n17851), .B(n17852), .Z(n17824) );
  XNOR U18049 ( .A(n17853), .B(n15163), .Z(n17852) );
  XNOR U18050 ( .A(n17854), .B(n17855), .Z(n17279) );
  XOR U18051 ( .A(n17856), .B(n17857), .Z(n17855) );
  XOR U18052 ( .A(n17858), .B(n17859), .Z(n17854) );
  XNOR U18053 ( .A(n17860), .B(n17861), .Z(n16219) );
  XNOR U18054 ( .A(n17862), .B(n17863), .Z(n17861) );
  XOR U18055 ( .A(key[631]), .B(n17264), .Z(n17851) );
  XNOR U18056 ( .A(n17864), .B(n17865), .Z(n17827) );
  XNOR U18057 ( .A(n15189), .B(n17278), .Z(n17865) );
  XNOR U18058 ( .A(n15177), .B(n15188), .Z(n17278) );
  XOR U18059 ( .A(n17866), .B(n17867), .Z(n15177) );
  XOR U18060 ( .A(n17868), .B(n17869), .Z(n16207) );
  XNOR U18061 ( .A(n17870), .B(n17857), .Z(n17869) );
  XNOR U18062 ( .A(n17871), .B(n17872), .Z(n17857) );
  XNOR U18063 ( .A(n17873), .B(n17874), .Z(n17872) );
  NANDN U18064 ( .A(n17875), .B(n17876), .Z(n17874) );
  XNOR U18065 ( .A(n17842), .B(n17877), .Z(n17868) );
  XOR U18066 ( .A(n17878), .B(n17879), .Z(n17877) );
  ANDN U18067 ( .B(n17880), .A(n17881), .Z(n17879) );
  XNOR U18068 ( .A(n17882), .B(n17883), .Z(n16177) );
  XNOR U18069 ( .A(n17843), .B(n17863), .Z(n17883) );
  XNOR U18070 ( .A(n17884), .B(n17885), .Z(n17863) );
  XNOR U18071 ( .A(n17886), .B(n17887), .Z(n17885) );
  NANDN U18072 ( .A(n17888), .B(n17889), .Z(n17887) );
  XNOR U18073 ( .A(n17890), .B(n17891), .Z(n17882) );
  XOR U18074 ( .A(n17892), .B(n17893), .Z(n17891) );
  ANDN U18075 ( .B(n17894), .A(n17895), .Z(n17893) );
  XNOR U18076 ( .A(key[629]), .B(n17284), .Z(n17864) );
  XOR U18077 ( .A(n17896), .B(n17897), .Z(n17284) );
  XOR U18078 ( .A(n17898), .B(n17899), .Z(n17897) );
  XNOR U18079 ( .A(n17900), .B(n17901), .Z(n17896) );
  XOR U18080 ( .A(n17902), .B(n17903), .Z(n17901) );
  ANDN U18081 ( .B(n17904), .A(n17905), .Z(n17903) );
  IV U18082 ( .A(n17847), .Z(n17752) );
  XNOR U18083 ( .A(n17821), .B(n17906), .Z(n17847) );
  XOR U18084 ( .A(n17907), .B(n17908), .Z(n17829) );
  XOR U18085 ( .A(n17596), .B(n17280), .Z(n17908) );
  XNOR U18086 ( .A(n17264), .B(n15164), .Z(n17280) );
  XNOR U18087 ( .A(n17909), .B(n17910), .Z(n15164) );
  XOR U18088 ( .A(n17867), .B(n17835), .Z(n17910) );
  XNOR U18089 ( .A(n17911), .B(n17912), .Z(n17835) );
  XNOR U18090 ( .A(n17913), .B(n17914), .Z(n17912) );
  NANDN U18091 ( .A(n17915), .B(n17916), .Z(n17914) );
  XNOR U18092 ( .A(n17917), .B(n17918), .Z(n17596) );
  XNOR U18093 ( .A(n15182), .B(n15152), .Z(n16195) );
  XNOR U18094 ( .A(n17867), .B(n17919), .Z(n15152) );
  XNOR U18095 ( .A(n17920), .B(n17921), .Z(n17919) );
  XOR U18096 ( .A(n17922), .B(n17923), .Z(n17867) );
  IV U18097 ( .A(n17924), .Z(n15182) );
  XOR U18098 ( .A(n15183), .B(n16216), .Z(n15162) );
  XOR U18099 ( .A(n17925), .B(n17843), .Z(n15183) );
  XNOR U18100 ( .A(n17884), .B(n17926), .Z(n17843) );
  XNOR U18101 ( .A(n17927), .B(n17928), .Z(n17926) );
  ANDN U18102 ( .B(n17929), .A(n17930), .Z(n17927) );
  XNOR U18103 ( .A(n17931), .B(n17932), .Z(n17884) );
  XNOR U18104 ( .A(n17933), .B(n17934), .Z(n17932) );
  NANDN U18105 ( .A(n17935), .B(n17936), .Z(n17934) );
  XNOR U18106 ( .A(key[624]), .B(n17254), .Z(n17917) );
  XOR U18107 ( .A(n17842), .B(n17937), .Z(n17254) );
  XNOR U18108 ( .A(n17871), .B(n17938), .Z(n17842) );
  XOR U18109 ( .A(n17939), .B(n17940), .Z(n17938) );
  NOR U18110 ( .A(n17941), .B(n17942), .Z(n17939) );
  XOR U18111 ( .A(n17943), .B(n17944), .Z(n17871) );
  XNOR U18112 ( .A(n17945), .B(n17946), .Z(n17944) );
  NAND U18113 ( .A(n17947), .B(n17948), .Z(n17946) );
  XNOR U18114 ( .A(n15188), .B(n17949), .Z(n17907) );
  XNOR U18115 ( .A(key[630]), .B(n15176), .Z(n17949) );
  XNOR U18116 ( .A(n16209), .B(n17853), .Z(n15176) );
  XNOR U18117 ( .A(n17950), .B(n17951), .Z(n17263) );
  XNOR U18118 ( .A(n17952), .B(n17899), .Z(n17951) );
  XNOR U18119 ( .A(n17953), .B(n17954), .Z(n17899) );
  XNOR U18120 ( .A(n17955), .B(n17956), .Z(n17954) );
  NANDN U18121 ( .A(n17957), .B(n17958), .Z(n17956) );
  XOR U18122 ( .A(n16217), .B(n15192), .Z(n16209) );
  XOR U18123 ( .A(n17862), .B(n17959), .Z(n15192) );
  XOR U18124 ( .A(n17858), .B(n17960), .Z(n16217) );
  XNOR U18125 ( .A(n17952), .B(n17961), .Z(n15188) );
  XOR U18126 ( .A(n17962), .B(n17963), .Z(n17826) );
  XOR U18127 ( .A(n17258), .B(n17964), .Z(n17963) );
  XNOR U18128 ( .A(n15137), .B(n17849), .Z(n17964) );
  IV U18129 ( .A(n17820), .Z(n17849) );
  XNOR U18130 ( .A(n17965), .B(n17966), .Z(n17820) );
  XOR U18131 ( .A(n15151), .B(n16186), .Z(n17966) );
  XOR U18132 ( .A(n15153), .B(n15135), .Z(n16186) );
  IV U18133 ( .A(n16215), .Z(n15151) );
  XNOR U18134 ( .A(n15185), .B(n16196), .Z(n16215) );
  XNOR U18135 ( .A(n17856), .B(n17967), .Z(n16196) );
  XOR U18136 ( .A(n17858), .B(n17968), .Z(n17967) );
  XOR U18137 ( .A(n17862), .B(n17970), .Z(n15185) );
  XOR U18138 ( .A(n17971), .B(n17972), .Z(n17970) );
  XOR U18139 ( .A(n17925), .B(n17973), .Z(n17862) );
  IV U18140 ( .A(n17974), .Z(n17925) );
  XNOR U18141 ( .A(key[625]), .B(n17924), .Z(n17965) );
  XNOR U18142 ( .A(n17952), .B(n17975), .Z(n17924) );
  XNOR U18143 ( .A(n17976), .B(n17977), .Z(n17975) );
  XNOR U18144 ( .A(n17978), .B(n17979), .Z(n17952) );
  XOR U18145 ( .A(n17264), .B(n15172), .Z(n17258) );
  XNOR U18146 ( .A(n17836), .B(n15135), .Z(n15172) );
  XOR U18147 ( .A(n17922), .B(n17920), .Z(n15135) );
  XNOR U18148 ( .A(n17911), .B(n17980), .Z(n17836) );
  XOR U18149 ( .A(n17981), .B(n17982), .Z(n17980) );
  XOR U18150 ( .A(n17985), .B(n17986), .Z(n17911) );
  XNOR U18151 ( .A(n17987), .B(n17988), .Z(n17986) );
  NANDN U18152 ( .A(n17989), .B(n17990), .Z(n17988) );
  XOR U18153 ( .A(n17992), .B(n17913), .Z(n17991) );
  OR U18154 ( .A(n17993), .B(n17994), .Z(n17913) );
  ANDN U18155 ( .B(n17995), .A(n17996), .Z(n17992) );
  XNOR U18156 ( .A(n15146), .B(n17997), .Z(n17962) );
  XOR U18157 ( .A(key[627]), .B(n15148), .Z(n17997) );
  XNOR U18158 ( .A(n16197), .B(n15139), .Z(n15148) );
  XOR U18159 ( .A(n17860), .B(n17998), .Z(n15139) );
  XNOR U18160 ( .A(n17973), .B(n17959), .Z(n17998) );
  XNOR U18161 ( .A(n17999), .B(n18000), .Z(n17959) );
  XNOR U18162 ( .A(n18001), .B(n17892), .Z(n18000) );
  ANDN U18163 ( .B(n18002), .A(n18003), .Z(n17892) );
  ANDN U18164 ( .B(n18004), .A(n17930), .Z(n18001) );
  IV U18165 ( .A(n18005), .Z(n17930) );
  XNOR U18166 ( .A(n17890), .B(n18006), .Z(n17973) );
  XNOR U18167 ( .A(n18007), .B(n18008), .Z(n18006) );
  NANDN U18168 ( .A(n18009), .B(n18010), .Z(n18008) );
  XNOR U18169 ( .A(n17971), .B(n17972), .Z(n17860) );
  XNOR U18170 ( .A(n18007), .B(n18012), .Z(n18011) );
  NANDN U18171 ( .A(n18013), .B(n17889), .Z(n18012) );
  OR U18172 ( .A(n18014), .B(n18015), .Z(n18007) );
  XNOR U18173 ( .A(n17890), .B(n18016), .Z(n17999) );
  XNOR U18174 ( .A(n18017), .B(n18018), .Z(n18016) );
  NANDN U18175 ( .A(n17935), .B(n18019), .Z(n18018) );
  XOR U18176 ( .A(n18020), .B(n18017), .Z(n17890) );
  NANDN U18177 ( .A(n18021), .B(n18022), .Z(n18017) );
  ANDN U18178 ( .B(n18023), .A(n18024), .Z(n18020) );
  XNOR U18179 ( .A(n18025), .B(n18026), .Z(n16197) );
  XOR U18180 ( .A(n17856), .B(n17960), .Z(n18026) );
  XNOR U18181 ( .A(n18027), .B(n18028), .Z(n17960) );
  XNOR U18182 ( .A(n18029), .B(n17878), .Z(n18028) );
  ANDN U18183 ( .B(n18030), .A(n18031), .Z(n17878) );
  NOR U18184 ( .A(n18032), .B(n17942), .Z(n18029) );
  XOR U18185 ( .A(n18027), .B(n18033), .Z(n17856) );
  XNOR U18186 ( .A(n18034), .B(n18035), .Z(n18033) );
  NANDN U18187 ( .A(n18036), .B(n17876), .Z(n18035) );
  XNOR U18188 ( .A(n17870), .B(n18037), .Z(n18027) );
  XNOR U18189 ( .A(n18038), .B(n18039), .Z(n18037) );
  NAND U18190 ( .A(n18040), .B(n17947), .Z(n18039) );
  XNOR U18191 ( .A(n17969), .B(n17859), .Z(n18025) );
  XOR U18192 ( .A(n17870), .B(n18041), .Z(n17969) );
  XNOR U18193 ( .A(n18034), .B(n18042), .Z(n18041) );
  NANDN U18194 ( .A(n18043), .B(n18044), .Z(n18042) );
  OR U18195 ( .A(n18045), .B(n18046), .Z(n18034) );
  XOR U18196 ( .A(n18047), .B(n18038), .Z(n17870) );
  NANDN U18197 ( .A(n18048), .B(n18049), .Z(n18038) );
  ANDN U18198 ( .B(n18050), .A(n18051), .Z(n18047) );
  XNOR U18199 ( .A(n16216), .B(n17269), .Z(n15146) );
  XOR U18200 ( .A(n15153), .B(n17898), .Z(n17269) );
  XOR U18201 ( .A(n17979), .B(n17898), .Z(n16216) );
  XOR U18202 ( .A(n17953), .B(n18052), .Z(n17898) );
  XOR U18203 ( .A(n18053), .B(n18054), .Z(n18052) );
  XOR U18204 ( .A(n18057), .B(n18058), .Z(n17953) );
  XNOR U18205 ( .A(n18059), .B(n18060), .Z(n18058) );
  NANDN U18206 ( .A(n18061), .B(n18062), .Z(n18060) );
  XOR U18207 ( .A(n18063), .B(n18064), .Z(n17821) );
  XNOR U18208 ( .A(n16194), .B(n16191), .Z(n18064) );
  XNOR U18209 ( .A(n15158), .B(n15137), .Z(n16191) );
  XOR U18210 ( .A(n17950), .B(n18065), .Z(n15137) );
  XNOR U18211 ( .A(n17978), .B(n17961), .Z(n18065) );
  XNOR U18212 ( .A(n18066), .B(n18067), .Z(n17961) );
  XNOR U18213 ( .A(n18068), .B(n17902), .Z(n18067) );
  NOR U18214 ( .A(n18069), .B(n18070), .Z(n17902) );
  ANDN U18215 ( .B(n18056), .A(n18071), .Z(n18068) );
  XNOR U18216 ( .A(n17900), .B(n18072), .Z(n17978) );
  XNOR U18217 ( .A(n18073), .B(n18074), .Z(n18072) );
  NANDN U18218 ( .A(n18075), .B(n18076), .Z(n18074) );
  XOR U18219 ( .A(n17976), .B(n17977), .Z(n17950) );
  XNOR U18220 ( .A(n18073), .B(n18078), .Z(n18077) );
  NAND U18221 ( .A(n18079), .B(n17958), .Z(n18078) );
  OR U18222 ( .A(n18080), .B(n18081), .Z(n18073) );
  XNOR U18223 ( .A(n17900), .B(n18082), .Z(n18066) );
  XNOR U18224 ( .A(n18083), .B(n18084), .Z(n18082) );
  OR U18225 ( .A(n18061), .B(n18085), .Z(n18084) );
  XOR U18226 ( .A(n18086), .B(n18083), .Z(n17900) );
  OR U18227 ( .A(n18087), .B(n18088), .Z(n18083) );
  ANDN U18228 ( .B(n18089), .A(n18090), .Z(n18086) );
  XOR U18229 ( .A(n17909), .B(n18091), .Z(n15158) );
  XOR U18230 ( .A(n17923), .B(n17866), .Z(n18091) );
  XNOR U18231 ( .A(n18092), .B(n18093), .Z(n17866) );
  XNOR U18232 ( .A(n18094), .B(n17838), .Z(n18093) );
  ANDN U18233 ( .B(n18095), .A(n18096), .Z(n17838) );
  ANDN U18234 ( .B(n17984), .A(n18097), .Z(n18094) );
  XNOR U18235 ( .A(n17834), .B(n18098), .Z(n17923) );
  XNOR U18236 ( .A(n18099), .B(n18100), .Z(n18098) );
  NANDN U18237 ( .A(n18101), .B(n18102), .Z(n18100) );
  XOR U18238 ( .A(n17920), .B(n17921), .Z(n17909) );
  XNOR U18239 ( .A(n18099), .B(n18104), .Z(n18103) );
  NANDN U18240 ( .A(n18105), .B(n17916), .Z(n18104) );
  OR U18241 ( .A(n17993), .B(n18106), .Z(n18099) );
  XNOR U18242 ( .A(n17916), .B(n18102), .Z(n17993) );
  XOR U18243 ( .A(n17834), .B(n18107), .Z(n18092) );
  XNOR U18244 ( .A(n18108), .B(n18109), .Z(n18107) );
  NANDN U18245 ( .A(n17989), .B(n18110), .Z(n18109) );
  XNOR U18246 ( .A(n18111), .B(n18108), .Z(n17834) );
  NANDN U18247 ( .A(n18112), .B(n18113), .Z(n18108) );
  ANDN U18248 ( .B(n18114), .A(n18115), .Z(n18111) );
  XNOR U18249 ( .A(n17985), .B(n18116), .Z(n17920) );
  XNOR U18250 ( .A(n17982), .B(n18117), .Z(n18116) );
  NANDN U18251 ( .A(n18118), .B(n17840), .Z(n18117) );
  XOR U18252 ( .A(n17984), .B(n17840), .Z(n18095) );
  XNOR U18253 ( .A(n18120), .B(n17987), .Z(n17985) );
  OR U18254 ( .A(n18112), .B(n18121), .Z(n17987) );
  XNOR U18255 ( .A(n18115), .B(n17989), .Z(n18112) );
  XNOR U18256 ( .A(n18102), .B(n17840), .Z(n17989) );
  XOR U18257 ( .A(n18122), .B(n18123), .Z(n17840) );
  NANDN U18258 ( .A(n18124), .B(n18125), .Z(n18123) );
  IV U18259 ( .A(n17996), .Z(n18102) );
  XNOR U18260 ( .A(n18126), .B(n18127), .Z(n17996) );
  NANDN U18261 ( .A(n18124), .B(n18128), .Z(n18127) );
  NOR U18262 ( .A(n18115), .B(n18129), .Z(n18120) );
  XNOR U18263 ( .A(n17984), .B(n17916), .Z(n18115) );
  XNOR U18264 ( .A(n18130), .B(n18126), .Z(n17916) );
  NANDN U18265 ( .A(n18131), .B(n18132), .Z(n18126) );
  XOR U18266 ( .A(n18128), .B(n18133), .Z(n18132) );
  ANDN U18267 ( .B(n18133), .A(n18134), .Z(n18130) );
  XNOR U18268 ( .A(n18135), .B(n18122), .Z(n17984) );
  NANDN U18269 ( .A(n18131), .B(n18136), .Z(n18122) );
  XOR U18270 ( .A(n18137), .B(n18125), .Z(n18136) );
  XNOR U18271 ( .A(n18138), .B(n18139), .Z(n18124) );
  XOR U18272 ( .A(n18140), .B(n18141), .Z(n18139) );
  XNOR U18273 ( .A(n18142), .B(n18143), .Z(n18138) );
  XNOR U18274 ( .A(n18144), .B(n18145), .Z(n18143) );
  ANDN U18275 ( .B(n18137), .A(n18141), .Z(n18144) );
  ANDN U18276 ( .B(n18137), .A(n18134), .Z(n18135) );
  XNOR U18277 ( .A(n18140), .B(n18146), .Z(n18134) );
  XOR U18278 ( .A(n18147), .B(n18145), .Z(n18146) );
  NAND U18279 ( .A(n18148), .B(n18149), .Z(n18145) );
  XNOR U18280 ( .A(n18142), .B(n18125), .Z(n18149) );
  IV U18281 ( .A(n18137), .Z(n18142) );
  XNOR U18282 ( .A(n18128), .B(n18141), .Z(n18148) );
  IV U18283 ( .A(n18133), .Z(n18141) );
  XOR U18284 ( .A(n18150), .B(n18151), .Z(n18133) );
  XNOR U18285 ( .A(n18152), .B(n18153), .Z(n18151) );
  XNOR U18286 ( .A(n18154), .B(n18155), .Z(n18150) );
  NOR U18287 ( .A(n18097), .B(n17983), .Z(n18154) );
  AND U18288 ( .A(n18125), .B(n18128), .Z(n18147) );
  XNOR U18289 ( .A(n18125), .B(n18128), .Z(n18140) );
  XNOR U18290 ( .A(n18156), .B(n18157), .Z(n18128) );
  XNOR U18291 ( .A(n18158), .B(n18153), .Z(n18157) );
  XOR U18292 ( .A(n18159), .B(n18160), .Z(n18156) );
  XNOR U18293 ( .A(n18161), .B(n18155), .Z(n18160) );
  OR U18294 ( .A(n18096), .B(n18119), .Z(n18155) );
  XNOR U18295 ( .A(n17983), .B(n18118), .Z(n18119) );
  XNOR U18296 ( .A(n18097), .B(n17841), .Z(n18096) );
  ANDN U18297 ( .B(n18162), .A(n18118), .Z(n18161) );
  XNOR U18298 ( .A(n18163), .B(n18164), .Z(n18125) );
  XNOR U18299 ( .A(n18153), .B(n18165), .Z(n18164) );
  XOR U18300 ( .A(n18105), .B(n18159), .Z(n18165) );
  XNOR U18301 ( .A(n17983), .B(n18166), .Z(n18153) );
  XNOR U18302 ( .A(n18167), .B(n18168), .Z(n18163) );
  XNOR U18303 ( .A(n18169), .B(n18170), .Z(n18168) );
  ANDN U18304 ( .B(n17995), .A(n18101), .Z(n18169) );
  XNOR U18305 ( .A(n18171), .B(n18172), .Z(n18137) );
  XNOR U18306 ( .A(n18158), .B(n18173), .Z(n18172) );
  XNOR U18307 ( .A(n18101), .B(n18152), .Z(n18173) );
  XOR U18308 ( .A(n18159), .B(n18174), .Z(n18152) );
  XNOR U18309 ( .A(n18175), .B(n18176), .Z(n18174) );
  NAND U18310 ( .A(n17990), .B(n18110), .Z(n18176) );
  XNOR U18311 ( .A(n18177), .B(n18175), .Z(n18159) );
  NANDN U18312 ( .A(n18121), .B(n18113), .Z(n18175) );
  XOR U18313 ( .A(n18114), .B(n18110), .Z(n18113) );
  XNOR U18314 ( .A(n18178), .B(n17841), .Z(n18110) );
  XOR U18315 ( .A(n18129), .B(n17990), .Z(n18121) );
  XOR U18316 ( .A(n17995), .B(n18179), .Z(n17990) );
  ANDN U18317 ( .B(n18114), .A(n18129), .Z(n18177) );
  XOR U18318 ( .A(n18167), .B(n17983), .Z(n18129) );
  XOR U18319 ( .A(n18180), .B(n18181), .Z(n17983) );
  XNOR U18320 ( .A(n18182), .B(n18183), .Z(n18181) );
  XOR U18321 ( .A(n18184), .B(n18166), .Z(n18114) );
  XOR U18322 ( .A(n18179), .B(n18162), .Z(n18158) );
  IV U18323 ( .A(n17841), .Z(n18162) );
  XOR U18324 ( .A(n18185), .B(n18186), .Z(n17841) );
  XNOR U18325 ( .A(n18187), .B(n18183), .Z(n18186) );
  IV U18326 ( .A(n18118), .Z(n18179) );
  XOR U18327 ( .A(n18183), .B(n18188), .Z(n18118) );
  XNOR U18328 ( .A(n17995), .B(n18189), .Z(n18171) );
  XNOR U18329 ( .A(n18190), .B(n18170), .Z(n18189) );
  OR U18330 ( .A(n18106), .B(n17994), .Z(n18170) );
  XNOR U18331 ( .A(n18167), .B(n17995), .Z(n17994) );
  XOR U18332 ( .A(n18105), .B(n18178), .Z(n18106) );
  IV U18333 ( .A(n18101), .Z(n18178) );
  XOR U18334 ( .A(n18166), .B(n18191), .Z(n18101) );
  XNOR U18335 ( .A(n18187), .B(n18180), .Z(n18191) );
  XOR U18336 ( .A(n18192), .B(n18193), .Z(n18180) );
  XOR U18337 ( .A(n18194), .B(n18195), .Z(n18193) );
  XOR U18338 ( .A(key[466]), .B(n18196), .Z(n18192) );
  IV U18339 ( .A(n18097), .Z(n18166) );
  XOR U18340 ( .A(n18185), .B(n18197), .Z(n18097) );
  XOR U18341 ( .A(n18183), .B(n18198), .Z(n18197) );
  ANDN U18342 ( .B(n18184), .A(n17915), .Z(n18190) );
  IV U18343 ( .A(n18105), .Z(n18184) );
  XOR U18344 ( .A(n18185), .B(n18199), .Z(n18105) );
  XOR U18345 ( .A(n18183), .B(n18200), .Z(n18199) );
  XOR U18346 ( .A(n18201), .B(n18202), .Z(n18183) );
  XNOR U18347 ( .A(n18203), .B(n17915), .Z(n18202) );
  IV U18348 ( .A(n18167), .Z(n17915) );
  XOR U18349 ( .A(n18204), .B(n18205), .Z(n18201) );
  XNOR U18350 ( .A(key[470]), .B(n18206), .Z(n18205) );
  IV U18351 ( .A(n18188), .Z(n18185) );
  XOR U18352 ( .A(n18207), .B(n18208), .Z(n18188) );
  XOR U18353 ( .A(n18209), .B(n18210), .Z(n18208) );
  XNOR U18354 ( .A(key[469]), .B(n18211), .Z(n18207) );
  XOR U18355 ( .A(n18212), .B(n18213), .Z(n17995) );
  XNOR U18356 ( .A(n18200), .B(n18198), .Z(n18213) );
  XNOR U18357 ( .A(n18214), .B(n18215), .Z(n18198) );
  XOR U18358 ( .A(n18216), .B(n18217), .Z(n18215) );
  XOR U18359 ( .A(key[471]), .B(n18218), .Z(n18214) );
  XNOR U18360 ( .A(n18219), .B(n18220), .Z(n18200) );
  XNOR U18361 ( .A(n18221), .B(n18222), .Z(n18220) );
  XOR U18362 ( .A(n18223), .B(n18224), .Z(n18219) );
  XNOR U18363 ( .A(key[468]), .B(n18225), .Z(n18224) );
  XOR U18364 ( .A(n18167), .B(n18182), .Z(n18212) );
  XOR U18365 ( .A(n18226), .B(n18227), .Z(n18182) );
  XNOR U18366 ( .A(n18187), .B(n18228), .Z(n18227) );
  XNOR U18367 ( .A(n18229), .B(n18230), .Z(n18228) );
  XOR U18368 ( .A(n18231), .B(n18232), .Z(n18187) );
  XNOR U18369 ( .A(n18233), .B(n18234), .Z(n18232) );
  XNOR U18370 ( .A(key[465]), .B(n18235), .Z(n18231) );
  XOR U18371 ( .A(n18236), .B(n18237), .Z(n18226) );
  XNOR U18372 ( .A(key[467]), .B(n18238), .Z(n18237) );
  XOR U18373 ( .A(n18239), .B(n18240), .Z(n18167) );
  IV U18374 ( .A(n15136), .Z(n16194) );
  XOR U18375 ( .A(n15155), .B(n16185), .Z(n15136) );
  XOR U18376 ( .A(n17937), .B(n17968), .Z(n16185) );
  IV U18377 ( .A(n17859), .Z(n17968) );
  XOR U18378 ( .A(n17943), .B(n18244), .Z(n17859) );
  XNOR U18379 ( .A(n17940), .B(n18245), .Z(n18244) );
  NANDN U18380 ( .A(n18246), .B(n17880), .Z(n18245) );
  XNOR U18381 ( .A(n17942), .B(n17880), .Z(n18030) );
  XOR U18382 ( .A(n18249), .B(n17873), .Z(n18248) );
  OR U18383 ( .A(n18045), .B(n18250), .Z(n17873) );
  XNOR U18384 ( .A(n17876), .B(n18044), .Z(n18045) );
  ANDN U18385 ( .B(n18251), .A(n18252), .Z(n18249) );
  XNOR U18386 ( .A(n18253), .B(n17945), .Z(n17943) );
  OR U18387 ( .A(n18048), .B(n18254), .Z(n17945) );
  XOR U18388 ( .A(n18051), .B(n17947), .Z(n18048) );
  XOR U18389 ( .A(n18044), .B(n17880), .Z(n17947) );
  XOR U18390 ( .A(n18255), .B(n18256), .Z(n17880) );
  NANDN U18391 ( .A(n18257), .B(n18258), .Z(n18256) );
  IV U18392 ( .A(n18252), .Z(n18044) );
  XNOR U18393 ( .A(n18259), .B(n18260), .Z(n18252) );
  NANDN U18394 ( .A(n18257), .B(n18261), .Z(n18260) );
  ANDN U18395 ( .B(n18262), .A(n18051), .Z(n18253) );
  XOR U18396 ( .A(n17942), .B(n17876), .Z(n18051) );
  XNOR U18397 ( .A(n18263), .B(n18259), .Z(n17876) );
  NANDN U18398 ( .A(n18264), .B(n18265), .Z(n18259) );
  XOR U18399 ( .A(n18261), .B(n18266), .Z(n18265) );
  ANDN U18400 ( .B(n18266), .A(n18267), .Z(n18263) );
  XOR U18401 ( .A(n18268), .B(n18255), .Z(n17942) );
  NANDN U18402 ( .A(n18264), .B(n18269), .Z(n18255) );
  XOR U18403 ( .A(n18270), .B(n18258), .Z(n18269) );
  XNOR U18404 ( .A(n18271), .B(n18272), .Z(n18257) );
  XOR U18405 ( .A(n18273), .B(n18274), .Z(n18272) );
  XNOR U18406 ( .A(n18275), .B(n18276), .Z(n18271) );
  XNOR U18407 ( .A(n18277), .B(n18278), .Z(n18276) );
  ANDN U18408 ( .B(n18270), .A(n18274), .Z(n18277) );
  ANDN U18409 ( .B(n18270), .A(n18267), .Z(n18268) );
  XNOR U18410 ( .A(n18273), .B(n18279), .Z(n18267) );
  XOR U18411 ( .A(n18280), .B(n18278), .Z(n18279) );
  NAND U18412 ( .A(n18281), .B(n18282), .Z(n18278) );
  XNOR U18413 ( .A(n18275), .B(n18258), .Z(n18282) );
  IV U18414 ( .A(n18270), .Z(n18275) );
  XNOR U18415 ( .A(n18261), .B(n18274), .Z(n18281) );
  IV U18416 ( .A(n18266), .Z(n18274) );
  XOR U18417 ( .A(n18283), .B(n18284), .Z(n18266) );
  XNOR U18418 ( .A(n18285), .B(n18286), .Z(n18284) );
  XNOR U18419 ( .A(n18287), .B(n18288), .Z(n18283) );
  NOR U18420 ( .A(n18032), .B(n17941), .Z(n18287) );
  AND U18421 ( .A(n18258), .B(n18261), .Z(n18280) );
  XNOR U18422 ( .A(n18258), .B(n18261), .Z(n18273) );
  XNOR U18423 ( .A(n18289), .B(n18290), .Z(n18261) );
  XNOR U18424 ( .A(n18291), .B(n18286), .Z(n18290) );
  XOR U18425 ( .A(n18292), .B(n18293), .Z(n18289) );
  XNOR U18426 ( .A(n18294), .B(n18288), .Z(n18293) );
  OR U18427 ( .A(n18031), .B(n18247), .Z(n18288) );
  XNOR U18428 ( .A(n17941), .B(n18246), .Z(n18247) );
  XNOR U18429 ( .A(n18032), .B(n17881), .Z(n18031) );
  ANDN U18430 ( .B(n18295), .A(n18246), .Z(n18294) );
  XNOR U18431 ( .A(n18296), .B(n18297), .Z(n18258) );
  XNOR U18432 ( .A(n18286), .B(n18298), .Z(n18297) );
  XOR U18433 ( .A(n18036), .B(n18292), .Z(n18298) );
  XNOR U18434 ( .A(n17941), .B(n18299), .Z(n18286) );
  XNOR U18435 ( .A(n18300), .B(n18301), .Z(n18296) );
  XNOR U18436 ( .A(n18302), .B(n18303), .Z(n18301) );
  ANDN U18437 ( .B(n18251), .A(n18043), .Z(n18302) );
  XNOR U18438 ( .A(n18304), .B(n18305), .Z(n18270) );
  XNOR U18439 ( .A(n18291), .B(n18306), .Z(n18305) );
  XNOR U18440 ( .A(n18043), .B(n18285), .Z(n18306) );
  XOR U18441 ( .A(n18292), .B(n18307), .Z(n18285) );
  XNOR U18442 ( .A(n18308), .B(n18309), .Z(n18307) );
  NAND U18443 ( .A(n17948), .B(n18040), .Z(n18309) );
  XNOR U18444 ( .A(n18310), .B(n18308), .Z(n18292) );
  NANDN U18445 ( .A(n18254), .B(n18049), .Z(n18308) );
  XOR U18446 ( .A(n18050), .B(n18040), .Z(n18049) );
  XNOR U18447 ( .A(n18311), .B(n17881), .Z(n18040) );
  XOR U18448 ( .A(n18312), .B(n17948), .Z(n18254) );
  XOR U18449 ( .A(n18251), .B(n18313), .Z(n17948) );
  ANDN U18450 ( .B(n18050), .A(n18312), .Z(n18310) );
  IV U18451 ( .A(n18262), .Z(n18312) );
  XOR U18452 ( .A(n18314), .B(n18299), .Z(n18050) );
  XOR U18453 ( .A(n18313), .B(n18295), .Z(n18291) );
  IV U18454 ( .A(n17881), .Z(n18295) );
  XOR U18455 ( .A(n18315), .B(n18316), .Z(n17881) );
  XNOR U18456 ( .A(n18317), .B(n18318), .Z(n18316) );
  IV U18457 ( .A(n18246), .Z(n18313) );
  XOR U18458 ( .A(n18318), .B(n18319), .Z(n18246) );
  XNOR U18459 ( .A(n18251), .B(n18320), .Z(n18304) );
  XNOR U18460 ( .A(n18321), .B(n18303), .Z(n18320) );
  OR U18461 ( .A(n18046), .B(n18250), .Z(n18303) );
  XNOR U18462 ( .A(n18300), .B(n18251), .Z(n18250) );
  XOR U18463 ( .A(n18036), .B(n18311), .Z(n18046) );
  IV U18464 ( .A(n18043), .Z(n18311) );
  XOR U18465 ( .A(n18299), .B(n18322), .Z(n18043) );
  XNOR U18466 ( .A(n18317), .B(n18323), .Z(n18322) );
  IV U18467 ( .A(n18032), .Z(n18299) );
  XOR U18468 ( .A(n18315), .B(n18324), .Z(n18032) );
  XOR U18469 ( .A(n18318), .B(n18325), .Z(n18324) );
  ANDN U18470 ( .B(n18314), .A(n17875), .Z(n18321) );
  IV U18471 ( .A(n18036), .Z(n18314) );
  XOR U18472 ( .A(n18315), .B(n18326), .Z(n18036) );
  XOR U18473 ( .A(n18318), .B(n18327), .Z(n18326) );
  IV U18474 ( .A(n18319), .Z(n18315) );
  XOR U18475 ( .A(n18328), .B(n18329), .Z(n18319) );
  XOR U18476 ( .A(n18330), .B(n18331), .Z(n18329) );
  XNOR U18477 ( .A(n18332), .B(n18333), .Z(n18328) );
  XNOR U18478 ( .A(key[509]), .B(n18334), .Z(n18333) );
  XOR U18479 ( .A(n18335), .B(n18336), .Z(n18251) );
  XNOR U18480 ( .A(n18327), .B(n18325), .Z(n18336) );
  XNOR U18481 ( .A(n18337), .B(n18338), .Z(n18325) );
  XNOR U18482 ( .A(n18339), .B(n18340), .Z(n18338) );
  XNOR U18483 ( .A(n18342), .B(n18343), .Z(n18327) );
  XOR U18484 ( .A(n18344), .B(n18345), .Z(n18343) );
  XNOR U18485 ( .A(n18346), .B(n18347), .Z(n18342) );
  XNOR U18486 ( .A(key[508]), .B(n18348), .Z(n18347) );
  XOR U18487 ( .A(n18300), .B(n18349), .Z(n18335) );
  XOR U18488 ( .A(n17875), .B(n17941), .Z(n18262) );
  XOR U18489 ( .A(n18323), .B(n18350), .Z(n17941) );
  XNOR U18490 ( .A(n18349), .B(n18318), .Z(n18350) );
  XOR U18491 ( .A(n18351), .B(n18352), .Z(n18318) );
  XOR U18492 ( .A(n18353), .B(n17875), .Z(n18352) );
  XOR U18493 ( .A(n18354), .B(n18355), .Z(n18351) );
  XOR U18494 ( .A(key[510]), .B(n18356), .Z(n18355) );
  XOR U18495 ( .A(n18357), .B(n18358), .Z(n18349) );
  XNOR U18496 ( .A(n18317), .B(n18359), .Z(n18358) );
  XNOR U18497 ( .A(n18360), .B(n18361), .Z(n18359) );
  XOR U18498 ( .A(n18362), .B(n18363), .Z(n18317) );
  XOR U18499 ( .A(n18364), .B(n18365), .Z(n18363) );
  XOR U18500 ( .A(n18366), .B(n18367), .Z(n18362) );
  XOR U18501 ( .A(key[505]), .B(n18368), .Z(n18367) );
  XNOR U18502 ( .A(n18369), .B(n18370), .Z(n18357) );
  XNOR U18503 ( .A(key[507]), .B(n18371), .Z(n18370) );
  XOR U18504 ( .A(n18372), .B(n18373), .Z(n18323) );
  XNOR U18505 ( .A(n18374), .B(n18375), .Z(n18373) );
  XOR U18506 ( .A(n18376), .B(n18377), .Z(n18372) );
  XNOR U18507 ( .A(key[506]), .B(n18378), .Z(n18377) );
  IV U18508 ( .A(n18300), .Z(n17875) );
  XOR U18509 ( .A(n18379), .B(n18380), .Z(n18300) );
  XOR U18510 ( .A(n18381), .B(n18382), .Z(n18380) );
  XNOR U18511 ( .A(n18383), .B(n18384), .Z(n18379) );
  XOR U18512 ( .A(n17971), .B(n17974), .Z(n15155) );
  XNOR U18513 ( .A(n17931), .B(n18386), .Z(n17974) );
  XOR U18514 ( .A(n18387), .B(n17886), .Z(n18386) );
  OR U18515 ( .A(n18388), .B(n18014), .Z(n17886) );
  XNOR U18516 ( .A(n17889), .B(n18010), .Z(n18014) );
  ANDN U18517 ( .B(n18389), .A(n18390), .Z(n18387) );
  XNOR U18518 ( .A(n17931), .B(n18391), .Z(n17971) );
  XOR U18519 ( .A(n17928), .B(n18392), .Z(n18391) );
  NANDN U18520 ( .A(n18393), .B(n17894), .Z(n18392) );
  XOR U18521 ( .A(n18005), .B(n17894), .Z(n18002) );
  XOR U18522 ( .A(n18395), .B(n17933), .Z(n17931) );
  OR U18523 ( .A(n18021), .B(n18396), .Z(n17933) );
  XNOR U18524 ( .A(n18024), .B(n17935), .Z(n18021) );
  XNOR U18525 ( .A(n18010), .B(n17894), .Z(n17935) );
  XOR U18526 ( .A(n18397), .B(n18398), .Z(n17894) );
  NANDN U18527 ( .A(n18399), .B(n18400), .Z(n18398) );
  IV U18528 ( .A(n18390), .Z(n18010) );
  XNOR U18529 ( .A(n18401), .B(n18402), .Z(n18390) );
  NANDN U18530 ( .A(n18399), .B(n18403), .Z(n18402) );
  NOR U18531 ( .A(n18024), .B(n18404), .Z(n18395) );
  XNOR U18532 ( .A(n18005), .B(n17889), .Z(n18024) );
  XNOR U18533 ( .A(n18405), .B(n18401), .Z(n17889) );
  NANDN U18534 ( .A(n18406), .B(n18407), .Z(n18401) );
  XOR U18535 ( .A(n18403), .B(n18408), .Z(n18407) );
  ANDN U18536 ( .B(n18408), .A(n18409), .Z(n18405) );
  XNOR U18537 ( .A(n18410), .B(n18397), .Z(n18005) );
  NANDN U18538 ( .A(n18406), .B(n18411), .Z(n18397) );
  XOR U18539 ( .A(n18412), .B(n18400), .Z(n18411) );
  XNOR U18540 ( .A(n18413), .B(n18414), .Z(n18399) );
  XOR U18541 ( .A(n18415), .B(n18416), .Z(n18414) );
  XNOR U18542 ( .A(n18417), .B(n18418), .Z(n18413) );
  XNOR U18543 ( .A(n18419), .B(n18420), .Z(n18418) );
  ANDN U18544 ( .B(n18412), .A(n18416), .Z(n18419) );
  ANDN U18545 ( .B(n18412), .A(n18409), .Z(n18410) );
  XNOR U18546 ( .A(n18415), .B(n18421), .Z(n18409) );
  XOR U18547 ( .A(n18422), .B(n18420), .Z(n18421) );
  NAND U18548 ( .A(n18423), .B(n18424), .Z(n18420) );
  XNOR U18549 ( .A(n18417), .B(n18400), .Z(n18424) );
  IV U18550 ( .A(n18412), .Z(n18417) );
  XNOR U18551 ( .A(n18403), .B(n18416), .Z(n18423) );
  IV U18552 ( .A(n18408), .Z(n18416) );
  XOR U18553 ( .A(n18425), .B(n18426), .Z(n18408) );
  XNOR U18554 ( .A(n18427), .B(n18428), .Z(n18426) );
  XNOR U18555 ( .A(n18429), .B(n18430), .Z(n18425) );
  ANDN U18556 ( .B(n17929), .A(n18431), .Z(n18429) );
  AND U18557 ( .A(n18400), .B(n18403), .Z(n18422) );
  XNOR U18558 ( .A(n18400), .B(n18403), .Z(n18415) );
  XNOR U18559 ( .A(n18432), .B(n18433), .Z(n18403) );
  XNOR U18560 ( .A(n18434), .B(n18428), .Z(n18433) );
  XOR U18561 ( .A(n18435), .B(n18436), .Z(n18432) );
  XNOR U18562 ( .A(n18437), .B(n18430), .Z(n18436) );
  OR U18563 ( .A(n18003), .B(n18394), .Z(n18430) );
  XNOR U18564 ( .A(n17929), .B(n18438), .Z(n18394) );
  XNOR U18565 ( .A(n18431), .B(n17895), .Z(n18003) );
  ANDN U18566 ( .B(n18439), .A(n18393), .Z(n18437) );
  XNOR U18567 ( .A(n18440), .B(n18441), .Z(n18400) );
  XNOR U18568 ( .A(n18428), .B(n18442), .Z(n18441) );
  XOR U18569 ( .A(n18013), .B(n18435), .Z(n18442) );
  XNOR U18570 ( .A(n17929), .B(n18431), .Z(n18428) );
  XNOR U18571 ( .A(n18443), .B(n18444), .Z(n18440) );
  XNOR U18572 ( .A(n18445), .B(n18446), .Z(n18444) );
  ANDN U18573 ( .B(n18389), .A(n18009), .Z(n18445) );
  XNOR U18574 ( .A(n18447), .B(n18448), .Z(n18412) );
  XNOR U18575 ( .A(n18434), .B(n18449), .Z(n18448) );
  XNOR U18576 ( .A(n18009), .B(n18427), .Z(n18449) );
  XOR U18577 ( .A(n18435), .B(n18450), .Z(n18427) );
  XNOR U18578 ( .A(n18451), .B(n18452), .Z(n18450) );
  NAND U18579 ( .A(n17936), .B(n18019), .Z(n18452) );
  XNOR U18580 ( .A(n18453), .B(n18451), .Z(n18435) );
  NANDN U18581 ( .A(n18396), .B(n18022), .Z(n18451) );
  XOR U18582 ( .A(n18023), .B(n18019), .Z(n18022) );
  XNOR U18583 ( .A(n18454), .B(n17895), .Z(n18019) );
  XOR U18584 ( .A(n18404), .B(n17936), .Z(n18396) );
  XOR U18585 ( .A(n18389), .B(n18438), .Z(n17936) );
  ANDN U18586 ( .B(n18023), .A(n18404), .Z(n18453) );
  XNOR U18587 ( .A(n18443), .B(n17929), .Z(n18404) );
  XNOR U18588 ( .A(n18455), .B(n18456), .Z(n17929) );
  XNOR U18589 ( .A(n18457), .B(n18458), .Z(n18456) );
  XOR U18590 ( .A(n18459), .B(n18004), .Z(n18023) );
  XOR U18591 ( .A(n18438), .B(n18439), .Z(n18434) );
  IV U18592 ( .A(n17895), .Z(n18439) );
  XOR U18593 ( .A(n18460), .B(n18461), .Z(n17895) );
  XNOR U18594 ( .A(n18462), .B(n18458), .Z(n18461) );
  IV U18595 ( .A(n18393), .Z(n18438) );
  XOR U18596 ( .A(n18458), .B(n18463), .Z(n18393) );
  XNOR U18597 ( .A(n18389), .B(n18464), .Z(n18447) );
  XNOR U18598 ( .A(n18465), .B(n18446), .Z(n18464) );
  OR U18599 ( .A(n18015), .B(n18388), .Z(n18446) );
  XNOR U18600 ( .A(n18443), .B(n18389), .Z(n18388) );
  XOR U18601 ( .A(n18013), .B(n18454), .Z(n18015) );
  IV U18602 ( .A(n18009), .Z(n18454) );
  XOR U18603 ( .A(n18004), .B(n18466), .Z(n18009) );
  XNOR U18604 ( .A(n18462), .B(n18455), .Z(n18466) );
  XOR U18605 ( .A(n18467), .B(n18468), .Z(n18455) );
  XOR U18606 ( .A(n18469), .B(n18470), .Z(n18468) );
  XOR U18607 ( .A(key[386]), .B(n18471), .Z(n18467) );
  IV U18608 ( .A(n18431), .Z(n18004) );
  XOR U18609 ( .A(n18460), .B(n18472), .Z(n18431) );
  XOR U18610 ( .A(n18458), .B(n18473), .Z(n18472) );
  ANDN U18611 ( .B(n18459), .A(n17888), .Z(n18465) );
  IV U18612 ( .A(n18013), .Z(n18459) );
  XOR U18613 ( .A(n18460), .B(n18474), .Z(n18013) );
  XOR U18614 ( .A(n18458), .B(n18475), .Z(n18474) );
  XOR U18615 ( .A(n18476), .B(n18477), .Z(n18458) );
  XNOR U18616 ( .A(n18478), .B(n17888), .Z(n18477) );
  IV U18617 ( .A(n18443), .Z(n17888) );
  XOR U18618 ( .A(n18479), .B(n18480), .Z(n18476) );
  XNOR U18619 ( .A(key[390]), .B(n18481), .Z(n18480) );
  IV U18620 ( .A(n18463), .Z(n18460) );
  XOR U18621 ( .A(n18482), .B(n18483), .Z(n18463) );
  XNOR U18622 ( .A(n18484), .B(n18485), .Z(n18483) );
  XNOR U18623 ( .A(key[389]), .B(n18486), .Z(n18482) );
  XOR U18624 ( .A(n18487), .B(n18488), .Z(n18389) );
  XNOR U18625 ( .A(n18475), .B(n18473), .Z(n18488) );
  XNOR U18626 ( .A(n18489), .B(n18490), .Z(n18473) );
  XOR U18627 ( .A(n18491), .B(n18492), .Z(n18490) );
  XNOR U18628 ( .A(key[391]), .B(n18493), .Z(n18489) );
  XNOR U18629 ( .A(n18494), .B(n18495), .Z(n18475) );
  XNOR U18630 ( .A(n18496), .B(n18497), .Z(n18495) );
  XOR U18631 ( .A(n18498), .B(n18499), .Z(n18494) );
  XOR U18632 ( .A(key[388]), .B(n18500), .Z(n18499) );
  XOR U18633 ( .A(n18443), .B(n18457), .Z(n18487) );
  XOR U18634 ( .A(n18501), .B(n18502), .Z(n18457) );
  XNOR U18635 ( .A(n18462), .B(n18503), .Z(n18502) );
  XNOR U18636 ( .A(n18504), .B(n18505), .Z(n18503) );
  XOR U18637 ( .A(n18506), .B(n18507), .Z(n18462) );
  XOR U18638 ( .A(n18508), .B(n18509), .Z(n18507) );
  XOR U18639 ( .A(key[385]), .B(n18510), .Z(n18506) );
  XNOR U18640 ( .A(n18511), .B(n18512), .Z(n18501) );
  XOR U18641 ( .A(key[387]), .B(n18513), .Z(n18512) );
  XOR U18642 ( .A(n18514), .B(n18515), .Z(n18443) );
  XNOR U18643 ( .A(n18516), .B(n18517), .Z(n18515) );
  XNOR U18644 ( .A(key[626]), .B(n15153), .Z(n18063) );
  XOR U18645 ( .A(n17977), .B(n17979), .Z(n15153) );
  XOR U18646 ( .A(n18520), .B(n17955), .Z(n18519) );
  OR U18647 ( .A(n18080), .B(n18521), .Z(n17955) );
  XNOR U18648 ( .A(n17958), .B(n18076), .Z(n18080) );
  ANDN U18649 ( .B(n18076), .A(n18522), .Z(n18520) );
  XNOR U18650 ( .A(n18057), .B(n18523), .Z(n17977) );
  XNOR U18651 ( .A(n18054), .B(n18524), .Z(n18523) );
  NANDN U18652 ( .A(n18525), .B(n17904), .Z(n18524) );
  OR U18653 ( .A(n18526), .B(n18069), .Z(n18054) );
  XNOR U18654 ( .A(n18056), .B(n17904), .Z(n18069) );
  XNOR U18655 ( .A(n18527), .B(n18059), .Z(n18057) );
  NANDN U18656 ( .A(n18088), .B(n18528), .Z(n18059) );
  XOR U18657 ( .A(n18089), .B(n18061), .Z(n18088) );
  XNOR U18658 ( .A(n18076), .B(n17904), .Z(n18061) );
  XNOR U18659 ( .A(n18529), .B(n18530), .Z(n17904) );
  NANDN U18660 ( .A(n18531), .B(n18532), .Z(n18530) );
  XOR U18661 ( .A(n18533), .B(n18534), .Z(n18076) );
  NANDN U18662 ( .A(n18531), .B(n18535), .Z(n18534) );
  XOR U18663 ( .A(n18056), .B(n17958), .Z(n18089) );
  XNOR U18664 ( .A(n18537), .B(n18533), .Z(n17958) );
  NANDN U18665 ( .A(n18538), .B(n18539), .Z(n18533) );
  XOR U18666 ( .A(n18535), .B(n18540), .Z(n18539) );
  ANDN U18667 ( .B(n18540), .A(n18541), .Z(n18537) );
  XOR U18668 ( .A(n18542), .B(n18529), .Z(n18056) );
  ANDN U18669 ( .B(n18543), .A(n18538), .Z(n18529) );
  XNOR U18670 ( .A(n18544), .B(n18545), .Z(n18531) );
  XOR U18671 ( .A(n18546), .B(n18547), .Z(n18545) );
  XNOR U18672 ( .A(n18548), .B(n18549), .Z(n18544) );
  XNOR U18673 ( .A(n18550), .B(n18551), .Z(n18549) );
  ANDN U18674 ( .B(n18552), .A(n18547), .Z(n18550) );
  XOR U18675 ( .A(n18552), .B(n18532), .Z(n18543) );
  ANDN U18676 ( .B(n18552), .A(n18541), .Z(n18542) );
  XNOR U18677 ( .A(n18546), .B(n18553), .Z(n18541) );
  XOR U18678 ( .A(n18554), .B(n18551), .Z(n18553) );
  NAND U18679 ( .A(n18555), .B(n18556), .Z(n18551) );
  XNOR U18680 ( .A(n18548), .B(n18532), .Z(n18556) );
  IV U18681 ( .A(n18552), .Z(n18548) );
  XNOR U18682 ( .A(n18535), .B(n18547), .Z(n18555) );
  IV U18683 ( .A(n18540), .Z(n18547) );
  XOR U18684 ( .A(n18557), .B(n18558), .Z(n18540) );
  XNOR U18685 ( .A(n18559), .B(n18560), .Z(n18558) );
  XNOR U18686 ( .A(n18561), .B(n18562), .Z(n18557) );
  ANDN U18687 ( .B(n18563), .A(n18564), .Z(n18561) );
  AND U18688 ( .A(n18532), .B(n18535), .Z(n18554) );
  XNOR U18689 ( .A(n18532), .B(n18535), .Z(n18546) );
  XNOR U18690 ( .A(n18565), .B(n18566), .Z(n18535) );
  XNOR U18691 ( .A(n18567), .B(n18560), .Z(n18566) );
  XOR U18692 ( .A(n18568), .B(n18569), .Z(n18565) );
  XNOR U18693 ( .A(n18570), .B(n18562), .Z(n18569) );
  OR U18694 ( .A(n18070), .B(n18526), .Z(n18562) );
  XNOR U18695 ( .A(n18055), .B(n18601), .Z(n18526) );
  XNOR U18696 ( .A(n18071), .B(n17905), .Z(n18070) );
  ANDN U18697 ( .B(n18571), .A(n18525), .Z(n18570) );
  XNOR U18698 ( .A(n18572), .B(n18573), .Z(n18532) );
  XNOR U18699 ( .A(n18560), .B(n18574), .Z(n18573) );
  XNOR U18700 ( .A(n18079), .B(n18568), .Z(n18574) );
  XNOR U18701 ( .A(n18071), .B(n18055), .Z(n18560) );
  XNOR U18702 ( .A(n18575), .B(n18576), .Z(n18572) );
  XNOR U18703 ( .A(n18577), .B(n18578), .Z(n18576) );
  ANDN U18704 ( .B(n18579), .A(n18522), .Z(n18577) );
  XNOR U18705 ( .A(n18580), .B(n18581), .Z(n18552) );
  XNOR U18706 ( .A(n18567), .B(n18582), .Z(n18581) );
  XNOR U18707 ( .A(n18583), .B(n18559), .Z(n18582) );
  XOR U18708 ( .A(n18568), .B(n18584), .Z(n18559) );
  XNOR U18709 ( .A(n18585), .B(n18586), .Z(n18584) );
  NANDN U18710 ( .A(n18085), .B(n18062), .Z(n18586) );
  XNOR U18711 ( .A(n18587), .B(n18585), .Z(n18568) );
  NANDN U18712 ( .A(n18087), .B(n18528), .Z(n18585) );
  XOR U18713 ( .A(n18536), .B(n18062), .Z(n18528) );
  XNOR U18714 ( .A(n18522), .B(n18601), .Z(n18062) );
  IV U18715 ( .A(n18583), .Z(n18522) );
  XOR U18716 ( .A(n18588), .B(n18085), .Z(n18087) );
  XNOR U18717 ( .A(n18571), .B(n18579), .Z(n18085) );
  IV U18718 ( .A(n17905), .Z(n18571) );
  ANDN U18719 ( .B(n18536), .A(n18090), .Z(n18587) );
  IV U18720 ( .A(n18588), .Z(n18090) );
  XOR U18721 ( .A(n18563), .B(n18079), .Z(n18588) );
  XOR U18722 ( .A(n17905), .B(n18525), .Z(n18567) );
  XOR U18723 ( .A(n18589), .B(n18590), .Z(n18525) );
  XOR U18724 ( .A(n18591), .B(n18592), .Z(n17905) );
  XOR U18725 ( .A(n18593), .B(n18590), .Z(n18592) );
  XNOR U18726 ( .A(n18075), .B(n18594), .Z(n18580) );
  XNOR U18727 ( .A(n18595), .B(n18578), .Z(n18594) );
  OR U18728 ( .A(n18081), .B(n18521), .Z(n18578) );
  XNOR U18729 ( .A(n18575), .B(n18583), .Z(n18521) );
  XOR U18730 ( .A(n18596), .B(n18597), .Z(n18583) );
  XNOR U18731 ( .A(n18598), .B(n18599), .Z(n18597) );
  XOR U18732 ( .A(n18575), .B(n18600), .Z(n18596) );
  XNOR U18733 ( .A(n18079), .B(n18579), .Z(n18081) );
  IV U18734 ( .A(n18075), .Z(n18579) );
  ANDN U18735 ( .B(n18079), .A(n17957), .Z(n18595) );
  XOR U18736 ( .A(n18598), .B(n18601), .Z(n18079) );
  XOR U18737 ( .A(n18602), .B(n18603), .Z(n18598) );
  XNOR U18738 ( .A(n18604), .B(n18605), .Z(n18603) );
  XNOR U18739 ( .A(n18606), .B(n18607), .Z(n18602) );
  XOR U18740 ( .A(key[428]), .B(n18608), .Z(n18607) );
  XNOR U18741 ( .A(n18609), .B(n18610), .Z(n18075) );
  XOR U18742 ( .A(n18071), .B(n18591), .Z(n18610) );
  IV U18743 ( .A(n18563), .Z(n18071) );
  XOR U18744 ( .A(n18600), .B(n18601), .Z(n18563) );
  XNOR U18745 ( .A(n18589), .B(n18590), .Z(n18601) );
  IV U18746 ( .A(n18593), .Z(n18589) );
  XNOR U18747 ( .A(n18611), .B(n18612), .Z(n18593) );
  XOR U18748 ( .A(n18613), .B(n18614), .Z(n18612) );
  XNOR U18749 ( .A(n18615), .B(n18616), .Z(n18611) );
  XNOR U18750 ( .A(key[429]), .B(n18617), .Z(n18616) );
  XOR U18751 ( .A(n18618), .B(n18619), .Z(n18600) );
  XNOR U18752 ( .A(n18620), .B(n18621), .Z(n18619) );
  XOR U18753 ( .A(key[431]), .B(n18622), .Z(n18618) );
  XOR U18754 ( .A(n17957), .B(n18564), .Z(n18536) );
  IV U18755 ( .A(n18055), .Z(n18564) );
  XNOR U18756 ( .A(n18599), .B(n18623), .Z(n18055) );
  XNOR U18757 ( .A(n18590), .B(n18609), .Z(n18623) );
  XOR U18758 ( .A(n18624), .B(n18625), .Z(n18609) );
  XOR U18759 ( .A(n18626), .B(n18627), .Z(n18625) );
  XOR U18760 ( .A(n18628), .B(n18629), .Z(n18624) );
  XNOR U18761 ( .A(key[426]), .B(n18630), .Z(n18629) );
  XOR U18762 ( .A(n18631), .B(n18632), .Z(n18590) );
  XOR U18763 ( .A(n18633), .B(n17957), .Z(n18632) );
  XNOR U18764 ( .A(n18634), .B(n18635), .Z(n18631) );
  XNOR U18765 ( .A(key[430]), .B(n18636), .Z(n18635) );
  XOR U18766 ( .A(n18637), .B(n18638), .Z(n18599) );
  XOR U18767 ( .A(n18591), .B(n18639), .Z(n18638) );
  XNOR U18768 ( .A(n18640), .B(n18641), .Z(n18639) );
  XNOR U18769 ( .A(n18642), .B(n18643), .Z(n18591) );
  XNOR U18770 ( .A(n18644), .B(n18645), .Z(n18643) );
  XOR U18771 ( .A(key[425]), .B(n18647), .Z(n18646) );
  XNOR U18772 ( .A(n18649), .B(n18650), .Z(n18637) );
  XOR U18773 ( .A(key[427]), .B(n18651), .Z(n18650) );
  IV U18774 ( .A(n18575), .Z(n17957) );
  XOR U18775 ( .A(n18652), .B(n18653), .Z(n18575) );
  XOR U18776 ( .A(n18654), .B(n18655), .Z(n18653) );
  XOR U18777 ( .A(n18656), .B(n18657), .Z(n18652) );
  XOR U18778 ( .A(n17621), .B(n17667), .Z(n13413) );
  XNOR U18779 ( .A(n17615), .B(n18659), .Z(n17621) );
  XOR U18780 ( .A(n18660), .B(n18661), .Z(n18659) );
  ANDN U18781 ( .B(n18662), .A(n17677), .Z(n18660) );
  XNOR U18782 ( .A(n18663), .B(n18664), .Z(n17615) );
  XNOR U18783 ( .A(n18665), .B(n18666), .Z(n18664) );
  NAND U18784 ( .A(n18667), .B(n18668), .Z(n18666) );
  XNOR U18785 ( .A(n14428), .B(n14422), .Z(n12286) );
  IV U18786 ( .A(n12309), .Z(n14422) );
  XOR U18787 ( .A(n17526), .B(n17544), .Z(n18669) );
  XOR U18788 ( .A(n17655), .B(n17527), .Z(n17544) );
  XNOR U18789 ( .A(n17630), .B(n18670), .Z(n17527) );
  XNOR U18790 ( .A(n18671), .B(n18672), .Z(n18670) );
  NANDN U18791 ( .A(n18673), .B(n18674), .Z(n18672) );
  IV U18792 ( .A(n17656), .Z(n17655) );
  XNOR U18793 ( .A(n17661), .B(n18675), .Z(n17656) );
  XOR U18794 ( .A(n18676), .B(n17633), .Z(n18675) );
  OR U18795 ( .A(n18677), .B(n18678), .Z(n17633) );
  ANDN U18796 ( .B(n18674), .A(n18679), .Z(n18676) );
  XNOR U18797 ( .A(n17569), .B(n18680), .Z(n17526) );
  XNOR U18798 ( .A(n18671), .B(n18681), .Z(n18680) );
  NANDN U18799 ( .A(n18682), .B(n17636), .Z(n18681) );
  OR U18800 ( .A(n18677), .B(n18683), .Z(n18671) );
  XNOR U18801 ( .A(n17636), .B(n18674), .Z(n18677) );
  XOR U18802 ( .A(n17630), .B(n18684), .Z(n17569) );
  XNOR U18803 ( .A(n18685), .B(n18686), .Z(n18684) );
  NAND U18804 ( .A(n18687), .B(n17665), .Z(n18686) );
  XOR U18805 ( .A(n18688), .B(n18685), .Z(n17630) );
  NANDN U18806 ( .A(n18689), .B(n18690), .Z(n18685) );
  ANDN U18807 ( .B(n18691), .A(n18692), .Z(n18688) );
  XNOR U18808 ( .A(n17661), .B(n18693), .Z(n17524) );
  XNOR U18809 ( .A(n17659), .B(n18694), .Z(n18693) );
  NANDN U18810 ( .A(n18695), .B(n17640), .Z(n18694) );
  NANDN U18811 ( .A(n18696), .B(n17643), .Z(n17659) );
  XNOR U18812 ( .A(n17574), .B(n17640), .Z(n17643) );
  XOR U18813 ( .A(n18697), .B(n17663), .Z(n17661) );
  OR U18814 ( .A(n18689), .B(n18698), .Z(n17663) );
  XNOR U18815 ( .A(n18699), .B(n17665), .Z(n18689) );
  XOR U18816 ( .A(n18674), .B(n17640), .Z(n17665) );
  XOR U18817 ( .A(n18700), .B(n18701), .Z(n17640) );
  NANDN U18818 ( .A(n18702), .B(n18703), .Z(n18701) );
  XOR U18819 ( .A(n18704), .B(n18705), .Z(n18674) );
  NANDN U18820 ( .A(n18702), .B(n18706), .Z(n18705) );
  ANDN U18821 ( .B(n18699), .A(n18707), .Z(n18697) );
  IV U18822 ( .A(n18692), .Z(n18699) );
  XOR U18823 ( .A(n17574), .B(n17636), .Z(n18692) );
  XNOR U18824 ( .A(n18708), .B(n18704), .Z(n17636) );
  NANDN U18825 ( .A(n18709), .B(n18710), .Z(n18704) );
  XOR U18826 ( .A(n18706), .B(n18711), .Z(n18710) );
  ANDN U18827 ( .B(n18711), .A(n18712), .Z(n18708) );
  XOR U18828 ( .A(n18713), .B(n18700), .Z(n17574) );
  NANDN U18829 ( .A(n18709), .B(n18714), .Z(n18700) );
  XOR U18830 ( .A(n18715), .B(n18703), .Z(n18714) );
  XNOR U18831 ( .A(n18716), .B(n18717), .Z(n18702) );
  XOR U18832 ( .A(n18718), .B(n18719), .Z(n18717) );
  XNOR U18833 ( .A(n18720), .B(n18721), .Z(n18716) );
  XNOR U18834 ( .A(n18722), .B(n18723), .Z(n18721) );
  ANDN U18835 ( .B(n18715), .A(n18719), .Z(n18722) );
  ANDN U18836 ( .B(n18715), .A(n18712), .Z(n18713) );
  XNOR U18837 ( .A(n18718), .B(n18724), .Z(n18712) );
  XOR U18838 ( .A(n18725), .B(n18723), .Z(n18724) );
  NAND U18839 ( .A(n18726), .B(n18727), .Z(n18723) );
  XNOR U18840 ( .A(n18720), .B(n18703), .Z(n18727) );
  IV U18841 ( .A(n18715), .Z(n18720) );
  XNOR U18842 ( .A(n18706), .B(n18719), .Z(n18726) );
  IV U18843 ( .A(n18711), .Z(n18719) );
  XOR U18844 ( .A(n18728), .B(n18729), .Z(n18711) );
  XNOR U18845 ( .A(n18730), .B(n18731), .Z(n18729) );
  XNOR U18846 ( .A(n18732), .B(n18733), .Z(n18728) );
  ANDN U18847 ( .B(n17660), .A(n17573), .Z(n18732) );
  AND U18848 ( .A(n18703), .B(n18706), .Z(n18725) );
  XNOR U18849 ( .A(n18703), .B(n18706), .Z(n18718) );
  XNOR U18850 ( .A(n18734), .B(n18735), .Z(n18706) );
  XNOR U18851 ( .A(n18736), .B(n18731), .Z(n18735) );
  XOR U18852 ( .A(n18737), .B(n18738), .Z(n18734) );
  XNOR U18853 ( .A(n18739), .B(n18733), .Z(n18738) );
  OR U18854 ( .A(n17642), .B(n18696), .Z(n18733) );
  XNOR U18855 ( .A(n17660), .B(n18740), .Z(n18696) );
  XNOR U18856 ( .A(n17573), .B(n17641), .Z(n17642) );
  ANDN U18857 ( .B(n18741), .A(n18695), .Z(n18739) );
  XNOR U18858 ( .A(n18742), .B(n18743), .Z(n18703) );
  XNOR U18859 ( .A(n18731), .B(n18744), .Z(n18743) );
  XOR U18860 ( .A(n18682), .B(n18737), .Z(n18744) );
  XNOR U18861 ( .A(n17660), .B(n17573), .Z(n18731) );
  XOR U18862 ( .A(n17635), .B(n18745), .Z(n18742) );
  XNOR U18863 ( .A(n18746), .B(n18747), .Z(n18745) );
  ANDN U18864 ( .B(n18748), .A(n18679), .Z(n18746) );
  XNOR U18865 ( .A(n18749), .B(n18750), .Z(n18715) );
  XNOR U18866 ( .A(n18736), .B(n18751), .Z(n18750) );
  XNOR U18867 ( .A(n18673), .B(n18730), .Z(n18751) );
  XOR U18868 ( .A(n18737), .B(n18752), .Z(n18730) );
  XNOR U18869 ( .A(n18753), .B(n18754), .Z(n18752) );
  NAND U18870 ( .A(n17666), .B(n18687), .Z(n18754) );
  XNOR U18871 ( .A(n18755), .B(n18753), .Z(n18737) );
  NANDN U18872 ( .A(n18698), .B(n18690), .Z(n18753) );
  XOR U18873 ( .A(n18691), .B(n18687), .Z(n18690) );
  XNOR U18874 ( .A(n18748), .B(n17641), .Z(n18687) );
  XOR U18875 ( .A(n18707), .B(n17666), .Z(n18698) );
  XNOR U18876 ( .A(n18679), .B(n18740), .Z(n17666) );
  ANDN U18877 ( .B(n18691), .A(n18707), .Z(n18755) );
  XOR U18878 ( .A(n17635), .B(n17660), .Z(n18707) );
  XNOR U18879 ( .A(n18756), .B(n18757), .Z(n17660) );
  XNOR U18880 ( .A(n18758), .B(n18759), .Z(n18757) );
  XOR U18881 ( .A(n18740), .B(n18741), .Z(n18736) );
  IV U18882 ( .A(n17641), .Z(n18741) );
  XOR U18883 ( .A(n18760), .B(n18761), .Z(n17641) );
  XOR U18884 ( .A(n18762), .B(n18759), .Z(n18761) );
  IV U18885 ( .A(n18695), .Z(n18740) );
  XOR U18886 ( .A(n18759), .B(n18763), .Z(n18695) );
  XNOR U18887 ( .A(n18764), .B(n18765), .Z(n18749) );
  XNOR U18888 ( .A(n18766), .B(n18747), .Z(n18765) );
  OR U18889 ( .A(n18683), .B(n18678), .Z(n18747) );
  XNOR U18890 ( .A(n17635), .B(n18679), .Z(n18678) );
  IV U18891 ( .A(n18764), .Z(n18679) );
  XOR U18892 ( .A(n18682), .B(n18748), .Z(n18683) );
  IV U18893 ( .A(n18673), .Z(n18748) );
  XNOR U18894 ( .A(n18768), .B(n18756), .Z(n18767) );
  XOR U18895 ( .A(n18769), .B(n18770), .Z(n18756) );
  XNOR U18896 ( .A(n15464), .B(n16527), .Z(n18770) );
  XNOR U18897 ( .A(n15463), .B(n15480), .Z(n16527) );
  XOR U18898 ( .A(n18771), .B(n18772), .Z(n15480) );
  XOR U18899 ( .A(n18773), .B(n18774), .Z(n18771) );
  XOR U18900 ( .A(n16495), .B(n18775), .Z(n15464) );
  XOR U18901 ( .A(key[546]), .B(n15486), .Z(n18769) );
  XOR U18902 ( .A(n18760), .B(n18776), .Z(n17573) );
  XOR U18903 ( .A(n18759), .B(n18777), .Z(n18776) );
  NOR U18904 ( .A(n18682), .B(n17635), .Z(n18766) );
  XOR U18905 ( .A(n18760), .B(n18778), .Z(n18682) );
  XOR U18906 ( .A(n18759), .B(n18779), .Z(n18778) );
  XOR U18907 ( .A(n18780), .B(n18781), .Z(n18759) );
  XOR U18908 ( .A(n17635), .B(n16983), .Z(n18781) );
  XNOR U18909 ( .A(n16969), .B(n15459), .Z(n16983) );
  XNOR U18910 ( .A(n18782), .B(n18772), .Z(n15459) );
  XNOR U18911 ( .A(n18783), .B(n18784), .Z(n18772) );
  XNOR U18912 ( .A(n18785), .B(n18786), .Z(n18782) );
  IV U18913 ( .A(n16980), .Z(n16969) );
  XNOR U18914 ( .A(n15470), .B(n18787), .Z(n18780) );
  XNOR U18915 ( .A(key[550]), .B(n15452), .Z(n18787) );
  XOR U18916 ( .A(n16509), .B(n18788), .Z(n15470) );
  XOR U18917 ( .A(n15450), .B(n16503), .Z(n16509) );
  XOR U18918 ( .A(n18789), .B(n18790), .Z(n16503) );
  XOR U18919 ( .A(n18791), .B(n18792), .Z(n15450) );
  IV U18920 ( .A(n18763), .Z(n18760) );
  XOR U18921 ( .A(n18793), .B(n18794), .Z(n18763) );
  XOR U18922 ( .A(n16972), .B(n16981), .Z(n18794) );
  XNOR U18923 ( .A(n15452), .B(n15471), .Z(n16981) );
  XOR U18924 ( .A(n18773), .B(n18795), .Z(n15471) );
  XNOR U18925 ( .A(n18797), .B(n18798), .Z(n18796) );
  ANDN U18926 ( .B(n18799), .A(n18800), .Z(n18797) );
  XNOR U18927 ( .A(n18802), .B(n18803), .Z(n15452) );
  XNOR U18928 ( .A(key[549]), .B(n15451), .Z(n18793) );
  XOR U18929 ( .A(n16511), .B(n16522), .Z(n15451) );
  XNOR U18930 ( .A(n18804), .B(n18805), .Z(n16522) );
  XNOR U18931 ( .A(n18806), .B(n18807), .Z(n18805) );
  XNOR U18932 ( .A(n18808), .B(n18809), .Z(n18804) );
  XOR U18933 ( .A(n18810), .B(n18811), .Z(n18809) );
  ANDN U18934 ( .B(n18812), .A(n18813), .Z(n18811) );
  XOR U18935 ( .A(n18814), .B(n18815), .Z(n16511) );
  XNOR U18936 ( .A(n18816), .B(n18817), .Z(n18815) );
  XNOR U18937 ( .A(n18818), .B(n18819), .Z(n18814) );
  XOR U18938 ( .A(n18820), .B(n18821), .Z(n18819) );
  ANDN U18939 ( .B(n18822), .A(n18823), .Z(n18821) );
  XOR U18940 ( .A(n18824), .B(n18825), .Z(n18764) );
  XNOR U18941 ( .A(n18779), .B(n18777), .Z(n18825) );
  XNOR U18942 ( .A(n18826), .B(n18827), .Z(n18777) );
  XOR U18943 ( .A(n16980), .B(n15458), .Z(n18827) );
  XNOR U18944 ( .A(n16506), .B(n16982), .Z(n15458) );
  XNOR U18945 ( .A(n18828), .B(n18829), .Z(n16982) );
  XOR U18946 ( .A(n18830), .B(n18831), .Z(n18829) );
  XNOR U18947 ( .A(n18817), .B(n18789), .Z(n18828) );
  XNOR U18948 ( .A(n18832), .B(n18833), .Z(n18817) );
  XNOR U18949 ( .A(n18834), .B(n18835), .Z(n18833) );
  OR U18950 ( .A(n18836), .B(n18837), .Z(n18835) );
  XOR U18951 ( .A(n18838), .B(n18839), .Z(n16506) );
  XNOR U18952 ( .A(n18791), .B(n18807), .Z(n18838) );
  XNOR U18953 ( .A(n18840), .B(n18841), .Z(n18807) );
  XNOR U18954 ( .A(n18842), .B(n18843), .Z(n18841) );
  OR U18955 ( .A(n18844), .B(n18845), .Z(n18843) );
  XNOR U18956 ( .A(key[551]), .B(n18788), .Z(n18826) );
  XNOR U18957 ( .A(n16538), .B(n16968), .Z(n18788) );
  XOR U18958 ( .A(n18846), .B(n18847), .Z(n16968) );
  XNOR U18959 ( .A(n18848), .B(n18849), .Z(n18847) );
  XOR U18960 ( .A(n18802), .B(n18850), .Z(n18846) );
  XNOR U18961 ( .A(n18851), .B(n18852), .Z(n18779) );
  XNOR U18962 ( .A(n16956), .B(n16958), .Z(n18852) );
  XNOR U18963 ( .A(n15454), .B(n16980), .Z(n16958) );
  XOR U18964 ( .A(n18853), .B(n18854), .Z(n15454) );
  XNOR U18965 ( .A(n18855), .B(n18785), .Z(n18854) );
  XNOR U18966 ( .A(n18856), .B(n18857), .Z(n18785) );
  XNOR U18967 ( .A(n18858), .B(n18859), .Z(n18857) );
  NANDN U18968 ( .A(n18860), .B(n18861), .Z(n18859) );
  XNOR U18969 ( .A(n18862), .B(n18863), .Z(n18853) );
  XOR U18970 ( .A(n18798), .B(n18864), .Z(n18863) );
  ANDN U18971 ( .B(n18865), .A(n18866), .Z(n18864) );
  NOR U18972 ( .A(n18867), .B(n18868), .Z(n18798) );
  XOR U18973 ( .A(n15440), .B(n18869), .Z(n18851) );
  XNOR U18974 ( .A(key[548]), .B(n15439), .Z(n18869) );
  XNOR U18975 ( .A(n18870), .B(n16972), .Z(n15439) );
  XNOR U18976 ( .A(n18871), .B(n18872), .Z(n16972) );
  XNOR U18977 ( .A(n18873), .B(n18849), .Z(n18872) );
  XNOR U18978 ( .A(n18874), .B(n18875), .Z(n18849) );
  XNOR U18979 ( .A(n18876), .B(n18877), .Z(n18875) );
  NANDN U18980 ( .A(n18878), .B(n18879), .Z(n18877) );
  XNOR U18981 ( .A(n18880), .B(n18881), .Z(n18871) );
  XOR U18982 ( .A(n18882), .B(n18883), .Z(n18881) );
  ANDN U18983 ( .B(n18884), .A(n18885), .Z(n18883) );
  XOR U18984 ( .A(n16520), .B(n16960), .Z(n15440) );
  XOR U18985 ( .A(n18806), .B(n15488), .Z(n16960) );
  IV U18986 ( .A(n18775), .Z(n15488) );
  XOR U18987 ( .A(n18816), .B(n16495), .Z(n16520) );
  XNOR U18988 ( .A(n18888), .B(n18831), .Z(n16495) );
  XNOR U18989 ( .A(n17635), .B(n18758), .Z(n18824) );
  XOR U18990 ( .A(n18889), .B(n18890), .Z(n18758) );
  XNOR U18991 ( .A(n16991), .B(n18891), .Z(n18890) );
  XNOR U18992 ( .A(n15476), .B(n18768), .Z(n18891) );
  IV U18993 ( .A(n18762), .Z(n18768) );
  XNOR U18994 ( .A(n18892), .B(n18893), .Z(n18762) );
  XOR U18995 ( .A(n16537), .B(n16995), .Z(n18893) );
  XNOR U18996 ( .A(n15467), .B(n15486), .Z(n16995) );
  IV U18997 ( .A(n15484), .Z(n16537) );
  XNOR U18998 ( .A(n15491), .B(n16531), .Z(n15484) );
  XNOR U18999 ( .A(n18831), .B(n18894), .Z(n16531) );
  XOR U19000 ( .A(n18789), .B(n18895), .Z(n18894) );
  XNOR U19001 ( .A(n18888), .B(n18896), .Z(n18789) );
  IV U19002 ( .A(n18897), .Z(n18888) );
  XOR U19003 ( .A(n18886), .B(n18898), .Z(n15491) );
  XOR U19004 ( .A(n18900), .B(n18887), .Z(n18791) );
  XOR U19005 ( .A(key[545]), .B(n15492), .Z(n18892) );
  XOR U19006 ( .A(n18870), .B(n16956), .Z(n15476) );
  XOR U19007 ( .A(n18873), .B(n15486), .Z(n16956) );
  XOR U19008 ( .A(n18901), .B(n18850), .Z(n15486) );
  XNOR U19009 ( .A(n16980), .B(n15441), .Z(n16991) );
  XNOR U19010 ( .A(n18862), .B(n15467), .Z(n15441) );
  XOR U19011 ( .A(n18862), .B(n18903), .Z(n16980) );
  XNOR U19012 ( .A(n18856), .B(n18904), .Z(n18862) );
  XOR U19013 ( .A(n18905), .B(n18906), .Z(n18904) );
  ANDN U19014 ( .B(n18907), .A(n18800), .Z(n18905) );
  IV U19015 ( .A(n18908), .Z(n18800) );
  XNOR U19016 ( .A(n18909), .B(n18910), .Z(n18856) );
  XNOR U19017 ( .A(n18911), .B(n18912), .Z(n18910) );
  NAND U19018 ( .A(n18913), .B(n18914), .Z(n18912) );
  XOR U19019 ( .A(n15478), .B(n18915), .Z(n18889) );
  XNOR U19020 ( .A(key[547]), .B(n15463), .Z(n18915) );
  XOR U19021 ( .A(n18916), .B(n18917), .Z(n15463) );
  XOR U19022 ( .A(n18850), .B(n18848), .Z(n18917) );
  XOR U19023 ( .A(n18918), .B(n18803), .Z(n18916) );
  XOR U19024 ( .A(n18919), .B(n18920), .Z(n18803) );
  XNOR U19025 ( .A(n18921), .B(n18882), .Z(n18920) );
  ANDN U19026 ( .B(n18922), .A(n18923), .Z(n18882) );
  NOR U19027 ( .A(n18924), .B(n18925), .Z(n18921) );
  IV U19028 ( .A(n16493), .Z(n15478) );
  XOR U19029 ( .A(n15465), .B(n16533), .Z(n16493) );
  XNOR U19030 ( .A(n18926), .B(n18927), .Z(n16533) );
  XNOR U19031 ( .A(n18895), .B(n18831), .Z(n18927) );
  XOR U19032 ( .A(n18928), .B(n18929), .Z(n18831) );
  XNOR U19033 ( .A(n18930), .B(n18931), .Z(n18929) );
  NANDN U19034 ( .A(n18932), .B(n18822), .Z(n18931) );
  IV U19035 ( .A(n18830), .Z(n18895) );
  XOR U19036 ( .A(n18933), .B(n18934), .Z(n18830) );
  XNOR U19037 ( .A(n18935), .B(n18936), .Z(n18934) );
  NANDN U19038 ( .A(n18836), .B(n18937), .Z(n18936) );
  XNOR U19039 ( .A(n18896), .B(n18790), .Z(n18926) );
  XNOR U19040 ( .A(n18933), .B(n18938), .Z(n18790) );
  XNOR U19041 ( .A(n18939), .B(n18820), .Z(n18938) );
  NOR U19042 ( .A(n18940), .B(n18941), .Z(n18820) );
  NOR U19043 ( .A(n18942), .B(n18943), .Z(n18939) );
  XNOR U19044 ( .A(n18818), .B(n18944), .Z(n18933) );
  XNOR U19045 ( .A(n18945), .B(n18946), .Z(n18944) );
  NAND U19046 ( .A(n18947), .B(n18948), .Z(n18946) );
  XOR U19047 ( .A(n18818), .B(n18949), .Z(n18896) );
  XNOR U19048 ( .A(n18935), .B(n18950), .Z(n18949) );
  NANDN U19049 ( .A(n18951), .B(n18952), .Z(n18950) );
  OR U19050 ( .A(n18953), .B(n18954), .Z(n18935) );
  XOR U19051 ( .A(n18955), .B(n18945), .Z(n18818) );
  OR U19052 ( .A(n18956), .B(n18957), .Z(n18945) );
  XOR U19053 ( .A(n18960), .B(n18839), .Z(n15465) );
  XOR U19054 ( .A(n18899), .B(n18886), .Z(n18839) );
  XOR U19055 ( .A(n18961), .B(n18962), .Z(n18886) );
  XNOR U19056 ( .A(n18963), .B(n18964), .Z(n18962) );
  NANDN U19057 ( .A(n18965), .B(n18812), .Z(n18964) );
  XOR U19058 ( .A(n18966), .B(n18967), .Z(n18899) );
  XNOR U19059 ( .A(n18968), .B(n18969), .Z(n18967) );
  NANDN U19060 ( .A(n18844), .B(n18970), .Z(n18969) );
  XNOR U19061 ( .A(n18900), .B(n18792), .Z(n18960) );
  XNOR U19062 ( .A(n18966), .B(n18971), .Z(n18792) );
  XNOR U19063 ( .A(n18972), .B(n18810), .Z(n18971) );
  ANDN U19064 ( .B(n18973), .A(n18974), .Z(n18810) );
  NOR U19065 ( .A(n18975), .B(n18976), .Z(n18972) );
  XNOR U19066 ( .A(n18808), .B(n18977), .Z(n18966) );
  XNOR U19067 ( .A(n18978), .B(n18979), .Z(n18977) );
  NAND U19068 ( .A(n18980), .B(n18981), .Z(n18979) );
  XOR U19069 ( .A(n18808), .B(n18982), .Z(n18900) );
  XNOR U19070 ( .A(n18968), .B(n18983), .Z(n18982) );
  NANDN U19071 ( .A(n18984), .B(n18985), .Z(n18983) );
  OR U19072 ( .A(n18986), .B(n18987), .Z(n18968) );
  XOR U19073 ( .A(n18988), .B(n18978), .Z(n18808) );
  OR U19074 ( .A(n18989), .B(n18990), .Z(n18978) );
  ANDN U19075 ( .B(n18991), .A(n18992), .Z(n18988) );
  XNOR U19076 ( .A(n18993), .B(n18994), .Z(n17635) );
  XNOR U19077 ( .A(n15492), .B(n15485), .Z(n16530) );
  XOR U19078 ( .A(n18784), .B(n18995), .Z(n15485) );
  XNOR U19079 ( .A(n18795), .B(n18783), .Z(n18995) );
  IV U19080 ( .A(n18902), .Z(n18783) );
  XOR U19081 ( .A(n18909), .B(n18996), .Z(n18902) );
  XNOR U19082 ( .A(n18906), .B(n18997), .Z(n18996) );
  NANDN U19083 ( .A(n18998), .B(n18865), .Z(n18997) );
  OR U19084 ( .A(n18999), .B(n18867), .Z(n18906) );
  XNOR U19085 ( .A(n18908), .B(n18865), .Z(n18867) );
  IV U19086 ( .A(n18786), .Z(n18795) );
  XOR U19087 ( .A(n18903), .B(n18774), .Z(n18786) );
  XOR U19088 ( .A(n18855), .B(n19000), .Z(n18774) );
  XNOR U19089 ( .A(n19001), .B(n19002), .Z(n19000) );
  NANDN U19090 ( .A(n19003), .B(n19004), .Z(n19002) );
  XOR U19091 ( .A(n18909), .B(n19005), .Z(n18903) );
  XOR U19092 ( .A(n19006), .B(n18858), .Z(n19005) );
  OR U19093 ( .A(n19007), .B(n19008), .Z(n18858) );
  ANDN U19094 ( .B(n19009), .A(n19010), .Z(n19006) );
  XOR U19095 ( .A(n19011), .B(n18911), .Z(n18909) );
  OR U19096 ( .A(n19012), .B(n19013), .Z(n18911) );
  ANDN U19097 ( .B(n19014), .A(n19015), .Z(n19011) );
  XNOR U19098 ( .A(n18801), .B(n19016), .Z(n18784) );
  XNOR U19099 ( .A(n19001), .B(n19017), .Z(n19016) );
  NANDN U19100 ( .A(n19018), .B(n18861), .Z(n19017) );
  OR U19101 ( .A(n19008), .B(n19019), .Z(n19001) );
  XNOR U19102 ( .A(n18861), .B(n19004), .Z(n19008) );
  XNOR U19103 ( .A(n18855), .B(n19020), .Z(n18801) );
  XNOR U19104 ( .A(n19021), .B(n19022), .Z(n19020) );
  NAND U19105 ( .A(n19023), .B(n18913), .Z(n19022) );
  XOR U19106 ( .A(n19024), .B(n19021), .Z(n18855) );
  NANDN U19107 ( .A(n19013), .B(n19025), .Z(n19021) );
  XOR U19108 ( .A(n19015), .B(n18913), .Z(n19013) );
  XOR U19109 ( .A(n19004), .B(n18865), .Z(n18913) );
  XOR U19110 ( .A(n19026), .B(n19027), .Z(n18865) );
  NANDN U19111 ( .A(n19028), .B(n19029), .Z(n19027) );
  IV U19112 ( .A(n19010), .Z(n19004) );
  XNOR U19113 ( .A(n19030), .B(n19031), .Z(n19010) );
  NANDN U19114 ( .A(n19028), .B(n19032), .Z(n19031) );
  ANDN U19115 ( .B(n19033), .A(n19015), .Z(n19024) );
  XNOR U19116 ( .A(n18908), .B(n18861), .Z(n19015) );
  XNOR U19117 ( .A(n19034), .B(n19030), .Z(n18861) );
  NANDN U19118 ( .A(n19035), .B(n19036), .Z(n19030) );
  XOR U19119 ( .A(n19032), .B(n19037), .Z(n19036) );
  ANDN U19120 ( .B(n19037), .A(n19038), .Z(n19034) );
  XNOR U19121 ( .A(n19039), .B(n19026), .Z(n18908) );
  NANDN U19122 ( .A(n19035), .B(n19040), .Z(n19026) );
  XOR U19123 ( .A(n19041), .B(n19029), .Z(n19040) );
  XNOR U19124 ( .A(n19042), .B(n19043), .Z(n19028) );
  XOR U19125 ( .A(n19044), .B(n19045), .Z(n19043) );
  XNOR U19126 ( .A(n19046), .B(n19047), .Z(n19042) );
  XNOR U19127 ( .A(n19048), .B(n19049), .Z(n19047) );
  ANDN U19128 ( .B(n19041), .A(n19045), .Z(n19048) );
  ANDN U19129 ( .B(n19041), .A(n19038), .Z(n19039) );
  XNOR U19130 ( .A(n19044), .B(n19050), .Z(n19038) );
  XOR U19131 ( .A(n19051), .B(n19049), .Z(n19050) );
  NAND U19132 ( .A(n19052), .B(n19053), .Z(n19049) );
  XNOR U19133 ( .A(n19046), .B(n19029), .Z(n19053) );
  IV U19134 ( .A(n19041), .Z(n19046) );
  XNOR U19135 ( .A(n19032), .B(n19045), .Z(n19052) );
  IV U19136 ( .A(n19037), .Z(n19045) );
  XOR U19137 ( .A(n19054), .B(n19055), .Z(n19037) );
  XNOR U19138 ( .A(n19056), .B(n19057), .Z(n19055) );
  XNOR U19139 ( .A(n19058), .B(n19059), .Z(n19054) );
  ANDN U19140 ( .B(n18907), .A(n19060), .Z(n19058) );
  AND U19141 ( .A(n19029), .B(n19032), .Z(n19051) );
  XNOR U19142 ( .A(n19029), .B(n19032), .Z(n19044) );
  XNOR U19143 ( .A(n19061), .B(n19062), .Z(n19032) );
  XNOR U19144 ( .A(n19063), .B(n19057), .Z(n19062) );
  XOR U19145 ( .A(n19064), .B(n19065), .Z(n19061) );
  XNOR U19146 ( .A(n19066), .B(n19059), .Z(n19065) );
  OR U19147 ( .A(n18868), .B(n18999), .Z(n19059) );
  XNOR U19148 ( .A(n18907), .B(n19067), .Z(n18999) );
  XNOR U19149 ( .A(n19060), .B(n18866), .Z(n18868) );
  ANDN U19150 ( .B(n19068), .A(n18998), .Z(n19066) );
  XNOR U19151 ( .A(n19069), .B(n19070), .Z(n19029) );
  XNOR U19152 ( .A(n19057), .B(n19071), .Z(n19070) );
  XOR U19153 ( .A(n19018), .B(n19064), .Z(n19071) );
  XNOR U19154 ( .A(n18907), .B(n19060), .Z(n19057) );
  XNOR U19155 ( .A(n19072), .B(n19073), .Z(n19069) );
  XNOR U19156 ( .A(n19074), .B(n19075), .Z(n19073) );
  ANDN U19157 ( .B(n19009), .A(n19003), .Z(n19074) );
  XNOR U19158 ( .A(n19076), .B(n19077), .Z(n19041) );
  XNOR U19159 ( .A(n19063), .B(n19078), .Z(n19077) );
  XNOR U19160 ( .A(n19003), .B(n19056), .Z(n19078) );
  XOR U19161 ( .A(n19064), .B(n19079), .Z(n19056) );
  XNOR U19162 ( .A(n19080), .B(n19081), .Z(n19079) );
  NAND U19163 ( .A(n18914), .B(n19023), .Z(n19081) );
  XNOR U19164 ( .A(n19082), .B(n19080), .Z(n19064) );
  NANDN U19165 ( .A(n19012), .B(n19025), .Z(n19080) );
  XOR U19166 ( .A(n19033), .B(n19023), .Z(n19025) );
  XNOR U19167 ( .A(n19083), .B(n18866), .Z(n19023) );
  XNOR U19168 ( .A(n19014), .B(n18914), .Z(n19012) );
  XOR U19169 ( .A(n19009), .B(n19067), .Z(n18914) );
  AND U19170 ( .A(n19033), .B(n19014), .Z(n19082) );
  XNOR U19171 ( .A(n18860), .B(n18907), .Z(n19014) );
  XNOR U19172 ( .A(n19084), .B(n19085), .Z(n18907) );
  XNOR U19173 ( .A(n19086), .B(n19087), .Z(n19085) );
  XOR U19174 ( .A(n19067), .B(n19068), .Z(n19063) );
  IV U19175 ( .A(n18866), .Z(n19068) );
  XOR U19176 ( .A(n19088), .B(n19089), .Z(n18866) );
  XNOR U19177 ( .A(n19090), .B(n19087), .Z(n19089) );
  IV U19178 ( .A(n18998), .Z(n19067) );
  XOR U19179 ( .A(n19087), .B(n19091), .Z(n18998) );
  XNOR U19180 ( .A(n19009), .B(n19092), .Z(n19076) );
  XNOR U19181 ( .A(n19093), .B(n19075), .Z(n19092) );
  OR U19182 ( .A(n19019), .B(n19007), .Z(n19075) );
  XNOR U19183 ( .A(n19072), .B(n19009), .Z(n19007) );
  XOR U19184 ( .A(n19018), .B(n19083), .Z(n19019) );
  IV U19185 ( .A(n19003), .Z(n19083) );
  XOR U19186 ( .A(n18799), .B(n19094), .Z(n19003) );
  XNOR U19187 ( .A(n19090), .B(n19084), .Z(n19094) );
  XOR U19188 ( .A(n19095), .B(n19096), .Z(n19084) );
  XNOR U19189 ( .A(n19097), .B(n18229), .Z(n19096) );
  XOR U19190 ( .A(key[450]), .B(n19098), .Z(n19095) );
  ANDN U19191 ( .B(n19099), .A(n18860), .Z(n19093) );
  XOR U19192 ( .A(n19100), .B(n19101), .Z(n19009) );
  XNOR U19193 ( .A(n19102), .B(n19103), .Z(n19101) );
  XOR U19194 ( .A(n19072), .B(n19086), .Z(n19100) );
  XOR U19195 ( .A(n19104), .B(n19105), .Z(n19086) );
  XNOR U19196 ( .A(n19090), .B(n19106), .Z(n19105) );
  XNOR U19197 ( .A(n19107), .B(n19108), .Z(n19106) );
  XOR U19198 ( .A(n19109), .B(n19110), .Z(n19090) );
  XOR U19199 ( .A(n18241), .B(n19111), .Z(n19110) );
  XOR U19200 ( .A(key[449]), .B(n19112), .Z(n19109) );
  XOR U19201 ( .A(n18196), .B(n19113), .Z(n19104) );
  XNOR U19202 ( .A(key[451]), .B(n19114), .Z(n19113) );
  XOR U19203 ( .A(n19099), .B(n18799), .Z(n19033) );
  IV U19204 ( .A(n19060), .Z(n18799) );
  XOR U19205 ( .A(n19088), .B(n19115), .Z(n19060) );
  XOR U19206 ( .A(n19087), .B(n19103), .Z(n19115) );
  XNOR U19207 ( .A(n19116), .B(n19117), .Z(n19103) );
  XNOR U19208 ( .A(n19118), .B(n19119), .Z(n19117) );
  XNOR U19209 ( .A(key[455]), .B(n19120), .Z(n19116) );
  IV U19210 ( .A(n19018), .Z(n19099) );
  XOR U19211 ( .A(n19088), .B(n19121), .Z(n19018) );
  XOR U19212 ( .A(n19087), .B(n19102), .Z(n19121) );
  XNOR U19213 ( .A(n19122), .B(n19123), .Z(n19102) );
  XOR U19214 ( .A(n19124), .B(n19125), .Z(n19123) );
  XNOR U19215 ( .A(n19126), .B(n19127), .Z(n19122) );
  XNOR U19216 ( .A(key[452]), .B(n19128), .Z(n19127) );
  XOR U19217 ( .A(n19129), .B(n19130), .Z(n19087) );
  XNOR U19218 ( .A(n19131), .B(n18860), .Z(n19130) );
  IV U19219 ( .A(n19072), .Z(n18860) );
  XOR U19220 ( .A(n19132), .B(n19133), .Z(n19072) );
  XOR U19221 ( .A(n19134), .B(n18234), .Z(n19133) );
  XNOR U19222 ( .A(key[448]), .B(n19135), .Z(n19132) );
  XOR U19223 ( .A(n19136), .B(n19137), .Z(n19129) );
  XNOR U19224 ( .A(key[454]), .B(n19138), .Z(n19137) );
  IV U19225 ( .A(n19091), .Z(n19088) );
  XOR U19226 ( .A(n19139), .B(n19140), .Z(n19091) );
  XOR U19227 ( .A(n19141), .B(n19142), .Z(n19140) );
  XNOR U19228 ( .A(key[453]), .B(n19143), .Z(n19139) );
  XOR U19229 ( .A(n18848), .B(n19144), .Z(n15492) );
  XNOR U19230 ( .A(n18802), .B(n18850), .Z(n19144) );
  XOR U19231 ( .A(n19145), .B(n19146), .Z(n18850) );
  XOR U19232 ( .A(n19147), .B(n19148), .Z(n19146) );
  NANDN U19233 ( .A(n19149), .B(n18884), .Z(n19148) );
  XOR U19234 ( .A(n18901), .B(n18918), .Z(n18802) );
  XOR U19235 ( .A(n18880), .B(n19150), .Z(n18918) );
  XNOR U19236 ( .A(n19151), .B(n19152), .Z(n19150) );
  NANDN U19237 ( .A(n19153), .B(n19154), .Z(n19152) );
  XNOR U19238 ( .A(n18919), .B(n19155), .Z(n18848) );
  XNOR U19239 ( .A(n19151), .B(n19156), .Z(n19155) );
  NANDN U19240 ( .A(n19157), .B(n18879), .Z(n19156) );
  OR U19241 ( .A(n19158), .B(n19159), .Z(n19151) );
  XNOR U19242 ( .A(n18880), .B(n19160), .Z(n18919) );
  XNOR U19243 ( .A(n19161), .B(n19162), .Z(n19160) );
  NAND U19244 ( .A(n19163), .B(n19164), .Z(n19162) );
  XOR U19245 ( .A(n19165), .B(n19161), .Z(n18880) );
  NANDN U19246 ( .A(n19166), .B(n19167), .Z(n19161) );
  ANDN U19247 ( .B(n19168), .A(n19169), .Z(n19165) );
  XNOR U19248 ( .A(n16505), .B(n16538), .Z(n15457) );
  IV U19249 ( .A(n18870), .Z(n16538) );
  XNOR U19250 ( .A(n18901), .B(n18873), .Z(n18870) );
  XNOR U19251 ( .A(n18874), .B(n19170), .Z(n18873) );
  XNOR U19252 ( .A(n19171), .B(n19147), .Z(n19170) );
  XNOR U19253 ( .A(n18925), .B(n18884), .Z(n18922) );
  ANDN U19254 ( .B(n19173), .A(n18925), .Z(n19171) );
  XNOR U19255 ( .A(n19145), .B(n19174), .Z(n18874) );
  XNOR U19256 ( .A(n19175), .B(n19176), .Z(n19174) );
  NAND U19257 ( .A(n19164), .B(n19177), .Z(n19176) );
  XOR U19258 ( .A(n19145), .B(n19178), .Z(n18901) );
  XOR U19259 ( .A(n19179), .B(n18876), .Z(n19178) );
  OR U19260 ( .A(n19180), .B(n19158), .Z(n18876) );
  XNOR U19261 ( .A(n18879), .B(n19154), .Z(n19158) );
  ANDN U19262 ( .B(n19181), .A(n19182), .Z(n19179) );
  XOR U19263 ( .A(n19183), .B(n19175), .Z(n19145) );
  OR U19264 ( .A(n19166), .B(n19184), .Z(n19175) );
  XNOR U19265 ( .A(n19185), .B(n19164), .Z(n19166) );
  XOR U19266 ( .A(n19154), .B(n18884), .Z(n19164) );
  XOR U19267 ( .A(n19186), .B(n19187), .Z(n18884) );
  NANDN U19268 ( .A(n19188), .B(n19189), .Z(n19187) );
  IV U19269 ( .A(n19182), .Z(n19154) );
  XNOR U19270 ( .A(n19190), .B(n19191), .Z(n19182) );
  NANDN U19271 ( .A(n19188), .B(n19192), .Z(n19191) );
  ANDN U19272 ( .B(n19185), .A(n19193), .Z(n19183) );
  IV U19273 ( .A(n19169), .Z(n19185) );
  XOR U19274 ( .A(n18925), .B(n18879), .Z(n19169) );
  XNOR U19275 ( .A(n19194), .B(n19190), .Z(n18879) );
  NANDN U19276 ( .A(n19195), .B(n19196), .Z(n19190) );
  XOR U19277 ( .A(n19192), .B(n19197), .Z(n19196) );
  ANDN U19278 ( .B(n19197), .A(n19198), .Z(n19194) );
  XOR U19279 ( .A(n19199), .B(n19186), .Z(n18925) );
  NANDN U19280 ( .A(n19195), .B(n19200), .Z(n19186) );
  XOR U19281 ( .A(n19201), .B(n19189), .Z(n19200) );
  XNOR U19282 ( .A(n19202), .B(n19203), .Z(n19188) );
  XOR U19283 ( .A(n19204), .B(n19205), .Z(n19203) );
  XNOR U19284 ( .A(n19206), .B(n19207), .Z(n19202) );
  XNOR U19285 ( .A(n19208), .B(n19209), .Z(n19207) );
  ANDN U19286 ( .B(n19201), .A(n19205), .Z(n19208) );
  ANDN U19287 ( .B(n19201), .A(n19198), .Z(n19199) );
  XNOR U19288 ( .A(n19204), .B(n19210), .Z(n19198) );
  XOR U19289 ( .A(n19211), .B(n19209), .Z(n19210) );
  NAND U19290 ( .A(n19212), .B(n19213), .Z(n19209) );
  XNOR U19291 ( .A(n19206), .B(n19189), .Z(n19213) );
  IV U19292 ( .A(n19201), .Z(n19206) );
  XNOR U19293 ( .A(n19192), .B(n19205), .Z(n19212) );
  IV U19294 ( .A(n19197), .Z(n19205) );
  XOR U19295 ( .A(n19214), .B(n19215), .Z(n19197) );
  XNOR U19296 ( .A(n19216), .B(n19217), .Z(n19215) );
  XNOR U19297 ( .A(n19218), .B(n19219), .Z(n19214) );
  ANDN U19298 ( .B(n19173), .A(n18924), .Z(n19218) );
  AND U19299 ( .A(n19189), .B(n19192), .Z(n19211) );
  XNOR U19300 ( .A(n19189), .B(n19192), .Z(n19204) );
  XNOR U19301 ( .A(n19220), .B(n19221), .Z(n19192) );
  XNOR U19302 ( .A(n19222), .B(n19217), .Z(n19221) );
  XOR U19303 ( .A(n19223), .B(n19224), .Z(n19220) );
  XNOR U19304 ( .A(n19225), .B(n19219), .Z(n19224) );
  OR U19305 ( .A(n18923), .B(n19172), .Z(n19219) );
  XNOR U19306 ( .A(n19173), .B(n19226), .Z(n19172) );
  XNOR U19307 ( .A(n18924), .B(n18885), .Z(n18923) );
  ANDN U19308 ( .B(n19227), .A(n19149), .Z(n19225) );
  XNOR U19309 ( .A(n19228), .B(n19229), .Z(n19189) );
  XNOR U19310 ( .A(n19217), .B(n19230), .Z(n19229) );
  XOR U19311 ( .A(n19157), .B(n19223), .Z(n19230) );
  XNOR U19312 ( .A(n19173), .B(n18924), .Z(n19217) );
  XNOR U19313 ( .A(n19231), .B(n19232), .Z(n19228) );
  XNOR U19314 ( .A(n19233), .B(n19234), .Z(n19232) );
  ANDN U19315 ( .B(n19181), .A(n19153), .Z(n19233) );
  XNOR U19316 ( .A(n19235), .B(n19236), .Z(n19201) );
  XNOR U19317 ( .A(n19222), .B(n19237), .Z(n19236) );
  XNOR U19318 ( .A(n19153), .B(n19216), .Z(n19237) );
  XOR U19319 ( .A(n19223), .B(n19238), .Z(n19216) );
  XNOR U19320 ( .A(n19239), .B(n19240), .Z(n19238) );
  NAND U19321 ( .A(n19177), .B(n19163), .Z(n19240) );
  XNOR U19322 ( .A(n19241), .B(n19239), .Z(n19223) );
  NANDN U19323 ( .A(n19184), .B(n19167), .Z(n19239) );
  XOR U19324 ( .A(n19168), .B(n19163), .Z(n19167) );
  XNOR U19325 ( .A(n19242), .B(n18885), .Z(n19163) );
  XOR U19326 ( .A(n19193), .B(n19177), .Z(n19184) );
  XOR U19327 ( .A(n19181), .B(n19226), .Z(n19177) );
  ANDN U19328 ( .B(n19168), .A(n19193), .Z(n19241) );
  XNOR U19329 ( .A(n19231), .B(n19173), .Z(n19193) );
  XNOR U19330 ( .A(n19243), .B(n19244), .Z(n19173) );
  XNOR U19331 ( .A(n19245), .B(n19246), .Z(n19244) );
  XOR U19332 ( .A(n19247), .B(n19248), .Z(n19168) );
  XOR U19333 ( .A(n19226), .B(n19227), .Z(n19222) );
  IV U19334 ( .A(n18885), .Z(n19227) );
  XOR U19335 ( .A(n19249), .B(n19250), .Z(n18885) );
  XNOR U19336 ( .A(n19251), .B(n19246), .Z(n19250) );
  IV U19337 ( .A(n19149), .Z(n19226) );
  XOR U19338 ( .A(n19246), .B(n19252), .Z(n19149) );
  XNOR U19339 ( .A(n19181), .B(n19253), .Z(n19235) );
  XNOR U19340 ( .A(n19254), .B(n19234), .Z(n19253) );
  OR U19341 ( .A(n19159), .B(n19180), .Z(n19234) );
  XNOR U19342 ( .A(n19231), .B(n19181), .Z(n19180) );
  XOR U19343 ( .A(n19157), .B(n19242), .Z(n19159) );
  IV U19344 ( .A(n19153), .Z(n19242) );
  XOR U19345 ( .A(n19248), .B(n19255), .Z(n19153) );
  XNOR U19346 ( .A(n19251), .B(n19243), .Z(n19255) );
  XOR U19347 ( .A(n19256), .B(n19257), .Z(n19243) );
  XOR U19348 ( .A(n18645), .B(n18640), .Z(n19257) );
  XOR U19349 ( .A(n19258), .B(n19259), .Z(n19256) );
  XNOR U19350 ( .A(key[442]), .B(n19260), .Z(n19259) );
  IV U19351 ( .A(n18924), .Z(n19248) );
  XOR U19352 ( .A(n19249), .B(n19261), .Z(n18924) );
  XOR U19353 ( .A(n19246), .B(n19262), .Z(n19261) );
  ANDN U19354 ( .B(n19247), .A(n18878), .Z(n19254) );
  IV U19355 ( .A(n19157), .Z(n19247) );
  XOR U19356 ( .A(n19249), .B(n19263), .Z(n19157) );
  XOR U19357 ( .A(n19246), .B(n19264), .Z(n19263) );
  XOR U19358 ( .A(n19265), .B(n19266), .Z(n19246) );
  XNOR U19359 ( .A(n19267), .B(n18878), .Z(n19266) );
  IV U19360 ( .A(n19231), .Z(n18878) );
  XOR U19361 ( .A(n19268), .B(n19269), .Z(n19265) );
  XNOR U19362 ( .A(key[446]), .B(n18617), .Z(n19269) );
  IV U19363 ( .A(n19252), .Z(n19249) );
  XOR U19364 ( .A(n19270), .B(n19271), .Z(n19252) );
  XOR U19365 ( .A(n18634), .B(n19272), .Z(n19271) );
  XOR U19366 ( .A(n19273), .B(n19274), .Z(n19270) );
  XNOR U19367 ( .A(key[445]), .B(n19275), .Z(n19274) );
  XOR U19368 ( .A(n19276), .B(n19277), .Z(n19181) );
  XNOR U19369 ( .A(n19264), .B(n19262), .Z(n19277) );
  XNOR U19370 ( .A(n19278), .B(n19279), .Z(n19262) );
  XOR U19371 ( .A(n18655), .B(n19280), .Z(n19279) );
  XNOR U19372 ( .A(key[447]), .B(n19281), .Z(n19278) );
  XNOR U19373 ( .A(n19282), .B(n19283), .Z(n19264) );
  XNOR U19374 ( .A(n19284), .B(n19285), .Z(n19282) );
  XOR U19375 ( .A(key[444]), .B(n19286), .Z(n19285) );
  XOR U19376 ( .A(n19231), .B(n19245), .Z(n19276) );
  XOR U19377 ( .A(n19287), .B(n19288), .Z(n19245) );
  XNOR U19378 ( .A(n19251), .B(n19289), .Z(n19288) );
  XNOR U19379 ( .A(n19290), .B(n19291), .Z(n19289) );
  XOR U19380 ( .A(n19292), .B(n19293), .Z(n19251) );
  XNOR U19381 ( .A(n18626), .B(n19294), .Z(n19293) );
  XNOR U19382 ( .A(n19295), .B(n19296), .Z(n19292) );
  XNOR U19383 ( .A(key[441]), .B(n19297), .Z(n19296) );
  XNOR U19384 ( .A(n19298), .B(n19299), .Z(n19287) );
  XNOR U19385 ( .A(key[443]), .B(n18630), .Z(n19299) );
  XOR U19386 ( .A(n19300), .B(n19301), .Z(n19231) );
  XNOR U19387 ( .A(n19302), .B(n19303), .Z(n19301) );
  XNOR U19388 ( .A(n19304), .B(n19305), .Z(n19300) );
  XNOR U19389 ( .A(key[440]), .B(n19306), .Z(n19305) );
  IV U19390 ( .A(n15495), .Z(n16505) );
  XOR U19391 ( .A(n18887), .B(n18806), .Z(n15495) );
  XNOR U19392 ( .A(n18840), .B(n19307), .Z(n18806) );
  XOR U19393 ( .A(n19308), .B(n18963), .Z(n19307) );
  XNOR U19394 ( .A(n18975), .B(n18812), .Z(n18973) );
  ANDN U19395 ( .B(n19310), .A(n18975), .Z(n19308) );
  XOR U19396 ( .A(n18961), .B(n19311), .Z(n18840) );
  XNOR U19397 ( .A(n19312), .B(n19313), .Z(n19311) );
  NAND U19398 ( .A(n18981), .B(n19314), .Z(n19313) );
  XOR U19399 ( .A(n19316), .B(n18842), .Z(n19315) );
  OR U19400 ( .A(n18986), .B(n19317), .Z(n18842) );
  XNOR U19401 ( .A(n18844), .B(n18984), .Z(n18986) );
  NOR U19402 ( .A(n19318), .B(n18984), .Z(n19316) );
  XNOR U19403 ( .A(n19319), .B(n19312), .Z(n18961) );
  OR U19404 ( .A(n18989), .B(n19320), .Z(n19312) );
  XNOR U19405 ( .A(n18991), .B(n18981), .Z(n18989) );
  XNOR U19406 ( .A(n18984), .B(n18812), .Z(n18981) );
  XOR U19407 ( .A(n19321), .B(n19322), .Z(n18812) );
  NANDN U19408 ( .A(n19323), .B(n19324), .Z(n19322) );
  XNOR U19409 ( .A(n19325), .B(n19326), .Z(n18984) );
  OR U19410 ( .A(n19323), .B(n19327), .Z(n19326) );
  XOR U19411 ( .A(n18844), .B(n18975), .Z(n18991) );
  XOR U19412 ( .A(n19329), .B(n19321), .Z(n18975) );
  NANDN U19413 ( .A(n19330), .B(n19331), .Z(n19321) );
  ANDN U19414 ( .B(n19332), .A(n19333), .Z(n19329) );
  NANDN U19415 ( .A(n19330), .B(n19335), .Z(n19325) );
  XOR U19416 ( .A(n19336), .B(n19323), .Z(n19330) );
  XNOR U19417 ( .A(n19337), .B(n19338), .Z(n19323) );
  XOR U19418 ( .A(n19339), .B(n19332), .Z(n19338) );
  XNOR U19419 ( .A(n19340), .B(n19341), .Z(n19337) );
  XNOR U19420 ( .A(n19342), .B(n19343), .Z(n19341) );
  ANDN U19421 ( .B(n19332), .A(n19344), .Z(n19342) );
  IV U19422 ( .A(n19345), .Z(n19332) );
  ANDN U19423 ( .B(n19336), .A(n19344), .Z(n19334) );
  IV U19424 ( .A(n19340), .Z(n19344) );
  IV U19425 ( .A(n19333), .Z(n19336) );
  XNOR U19426 ( .A(n19339), .B(n19346), .Z(n19333) );
  XOR U19427 ( .A(n19347), .B(n19343), .Z(n19346) );
  NAND U19428 ( .A(n19335), .B(n19331), .Z(n19343) );
  XNOR U19429 ( .A(n19324), .B(n19345), .Z(n19331) );
  XOR U19430 ( .A(n19348), .B(n19349), .Z(n19345) );
  XOR U19431 ( .A(n19350), .B(n19351), .Z(n19349) );
  XOR U19432 ( .A(n19352), .B(n19353), .Z(n19351) );
  XOR U19433 ( .A(n18985), .B(n19354), .Z(n19348) );
  XNOR U19434 ( .A(n19355), .B(n19356), .Z(n19354) );
  ANDN U19435 ( .B(n18970), .A(n18845), .Z(n19355) );
  XNOR U19436 ( .A(n19340), .B(n19327), .Z(n19335) );
  XOR U19437 ( .A(n19357), .B(n19358), .Z(n19340) );
  XNOR U19438 ( .A(n19359), .B(n19353), .Z(n19358) );
  XOR U19439 ( .A(n19360), .B(n19361), .Z(n19353) );
  XNOR U19440 ( .A(n19362), .B(n19363), .Z(n19361) );
  NAND U19441 ( .A(n19314), .B(n18980), .Z(n19363) );
  XNOR U19442 ( .A(n19364), .B(n19365), .Z(n19357) );
  ANDN U19443 ( .B(n19310), .A(n18976), .Z(n19364) );
  ANDN U19444 ( .B(n19324), .A(n19327), .Z(n19347) );
  XOR U19445 ( .A(n19327), .B(n19324), .Z(n19339) );
  XNOR U19446 ( .A(n19366), .B(n19367), .Z(n19324) );
  XNOR U19447 ( .A(n19360), .B(n19368), .Z(n19367) );
  XNOR U19448 ( .A(n18970), .B(n19359), .Z(n19368) );
  XNOR U19449 ( .A(n19369), .B(n19370), .Z(n19366) );
  XNOR U19450 ( .A(n19371), .B(n19356), .Z(n19370) );
  OR U19451 ( .A(n18987), .B(n19317), .Z(n19356) );
  XNOR U19452 ( .A(n19369), .B(n19352), .Z(n19317) );
  XNOR U19453 ( .A(n18970), .B(n18985), .Z(n18987) );
  ANDN U19454 ( .B(n18985), .A(n19318), .Z(n19371) );
  IV U19455 ( .A(n19352), .Z(n19318) );
  XOR U19456 ( .A(n19372), .B(n19373), .Z(n19327) );
  XOR U19457 ( .A(n19360), .B(n19350), .Z(n19373) );
  XOR U19458 ( .A(n19374), .B(n18965), .Z(n19350) );
  XOR U19459 ( .A(n19375), .B(n19362), .Z(n19360) );
  OR U19460 ( .A(n19320), .B(n18990), .Z(n19362) );
  XOR U19461 ( .A(n18992), .B(n18980), .Z(n18990) );
  XOR U19462 ( .A(n19374), .B(n18985), .Z(n18980) );
  XOR U19463 ( .A(n19376), .B(n19377), .Z(n18985) );
  XNOR U19464 ( .A(n18976), .B(n19378), .Z(n19377) );
  XNOR U19465 ( .A(n19328), .B(n19314), .Z(n19320) );
  XNOR U19466 ( .A(n18965), .B(n19352), .Z(n19314) );
  XOR U19467 ( .A(n19379), .B(n19380), .Z(n19352) );
  XNOR U19468 ( .A(n19381), .B(n19382), .Z(n19380) );
  XOR U19469 ( .A(n19369), .B(n19383), .Z(n19379) );
  ANDN U19470 ( .B(n19328), .A(n18992), .Z(n19375) );
  XOR U19471 ( .A(n18976), .B(n18970), .Z(n18992) );
  XOR U19472 ( .A(n19381), .B(n19384), .Z(n18970) );
  XOR U19473 ( .A(n19385), .B(n19386), .Z(n19384) );
  XOR U19474 ( .A(n19387), .B(n19388), .Z(n19381) );
  XNOR U19475 ( .A(n19389), .B(n19390), .Z(n19388) );
  XOR U19476 ( .A(key[404]), .B(n19391), .Z(n19387) );
  XOR U19477 ( .A(n19359), .B(n19392), .Z(n19372) );
  XNOR U19478 ( .A(n19393), .B(n19365), .Z(n19392) );
  OR U19479 ( .A(n19309), .B(n18974), .Z(n19365) );
  XOR U19480 ( .A(n18976), .B(n19374), .Z(n18974) );
  XNOR U19481 ( .A(n19310), .B(n19395), .Z(n19309) );
  ANDN U19482 ( .B(n19374), .A(n18965), .Z(n19393) );
  XOR U19483 ( .A(n19394), .B(n19386), .Z(n18965) );
  IV U19484 ( .A(n18813), .Z(n19374) );
  XNOR U19485 ( .A(n19378), .B(n19395), .Z(n18813) );
  XOR U19486 ( .A(n18976), .B(n19310), .Z(n19359) );
  XNOR U19487 ( .A(n19383), .B(n19395), .Z(n18976) );
  XNOR U19488 ( .A(n19394), .B(n19386), .Z(n19395) );
  IV U19489 ( .A(n19385), .Z(n19394) );
  XNOR U19490 ( .A(n19396), .B(n19397), .Z(n19385) );
  XOR U19491 ( .A(n19398), .B(n19399), .Z(n19397) );
  XOR U19492 ( .A(key[405]), .B(n19400), .Z(n19396) );
  XOR U19493 ( .A(n19401), .B(n19402), .Z(n19383) );
  XNOR U19494 ( .A(n19403), .B(n19404), .Z(n19402) );
  XNOR U19495 ( .A(key[407]), .B(n19405), .Z(n19401) );
  XOR U19496 ( .A(n19369), .B(n19310), .Z(n19328) );
  XNOR U19497 ( .A(n19382), .B(n19406), .Z(n19310) );
  XNOR U19498 ( .A(n19386), .B(n19376), .Z(n19406) );
  XOR U19499 ( .A(n19407), .B(n19408), .Z(n19376) );
  XNOR U19500 ( .A(n19409), .B(n19410), .Z(n19408) );
  XOR U19501 ( .A(key[402]), .B(n18510), .Z(n19407) );
  XOR U19502 ( .A(n19411), .B(n19412), .Z(n19386) );
  XOR U19503 ( .A(n19413), .B(n18845), .Z(n19412) );
  IV U19504 ( .A(n19369), .Z(n18845) );
  XOR U19505 ( .A(n19414), .B(n19415), .Z(n19411) );
  XNOR U19506 ( .A(key[406]), .B(n19416), .Z(n19415) );
  XOR U19507 ( .A(n19417), .B(n19418), .Z(n19382) );
  XNOR U19508 ( .A(n19378), .B(n19419), .Z(n19418) );
  XOR U19509 ( .A(n19420), .B(n19421), .Z(n19419) );
  XOR U19510 ( .A(n19422), .B(n19423), .Z(n19378) );
  XNOR U19511 ( .A(n18517), .B(n19424), .Z(n19423) );
  XOR U19512 ( .A(key[401]), .B(n19425), .Z(n19422) );
  XOR U19513 ( .A(n18469), .B(n19426), .Z(n19417) );
  XOR U19514 ( .A(key[403]), .B(n19427), .Z(n19426) );
  XOR U19515 ( .A(n19428), .B(n19429), .Z(n19369) );
  XNOR U19516 ( .A(n19430), .B(n18509), .Z(n19429) );
  XNOR U19517 ( .A(key[400]), .B(n19431), .Z(n19428) );
  XNOR U19518 ( .A(key[544]), .B(n16957), .Z(n18993) );
  XOR U19519 ( .A(n18816), .B(n18897), .Z(n16957) );
  XOR U19520 ( .A(n19433), .B(n18834), .Z(n19432) );
  OR U19521 ( .A(n19434), .B(n18953), .Z(n18834) );
  XNOR U19522 ( .A(n18836), .B(n18951), .Z(n18953) );
  NOR U19523 ( .A(n19435), .B(n18951), .Z(n19433) );
  XNOR U19524 ( .A(n18832), .B(n19436), .Z(n18816) );
  XOR U19525 ( .A(n19437), .B(n18930), .Z(n19436) );
  OR U19526 ( .A(n19438), .B(n18940), .Z(n18930) );
  XNOR U19527 ( .A(n19439), .B(n18822), .Z(n18940) );
  ANDN U19528 ( .B(n19440), .A(n18942), .Z(n19437) );
  IV U19529 ( .A(n19439), .Z(n18942) );
  XOR U19530 ( .A(n18928), .B(n19441), .Z(n18832) );
  XNOR U19531 ( .A(n19442), .B(n19443), .Z(n19441) );
  NAND U19532 ( .A(n18948), .B(n19444), .Z(n19443) );
  XNOR U19533 ( .A(n19445), .B(n19442), .Z(n18928) );
  NANDN U19534 ( .A(n18956), .B(n19446), .Z(n19442) );
  XOR U19535 ( .A(n18959), .B(n18948), .Z(n18956) );
  XNOR U19536 ( .A(n18951), .B(n18822), .Z(n18948) );
  XOR U19537 ( .A(n19447), .B(n19448), .Z(n18822) );
  NANDN U19538 ( .A(n19449), .B(n19450), .Z(n19448) );
  XNOR U19539 ( .A(n19451), .B(n19452), .Z(n18951) );
  OR U19540 ( .A(n19449), .B(n19453), .Z(n19452) );
  ANDN U19541 ( .B(n19454), .A(n18959), .Z(n19445) );
  XOR U19542 ( .A(n18836), .B(n19439), .Z(n18959) );
  XNOR U19543 ( .A(n19455), .B(n19447), .Z(n19439) );
  NANDN U19544 ( .A(n19456), .B(n19457), .Z(n19447) );
  ANDN U19545 ( .B(n19458), .A(n19459), .Z(n19455) );
  NANDN U19546 ( .A(n19456), .B(n19461), .Z(n19451) );
  XOR U19547 ( .A(n19462), .B(n19449), .Z(n19456) );
  XNOR U19548 ( .A(n19463), .B(n19464), .Z(n19449) );
  XOR U19549 ( .A(n19465), .B(n19458), .Z(n19464) );
  XNOR U19550 ( .A(n19466), .B(n19467), .Z(n19463) );
  XNOR U19551 ( .A(n19468), .B(n19469), .Z(n19467) );
  ANDN U19552 ( .B(n19458), .A(n19470), .Z(n19468) );
  IV U19553 ( .A(n19471), .Z(n19458) );
  ANDN U19554 ( .B(n19462), .A(n19470), .Z(n19460) );
  IV U19555 ( .A(n19466), .Z(n19470) );
  IV U19556 ( .A(n19459), .Z(n19462) );
  XNOR U19557 ( .A(n19465), .B(n19472), .Z(n19459) );
  XOR U19558 ( .A(n19473), .B(n19469), .Z(n19472) );
  NAND U19559 ( .A(n19461), .B(n19457), .Z(n19469) );
  XNOR U19560 ( .A(n19450), .B(n19471), .Z(n19457) );
  XOR U19561 ( .A(n19474), .B(n19475), .Z(n19471) );
  XOR U19562 ( .A(n19476), .B(n19477), .Z(n19475) );
  XOR U19563 ( .A(n19478), .B(n19479), .Z(n19477) );
  XOR U19564 ( .A(n18952), .B(n19480), .Z(n19474) );
  XNOR U19565 ( .A(n19481), .B(n19482), .Z(n19480) );
  ANDN U19566 ( .B(n18937), .A(n18837), .Z(n19481) );
  XNOR U19567 ( .A(n19466), .B(n19453), .Z(n19461) );
  XOR U19568 ( .A(n19483), .B(n19484), .Z(n19466) );
  XNOR U19569 ( .A(n19485), .B(n19479), .Z(n19484) );
  XOR U19570 ( .A(n19486), .B(n19487), .Z(n19479) );
  XNOR U19571 ( .A(n19488), .B(n19489), .Z(n19487) );
  NAND U19572 ( .A(n19444), .B(n18947), .Z(n19489) );
  XNOR U19573 ( .A(n19490), .B(n19491), .Z(n19483) );
  ANDN U19574 ( .B(n19440), .A(n18943), .Z(n19490) );
  ANDN U19575 ( .B(n19450), .A(n19453), .Z(n19473) );
  XOR U19576 ( .A(n19453), .B(n19450), .Z(n19465) );
  XNOR U19577 ( .A(n19492), .B(n19493), .Z(n19450) );
  XNOR U19578 ( .A(n19486), .B(n19494), .Z(n19493) );
  XNOR U19579 ( .A(n18937), .B(n19485), .Z(n19494) );
  XNOR U19580 ( .A(n19495), .B(n19496), .Z(n19492) );
  XNOR U19581 ( .A(n19497), .B(n19482), .Z(n19496) );
  OR U19582 ( .A(n18954), .B(n19434), .Z(n19482) );
  XNOR U19583 ( .A(n19495), .B(n19478), .Z(n19434) );
  XNOR U19584 ( .A(n18937), .B(n18952), .Z(n18954) );
  ANDN U19585 ( .B(n18952), .A(n19435), .Z(n19497) );
  IV U19586 ( .A(n19478), .Z(n19435) );
  XOR U19587 ( .A(n19498), .B(n19499), .Z(n19453) );
  XOR U19588 ( .A(n19486), .B(n19476), .Z(n19499) );
  XOR U19589 ( .A(n19500), .B(n18932), .Z(n19476) );
  XOR U19590 ( .A(n19501), .B(n19488), .Z(n19486) );
  NANDN U19591 ( .A(n18957), .B(n19446), .Z(n19488) );
  XOR U19592 ( .A(n19454), .B(n19444), .Z(n19446) );
  XNOR U19593 ( .A(n18932), .B(n19478), .Z(n19444) );
  XOR U19594 ( .A(n19502), .B(n19503), .Z(n19478) );
  XNOR U19595 ( .A(n19504), .B(n19505), .Z(n19503) );
  XOR U19596 ( .A(n19495), .B(n19506), .Z(n19502) );
  XOR U19597 ( .A(n18958), .B(n18947), .Z(n18957) );
  XOR U19598 ( .A(n19500), .B(n18952), .Z(n18947) );
  XOR U19599 ( .A(n19507), .B(n19508), .Z(n18952) );
  XNOR U19600 ( .A(n18943), .B(n19509), .Z(n19508) );
  ANDN U19601 ( .B(n19454), .A(n18958), .Z(n19501) );
  XOR U19602 ( .A(n18943), .B(n18937), .Z(n18958) );
  XOR U19603 ( .A(n19504), .B(n19510), .Z(n18937) );
  XOR U19604 ( .A(n19511), .B(n19512), .Z(n19510) );
  XOR U19605 ( .A(n19513), .B(n19514), .Z(n19504) );
  XOR U19606 ( .A(n19515), .B(n19516), .Z(n19513) );
  XNOR U19607 ( .A(key[492]), .B(n19517), .Z(n19516) );
  XOR U19608 ( .A(n19485), .B(n19518), .Z(n19498) );
  XNOR U19609 ( .A(n19519), .B(n19491), .Z(n19518) );
  OR U19610 ( .A(n19438), .B(n18941), .Z(n19491) );
  XOR U19611 ( .A(n18943), .B(n19500), .Z(n18941) );
  XNOR U19612 ( .A(n19440), .B(n19521), .Z(n19438) );
  ANDN U19613 ( .B(n19500), .A(n18932), .Z(n19519) );
  XOR U19614 ( .A(n19520), .B(n19512), .Z(n18932) );
  IV U19615 ( .A(n18823), .Z(n19500) );
  XNOR U19616 ( .A(n19509), .B(n19521), .Z(n18823) );
  XOR U19617 ( .A(n18943), .B(n19440), .Z(n19485) );
  XNOR U19618 ( .A(n19506), .B(n19521), .Z(n18943) );
  XNOR U19619 ( .A(n19520), .B(n19512), .Z(n19521) );
  IV U19620 ( .A(n19511), .Z(n19520) );
  XNOR U19621 ( .A(n19522), .B(n19523), .Z(n19511) );
  XOR U19622 ( .A(n19524), .B(n19525), .Z(n19523) );
  XOR U19623 ( .A(n19526), .B(n19527), .Z(n19522) );
  XNOR U19624 ( .A(key[493]), .B(n19528), .Z(n19527) );
  XOR U19625 ( .A(n19529), .B(n19530), .Z(n19506) );
  XOR U19626 ( .A(n18382), .B(n19531), .Z(n19530) );
  XNOR U19627 ( .A(key[495]), .B(n19532), .Z(n19529) );
  XOR U19628 ( .A(n19495), .B(n19440), .Z(n19454) );
  XNOR U19629 ( .A(n19505), .B(n19533), .Z(n19440) );
  XNOR U19630 ( .A(n19512), .B(n19507), .Z(n19533) );
  XOR U19631 ( .A(n19534), .B(n19535), .Z(n19507) );
  XNOR U19632 ( .A(n19536), .B(n19537), .Z(n19535) );
  XOR U19633 ( .A(n18364), .B(n19538), .Z(n19534) );
  XNOR U19634 ( .A(key[490]), .B(n18371), .Z(n19538) );
  XOR U19635 ( .A(n19539), .B(n19540), .Z(n19512) );
  XNOR U19636 ( .A(n19541), .B(n18837), .Z(n19540) );
  IV U19637 ( .A(n19495), .Z(n18837) );
  XNOR U19638 ( .A(n18334), .B(n19542), .Z(n19539) );
  XNOR U19639 ( .A(key[494]), .B(n19543), .Z(n19542) );
  XOR U19640 ( .A(n19544), .B(n19545), .Z(n19505) );
  XNOR U19641 ( .A(n19509), .B(n19546), .Z(n19545) );
  XNOR U19642 ( .A(n18375), .B(n19547), .Z(n19546) );
  XOR U19643 ( .A(n19548), .B(n19549), .Z(n19509) );
  XNOR U19644 ( .A(n18374), .B(n18381), .Z(n19549) );
  XNOR U19645 ( .A(n19550), .B(n19551), .Z(n19548) );
  XNOR U19646 ( .A(key[489]), .B(n19552), .Z(n19551) );
  XNOR U19647 ( .A(n19553), .B(n19554), .Z(n19544) );
  XOR U19648 ( .A(key[491]), .B(n19555), .Z(n19554) );
  XOR U19649 ( .A(n19556), .B(n19557), .Z(n19495) );
  XNOR U19650 ( .A(n19558), .B(n19559), .Z(n19557) );
  XNOR U19651 ( .A(n18341), .B(n19560), .Z(n19556) );
  XNOR U19652 ( .A(key[488]), .B(n19561), .Z(n19560) );
  IV U19653 ( .A(n17649), .Z(n14428) );
  XNOR U19654 ( .A(n17604), .B(n17567), .Z(n19562) );
  XOR U19655 ( .A(n17667), .B(n17678), .Z(n17567) );
  XNOR U19656 ( .A(n17614), .B(n19563), .Z(n17678) );
  XNOR U19657 ( .A(n19564), .B(n19565), .Z(n19563) );
  NANDN U19658 ( .A(n19566), .B(n19567), .Z(n19565) );
  XNOR U19659 ( .A(n18663), .B(n19568), .Z(n17667) );
  XOR U19660 ( .A(n19569), .B(n17617), .Z(n19568) );
  OR U19661 ( .A(n19570), .B(n19571), .Z(n17617) );
  ANDN U19662 ( .B(n19567), .A(n19572), .Z(n19569) );
  XNOR U19663 ( .A(n19564), .B(n19574), .Z(n19573) );
  NANDN U19664 ( .A(n19575), .B(n17620), .Z(n19574) );
  OR U19665 ( .A(n19570), .B(n19576), .Z(n19564) );
  XNOR U19666 ( .A(n17620), .B(n19567), .Z(n19570) );
  XNOR U19667 ( .A(n17614), .B(n19577), .Z(n17671) );
  XNOR U19668 ( .A(n19578), .B(n19579), .Z(n19577) );
  NAND U19669 ( .A(n19580), .B(n18667), .Z(n19579) );
  XOR U19670 ( .A(n19581), .B(n19578), .Z(n17614) );
  NANDN U19671 ( .A(n19582), .B(n19583), .Z(n19578) );
  ANDN U19672 ( .B(n19584), .A(n19585), .Z(n19581) );
  XNOR U19673 ( .A(n18663), .B(n19586), .Z(n17602) );
  XNOR U19674 ( .A(n18661), .B(n19587), .Z(n19586) );
  NANDN U19675 ( .A(n19588), .B(n17625), .Z(n19587) );
  XNOR U19676 ( .A(n17677), .B(n17625), .Z(n17674) );
  XOR U19677 ( .A(n19590), .B(n18665), .Z(n18663) );
  OR U19678 ( .A(n19582), .B(n19591), .Z(n18665) );
  XNOR U19679 ( .A(n19592), .B(n18667), .Z(n19582) );
  XOR U19680 ( .A(n19567), .B(n17625), .Z(n18667) );
  XOR U19681 ( .A(n19593), .B(n19594), .Z(n17625) );
  NANDN U19682 ( .A(n19595), .B(n19596), .Z(n19594) );
  XOR U19683 ( .A(n19597), .B(n19598), .Z(n19567) );
  NANDN U19684 ( .A(n19595), .B(n19599), .Z(n19598) );
  ANDN U19685 ( .B(n19592), .A(n19600), .Z(n19590) );
  IV U19686 ( .A(n19585), .Z(n19592) );
  XOR U19687 ( .A(n17677), .B(n17620), .Z(n19585) );
  XNOR U19688 ( .A(n19601), .B(n19597), .Z(n17620) );
  NANDN U19689 ( .A(n19602), .B(n19603), .Z(n19597) );
  XOR U19690 ( .A(n19599), .B(n19604), .Z(n19603) );
  ANDN U19691 ( .B(n19604), .A(n19605), .Z(n19601) );
  XOR U19692 ( .A(n19606), .B(n19593), .Z(n17677) );
  NANDN U19693 ( .A(n19602), .B(n19607), .Z(n19593) );
  XOR U19694 ( .A(n19608), .B(n19596), .Z(n19607) );
  XNOR U19695 ( .A(n19609), .B(n19610), .Z(n19595) );
  XOR U19696 ( .A(n19611), .B(n19612), .Z(n19610) );
  XNOR U19697 ( .A(n19613), .B(n19614), .Z(n19609) );
  XNOR U19698 ( .A(n19615), .B(n19616), .Z(n19614) );
  ANDN U19699 ( .B(n19608), .A(n19612), .Z(n19615) );
  ANDN U19700 ( .B(n19608), .A(n19605), .Z(n19606) );
  XNOR U19701 ( .A(n19611), .B(n19617), .Z(n19605) );
  XOR U19702 ( .A(n19618), .B(n19616), .Z(n19617) );
  NAND U19703 ( .A(n19619), .B(n19620), .Z(n19616) );
  XNOR U19704 ( .A(n19613), .B(n19596), .Z(n19620) );
  IV U19705 ( .A(n19608), .Z(n19613) );
  XNOR U19706 ( .A(n19599), .B(n19612), .Z(n19619) );
  IV U19707 ( .A(n19604), .Z(n19612) );
  XOR U19708 ( .A(n19621), .B(n19622), .Z(n19604) );
  XNOR U19709 ( .A(n19623), .B(n19624), .Z(n19622) );
  XNOR U19710 ( .A(n19625), .B(n19626), .Z(n19621) );
  ANDN U19711 ( .B(n18662), .A(n17676), .Z(n19625) );
  AND U19712 ( .A(n19596), .B(n19599), .Z(n19618) );
  XNOR U19713 ( .A(n19596), .B(n19599), .Z(n19611) );
  XNOR U19714 ( .A(n19627), .B(n19628), .Z(n19599) );
  XNOR U19715 ( .A(n19629), .B(n19624), .Z(n19628) );
  XOR U19716 ( .A(n19630), .B(n19631), .Z(n19627) );
  XNOR U19717 ( .A(n19632), .B(n19626), .Z(n19631) );
  OR U19718 ( .A(n17675), .B(n19589), .Z(n19626) );
  XNOR U19719 ( .A(n18662), .B(n19633), .Z(n19589) );
  XNOR U19720 ( .A(n17676), .B(n17626), .Z(n17675) );
  ANDN U19721 ( .B(n19634), .A(n19588), .Z(n19632) );
  XNOR U19722 ( .A(n19635), .B(n19636), .Z(n19596) );
  XNOR U19723 ( .A(n19624), .B(n19637), .Z(n19636) );
  XOR U19724 ( .A(n19575), .B(n19630), .Z(n19637) );
  XNOR U19725 ( .A(n18662), .B(n17676), .Z(n19624) );
  XOR U19726 ( .A(n17619), .B(n19638), .Z(n19635) );
  XNOR U19727 ( .A(n19639), .B(n19640), .Z(n19638) );
  ANDN U19728 ( .B(n19641), .A(n19572), .Z(n19639) );
  XNOR U19729 ( .A(n19642), .B(n19643), .Z(n19608) );
  XNOR U19730 ( .A(n19629), .B(n19644), .Z(n19643) );
  XNOR U19731 ( .A(n19566), .B(n19623), .Z(n19644) );
  XOR U19732 ( .A(n19630), .B(n19645), .Z(n19623) );
  XNOR U19733 ( .A(n19646), .B(n19647), .Z(n19645) );
  NAND U19734 ( .A(n18668), .B(n19580), .Z(n19647) );
  XNOR U19735 ( .A(n19648), .B(n19646), .Z(n19630) );
  NANDN U19736 ( .A(n19591), .B(n19583), .Z(n19646) );
  XOR U19737 ( .A(n19584), .B(n19580), .Z(n19583) );
  XNOR U19738 ( .A(n19641), .B(n17626), .Z(n19580) );
  XOR U19739 ( .A(n19600), .B(n18668), .Z(n19591) );
  XNOR U19740 ( .A(n19572), .B(n19633), .Z(n18668) );
  ANDN U19741 ( .B(n19584), .A(n19600), .Z(n19648) );
  XOR U19742 ( .A(n17619), .B(n18662), .Z(n19600) );
  XNOR U19743 ( .A(n19649), .B(n19650), .Z(n18662) );
  XNOR U19744 ( .A(n19651), .B(n19652), .Z(n19650) );
  XOR U19745 ( .A(n19633), .B(n19634), .Z(n19629) );
  IV U19746 ( .A(n17626), .Z(n19634) );
  XOR U19747 ( .A(n19654), .B(n19655), .Z(n17626) );
  XOR U19748 ( .A(n19656), .B(n19652), .Z(n19655) );
  IV U19749 ( .A(n19588), .Z(n19633) );
  XOR U19750 ( .A(n19652), .B(n19657), .Z(n19588) );
  XNOR U19751 ( .A(n19658), .B(n19659), .Z(n19642) );
  XNOR U19752 ( .A(n19660), .B(n19640), .Z(n19659) );
  OR U19753 ( .A(n19576), .B(n19571), .Z(n19640) );
  XNOR U19754 ( .A(n17619), .B(n19572), .Z(n19571) );
  IV U19755 ( .A(n19658), .Z(n19572) );
  XOR U19756 ( .A(n19575), .B(n19641), .Z(n19576) );
  IV U19757 ( .A(n19566), .Z(n19641) );
  XOR U19758 ( .A(n19653), .B(n19661), .Z(n19566) );
  XNOR U19759 ( .A(n19662), .B(n19649), .Z(n19661) );
  XOR U19760 ( .A(n19663), .B(n19664), .Z(n19649) );
  XOR U19761 ( .A(n19665), .B(n16345), .Z(n19664) );
  XOR U19762 ( .A(n15620), .B(n19666), .Z(n19663) );
  XNOR U19763 ( .A(key[538]), .B(n17399), .Z(n19666) );
  XOR U19764 ( .A(n19667), .B(n19668), .Z(n17399) );
  XOR U19765 ( .A(n19669), .B(n19670), .Z(n19668) );
  XNOR U19766 ( .A(n15584), .B(n16356), .Z(n15620) );
  IV U19767 ( .A(n17676), .Z(n19653) );
  XOR U19768 ( .A(n19654), .B(n19673), .Z(n17676) );
  XOR U19769 ( .A(n19652), .B(n19674), .Z(n19673) );
  NOR U19770 ( .A(n19575), .B(n17619), .Z(n19660) );
  XOR U19771 ( .A(n19654), .B(n19675), .Z(n19575) );
  XOR U19772 ( .A(n19652), .B(n19676), .Z(n19675) );
  XOR U19773 ( .A(n19677), .B(n19678), .Z(n19652) );
  XNOR U19774 ( .A(n17619), .B(n17389), .Z(n19678) );
  XOR U19775 ( .A(n15598), .B(n17376), .Z(n17389) );
  XOR U19776 ( .A(n15627), .B(n16374), .Z(n17376) );
  XNOR U19777 ( .A(n19679), .B(n19680), .Z(n16374) );
  XNOR U19778 ( .A(n19681), .B(n19682), .Z(n19680) );
  XOR U19779 ( .A(n19672), .B(n19671), .Z(n19679) );
  XOR U19780 ( .A(n15593), .B(n16385), .Z(n15598) );
  XOR U19781 ( .A(n19683), .B(n19684), .Z(n15593) );
  XNOR U19782 ( .A(n15592), .B(n19685), .Z(n19677) );
  XNOR U19783 ( .A(key[542]), .B(n16394), .Z(n19685) );
  XOR U19784 ( .A(n19686), .B(n19687), .Z(n16394) );
  XNOR U19785 ( .A(n15606), .B(n16372), .Z(n15592) );
  IV U19786 ( .A(n19657), .Z(n19654) );
  XOR U19787 ( .A(n19688), .B(n19689), .Z(n19657) );
  XNOR U19788 ( .A(n16385), .B(n17380), .Z(n19689) );
  XNOR U19789 ( .A(n19690), .B(n19691), .Z(n15599) );
  XNOR U19790 ( .A(n19692), .B(n19693), .Z(n19691) );
  XNOR U19791 ( .A(n19694), .B(n19695), .Z(n19690) );
  XOR U19792 ( .A(n19696), .B(n19697), .Z(n19695) );
  ANDN U19793 ( .B(n19698), .A(n19699), .Z(n19697) );
  XOR U19794 ( .A(n19700), .B(n19701), .Z(n16385) );
  XOR U19795 ( .A(n16392), .B(n19702), .Z(n19688) );
  XNOR U19796 ( .A(key[541]), .B(n17381), .Z(n19702) );
  XOR U19797 ( .A(n19670), .B(n19681), .Z(n17381) );
  XNOR U19798 ( .A(n19703), .B(n19704), .Z(n19670) );
  XNOR U19799 ( .A(n19705), .B(n19706), .Z(n19704) );
  ANDN U19800 ( .B(n19707), .A(n19708), .Z(n19705) );
  XNOR U19801 ( .A(n19709), .B(n19710), .Z(n16392) );
  XNOR U19802 ( .A(n19711), .B(n19712), .Z(n19710) );
  XNOR U19803 ( .A(n19713), .B(n19714), .Z(n19709) );
  XOR U19804 ( .A(n19715), .B(n19716), .Z(n19714) );
  ANDN U19805 ( .B(n19717), .A(n19718), .Z(n19716) );
  XOR U19806 ( .A(n19719), .B(n19720), .Z(n19658) );
  XNOR U19807 ( .A(n19676), .B(n19674), .Z(n19720) );
  XNOR U19808 ( .A(n19721), .B(n19722), .Z(n19674) );
  XNOR U19809 ( .A(n16381), .B(n17377), .Z(n19722) );
  XOR U19810 ( .A(n16388), .B(n16372), .Z(n17377) );
  XNOR U19811 ( .A(n19723), .B(n19724), .Z(n16372) );
  XNOR U19812 ( .A(n19700), .B(n19725), .Z(n19724) );
  XOR U19813 ( .A(n19726), .B(n19727), .Z(n16388) );
  XNOR U19814 ( .A(n19683), .B(n19693), .Z(n19727) );
  XNOR U19815 ( .A(n19728), .B(n19729), .Z(n19693) );
  XNOR U19816 ( .A(n19730), .B(n19731), .Z(n19729) );
  NANDN U19817 ( .A(n19732), .B(n19733), .Z(n19731) );
  XOR U19818 ( .A(n15627), .B(n15606), .Z(n16381) );
  XNOR U19819 ( .A(key[543]), .B(n16373), .Z(n19721) );
  XOR U19820 ( .A(n19734), .B(n19735), .Z(n16373) );
  XNOR U19821 ( .A(n19687), .B(n19712), .Z(n19735) );
  XNOR U19822 ( .A(n19736), .B(n19737), .Z(n19712) );
  XNOR U19823 ( .A(n19738), .B(n19739), .Z(n19737) );
  NANDN U19824 ( .A(n19740), .B(n19741), .Z(n19739) );
  XNOR U19825 ( .A(n19742), .B(n19743), .Z(n19676) );
  XOR U19826 ( .A(n17367), .B(n17365), .Z(n19743) );
  XOR U19827 ( .A(n15611), .B(n16368), .Z(n17365) );
  XNOR U19828 ( .A(n19694), .B(n15584), .Z(n15611) );
  XOR U19829 ( .A(n15627), .B(n16393), .Z(n17367) );
  XNOR U19830 ( .A(n19746), .B(n19747), .Z(n16393) );
  XNOR U19831 ( .A(n19748), .B(n19682), .Z(n19747) );
  XNOR U19832 ( .A(n19749), .B(n19750), .Z(n19682) );
  XNOR U19833 ( .A(n19751), .B(n19752), .Z(n19750) );
  NANDN U19834 ( .A(n19753), .B(n19754), .Z(n19752) );
  XOR U19835 ( .A(n19755), .B(n19756), .Z(n19746) );
  XOR U19836 ( .A(n19706), .B(n19757), .Z(n19756) );
  ANDN U19837 ( .B(n19758), .A(n19759), .Z(n19757) );
  NOR U19838 ( .A(n19760), .B(n19761), .Z(n19706) );
  XNOR U19839 ( .A(n15610), .B(n19762), .Z(n19742) );
  XNOR U19840 ( .A(key[540]), .B(n16365), .Z(n19762) );
  XNOR U19841 ( .A(n19713), .B(n19665), .Z(n16365) );
  IV U19842 ( .A(n16348), .Z(n19665) );
  XOR U19843 ( .A(n19763), .B(n19764), .Z(n16348) );
  XNOR U19844 ( .A(n15606), .B(n16391), .Z(n15610) );
  XNOR U19845 ( .A(n19765), .B(n19766), .Z(n16391) );
  XOR U19846 ( .A(n19767), .B(n19725), .Z(n19766) );
  XNOR U19847 ( .A(n19768), .B(n19769), .Z(n19725) );
  XNOR U19848 ( .A(n19770), .B(n19771), .Z(n19769) );
  NANDN U19849 ( .A(n19772), .B(n19773), .Z(n19771) );
  XNOR U19850 ( .A(n19774), .B(n19775), .Z(n19765) );
  XNOR U19851 ( .A(n19776), .B(n19777), .Z(n19775) );
  ANDN U19852 ( .B(n19778), .A(n19779), .Z(n19777) );
  XNOR U19853 ( .A(n17619), .B(n19651), .Z(n19719) );
  XOR U19854 ( .A(n19780), .B(n19781), .Z(n19651) );
  XNOR U19855 ( .A(n17394), .B(n19782), .Z(n19781) );
  XOR U19856 ( .A(n15583), .B(n19662), .Z(n19782) );
  IV U19857 ( .A(n19656), .Z(n19662) );
  XNOR U19858 ( .A(n19783), .B(n19784), .Z(n19656) );
  XNOR U19859 ( .A(n16356), .B(n17397), .Z(n19784) );
  XOR U19860 ( .A(n17387), .B(n19785), .Z(n19783) );
  XOR U19861 ( .A(key[537]), .B(n15628), .Z(n19785) );
  XOR U19862 ( .A(n15621), .B(n16350), .Z(n15628) );
  IV U19863 ( .A(n16382), .Z(n15621) );
  XNOR U19864 ( .A(n19744), .B(n19787), .Z(n19786) );
  XOR U19865 ( .A(n19745), .B(n19788), .Z(n19683) );
  IV U19866 ( .A(n16380), .Z(n17387) );
  XNOR U19867 ( .A(n19687), .B(n19789), .Z(n16380) );
  XNOR U19868 ( .A(n19764), .B(n19790), .Z(n19789) );
  XOR U19869 ( .A(n19763), .B(n19791), .Z(n19687) );
  XOR U19870 ( .A(n15616), .B(n16345), .Z(n15583) );
  XNOR U19871 ( .A(n19723), .B(n19792), .Z(n16345) );
  XNOR U19872 ( .A(n19793), .B(n19701), .Z(n19792) );
  XOR U19873 ( .A(n19794), .B(n19795), .Z(n19701) );
  XOR U19874 ( .A(n19796), .B(n19776), .Z(n19795) );
  OR U19875 ( .A(n19797), .B(n19798), .Z(n19776) );
  NOR U19876 ( .A(n19799), .B(n19800), .Z(n19796) );
  IV U19877 ( .A(n16355), .Z(n15616) );
  XOR U19878 ( .A(n19726), .B(n19803), .Z(n16355) );
  XNOR U19879 ( .A(n19788), .B(n19684), .Z(n19803) );
  XNOR U19880 ( .A(n19804), .B(n19805), .Z(n19684) );
  XNOR U19881 ( .A(n19806), .B(n19696), .Z(n19805) );
  ANDN U19882 ( .B(n19807), .A(n19808), .Z(n19696) );
  NOR U19883 ( .A(n19809), .B(n19810), .Z(n19806) );
  XNOR U19884 ( .A(n19692), .B(n19811), .Z(n19788) );
  XNOR U19885 ( .A(n19812), .B(n19813), .Z(n19811) );
  NANDN U19886 ( .A(n19814), .B(n19815), .Z(n19813) );
  XOR U19887 ( .A(n19744), .B(n19787), .Z(n19726) );
  XNOR U19888 ( .A(n19812), .B(n19817), .Z(n19816) );
  NANDN U19889 ( .A(n19818), .B(n19733), .Z(n19817) );
  OR U19890 ( .A(n19819), .B(n19820), .Z(n19812) );
  XNOR U19891 ( .A(n19692), .B(n19821), .Z(n19804) );
  XNOR U19892 ( .A(n19822), .B(n19823), .Z(n19821) );
  NAND U19893 ( .A(n19824), .B(n19825), .Z(n19823) );
  XOR U19894 ( .A(n19826), .B(n19822), .Z(n19692) );
  NANDN U19895 ( .A(n19827), .B(n19828), .Z(n19822) );
  ANDN U19896 ( .B(n19829), .A(n19830), .Z(n19826) );
  XOR U19897 ( .A(n19831), .B(n19832), .Z(n19744) );
  XOR U19898 ( .A(n19833), .B(n19834), .Z(n19832) );
  NANDN U19899 ( .A(n19835), .B(n19698), .Z(n19834) );
  XNOR U19900 ( .A(n15627), .B(n16366), .Z(n17394) );
  XNOR U19901 ( .A(n19755), .B(n17397), .Z(n16366) );
  XOR U19902 ( .A(n19836), .B(n19672), .Z(n17397) );
  XNOR U19903 ( .A(n19836), .B(n19755), .Z(n15627) );
  XOR U19904 ( .A(n19749), .B(n19837), .Z(n19755) );
  XNOR U19905 ( .A(n19838), .B(n19839), .Z(n19837) );
  ANDN U19906 ( .B(n19707), .A(n19840), .Z(n19838) );
  XOR U19907 ( .A(n19841), .B(n19842), .Z(n19749) );
  XNOR U19908 ( .A(n19843), .B(n19844), .Z(n19842) );
  NAND U19909 ( .A(n19845), .B(n19846), .Z(n19844) );
  XNOR U19910 ( .A(n15614), .B(n19847), .Z(n19780) );
  XOR U19911 ( .A(key[539]), .B(n17402), .Z(n19847) );
  XNOR U19912 ( .A(n19734), .B(n19848), .Z(n17402) );
  XOR U19913 ( .A(n19791), .B(n19686), .Z(n19848) );
  XNOR U19914 ( .A(n19849), .B(n19850), .Z(n19686) );
  XNOR U19915 ( .A(n19851), .B(n19715), .Z(n19850) );
  NOR U19916 ( .A(n19852), .B(n19853), .Z(n19715) );
  ANDN U19917 ( .B(n19854), .A(n19855), .Z(n19851) );
  XNOR U19918 ( .A(n19711), .B(n19856), .Z(n19791) );
  XNOR U19919 ( .A(n19857), .B(n19858), .Z(n19856) );
  NANDN U19920 ( .A(n19859), .B(n19860), .Z(n19858) );
  XOR U19921 ( .A(n19764), .B(n19790), .Z(n19734) );
  XNOR U19922 ( .A(n19849), .B(n19861), .Z(n19790) );
  XNOR U19923 ( .A(n19857), .B(n19862), .Z(n19861) );
  NANDN U19924 ( .A(n19863), .B(n19741), .Z(n19862) );
  OR U19925 ( .A(n19864), .B(n19865), .Z(n19857) );
  XOR U19926 ( .A(n19711), .B(n19866), .Z(n19849) );
  XNOR U19927 ( .A(n19867), .B(n19868), .Z(n19866) );
  NAND U19928 ( .A(n19869), .B(n19870), .Z(n19868) );
  XOR U19929 ( .A(n19871), .B(n19867), .Z(n19711) );
  NANDN U19930 ( .A(n19872), .B(n19873), .Z(n19867) );
  ANDN U19931 ( .B(n19874), .A(n19875), .Z(n19871) );
  XOR U19932 ( .A(n19877), .B(n19878), .Z(n19876) );
  NANDN U19933 ( .A(n19879), .B(n19717), .Z(n19878) );
  XOR U19934 ( .A(n15606), .B(n16368), .Z(n15614) );
  XNOR U19935 ( .A(n16356), .B(n19767), .Z(n16368) );
  XOR U19936 ( .A(n19802), .B(n19881), .Z(n16356) );
  XNOR U19937 ( .A(n19882), .B(n19883), .Z(n17619) );
  XNOR U19938 ( .A(n17388), .B(n15606), .Z(n19883) );
  XOR U19939 ( .A(n19881), .B(n19767), .Z(n15606) );
  XOR U19940 ( .A(n19768), .B(n19884), .Z(n19767) );
  XNOR U19941 ( .A(n19885), .B(n19886), .Z(n19884) );
  ANDN U19942 ( .B(n19887), .A(n19800), .Z(n19885) );
  XOR U19943 ( .A(n19888), .B(n19889), .Z(n19768) );
  XNOR U19944 ( .A(n19890), .B(n19891), .Z(n19889) );
  NANDN U19945 ( .A(n19892), .B(n19893), .Z(n19891) );
  XOR U19946 ( .A(n19681), .B(n19894), .Z(n17388) );
  XNOR U19947 ( .A(n19672), .B(n19671), .Z(n19894) );
  XNOR U19948 ( .A(n19703), .B(n19895), .Z(n19671) );
  XNOR U19949 ( .A(n19896), .B(n19897), .Z(n19895) );
  NANDN U19950 ( .A(n19898), .B(n19754), .Z(n19897) );
  XOR U19951 ( .A(n19748), .B(n19899), .Z(n19703) );
  XNOR U19952 ( .A(n19900), .B(n19901), .Z(n19899) );
  NAND U19953 ( .A(n19902), .B(n19845), .Z(n19901) );
  XOR U19954 ( .A(n19839), .B(n19904), .Z(n19903) );
  NANDN U19955 ( .A(n19905), .B(n19758), .Z(n19904) );
  XNOR U19956 ( .A(n19707), .B(n19758), .Z(n19760) );
  XOR U19957 ( .A(n19836), .B(n19669), .Z(n19681) );
  XNOR U19958 ( .A(n19748), .B(n19907), .Z(n19669) );
  XNOR U19959 ( .A(n19896), .B(n19908), .Z(n19907) );
  NANDN U19960 ( .A(n19909), .B(n19910), .Z(n19908) );
  OR U19961 ( .A(n19911), .B(n19912), .Z(n19896) );
  XOR U19962 ( .A(n19913), .B(n19900), .Z(n19748) );
  NANDN U19963 ( .A(n19914), .B(n19915), .Z(n19900) );
  ANDN U19964 ( .B(n19916), .A(n19917), .Z(n19913) );
  XNOR U19965 ( .A(n19841), .B(n19918), .Z(n19836) );
  XOR U19966 ( .A(n19919), .B(n19751), .Z(n19918) );
  OR U19967 ( .A(n19920), .B(n19911), .Z(n19751) );
  XNOR U19968 ( .A(n19754), .B(n19910), .Z(n19911) );
  ANDN U19969 ( .B(n19910), .A(n19921), .Z(n19919) );
  XNOR U19970 ( .A(n19922), .B(n19843), .Z(n19841) );
  OR U19971 ( .A(n19914), .B(n19923), .Z(n19843) );
  XNOR U19972 ( .A(n19924), .B(n19845), .Z(n19914) );
  XOR U19973 ( .A(n19910), .B(n19758), .Z(n19845) );
  XOR U19974 ( .A(n19925), .B(n19926), .Z(n19758) );
  NANDN U19975 ( .A(n19927), .B(n19928), .Z(n19926) );
  XOR U19976 ( .A(n19929), .B(n19930), .Z(n19910) );
  NANDN U19977 ( .A(n19927), .B(n19931), .Z(n19930) );
  ANDN U19978 ( .B(n19924), .A(n19932), .Z(n19922) );
  IV U19979 ( .A(n19917), .Z(n19924) );
  XNOR U19980 ( .A(n19707), .B(n19754), .Z(n19917) );
  XNOR U19981 ( .A(n19933), .B(n19929), .Z(n19754) );
  NANDN U19982 ( .A(n19934), .B(n19935), .Z(n19929) );
  XOR U19983 ( .A(n19931), .B(n19936), .Z(n19935) );
  ANDN U19984 ( .B(n19936), .A(n19937), .Z(n19933) );
  XNOR U19985 ( .A(n19938), .B(n19925), .Z(n19707) );
  NANDN U19986 ( .A(n19934), .B(n19939), .Z(n19925) );
  XOR U19987 ( .A(n19940), .B(n19928), .Z(n19939) );
  XNOR U19988 ( .A(n19941), .B(n19942), .Z(n19927) );
  XOR U19989 ( .A(n19943), .B(n19944), .Z(n19942) );
  XNOR U19990 ( .A(n19945), .B(n19946), .Z(n19941) );
  XNOR U19991 ( .A(n19947), .B(n19948), .Z(n19946) );
  ANDN U19992 ( .B(n19940), .A(n19944), .Z(n19947) );
  ANDN U19993 ( .B(n19940), .A(n19937), .Z(n19938) );
  XNOR U19994 ( .A(n19943), .B(n19949), .Z(n19937) );
  XOR U19995 ( .A(n19950), .B(n19948), .Z(n19949) );
  NAND U19996 ( .A(n19951), .B(n19952), .Z(n19948) );
  XNOR U19997 ( .A(n19945), .B(n19928), .Z(n19952) );
  IV U19998 ( .A(n19940), .Z(n19945) );
  XNOR U19999 ( .A(n19931), .B(n19944), .Z(n19951) );
  IV U20000 ( .A(n19936), .Z(n19944) );
  XOR U20001 ( .A(n19953), .B(n19954), .Z(n19936) );
  XNOR U20002 ( .A(n19955), .B(n19956), .Z(n19954) );
  XNOR U20003 ( .A(n19957), .B(n19958), .Z(n19953) );
  NOR U20004 ( .A(n19708), .B(n19840), .Z(n19957) );
  AND U20005 ( .A(n19928), .B(n19931), .Z(n19950) );
  XNOR U20006 ( .A(n19928), .B(n19931), .Z(n19943) );
  XNOR U20007 ( .A(n19959), .B(n19960), .Z(n19931) );
  XNOR U20008 ( .A(n19961), .B(n19956), .Z(n19960) );
  XOR U20009 ( .A(n19962), .B(n19963), .Z(n19959) );
  XNOR U20010 ( .A(n19964), .B(n19958), .Z(n19963) );
  OR U20011 ( .A(n19761), .B(n19906), .Z(n19958) );
  XNOR U20012 ( .A(n19840), .B(n19905), .Z(n19906) );
  XNOR U20013 ( .A(n19708), .B(n19759), .Z(n19761) );
  ANDN U20014 ( .B(n19965), .A(n19905), .Z(n19964) );
  XNOR U20015 ( .A(n19966), .B(n19967), .Z(n19928) );
  XNOR U20016 ( .A(n19956), .B(n19968), .Z(n19967) );
  XOR U20017 ( .A(n19898), .B(n19962), .Z(n19968) );
  XNOR U20018 ( .A(n19840), .B(n19969), .Z(n19956) );
  XOR U20019 ( .A(n19753), .B(n19970), .Z(n19966) );
  XNOR U20020 ( .A(n19971), .B(n19972), .Z(n19970) );
  ANDN U20021 ( .B(n19973), .A(n19921), .Z(n19971) );
  XNOR U20022 ( .A(n19974), .B(n19975), .Z(n19940) );
  XNOR U20023 ( .A(n19961), .B(n19976), .Z(n19975) );
  XNOR U20024 ( .A(n19909), .B(n19955), .Z(n19976) );
  XOR U20025 ( .A(n19962), .B(n19977), .Z(n19955) );
  XNOR U20026 ( .A(n19978), .B(n19979), .Z(n19977) );
  NAND U20027 ( .A(n19846), .B(n19902), .Z(n19979) );
  XNOR U20028 ( .A(n19980), .B(n19978), .Z(n19962) );
  NANDN U20029 ( .A(n19923), .B(n19915), .Z(n19978) );
  XOR U20030 ( .A(n19916), .B(n19902), .Z(n19915) );
  XNOR U20031 ( .A(n19973), .B(n19759), .Z(n19902) );
  XOR U20032 ( .A(n19932), .B(n19846), .Z(n19923) );
  XNOR U20033 ( .A(n19921), .B(n19981), .Z(n19846) );
  ANDN U20034 ( .B(n19916), .A(n19932), .Z(n19980) );
  XNOR U20035 ( .A(n19753), .B(n19840), .Z(n19932) );
  XOR U20036 ( .A(n19982), .B(n19983), .Z(n19840) );
  XNOR U20037 ( .A(n19984), .B(n19985), .Z(n19983) );
  XOR U20038 ( .A(n19981), .B(n19965), .Z(n19961) );
  IV U20039 ( .A(n19759), .Z(n19965) );
  XOR U20040 ( .A(n19986), .B(n19987), .Z(n19759) );
  XNOR U20041 ( .A(n19988), .B(n19985), .Z(n19987) );
  IV U20042 ( .A(n19905), .Z(n19981) );
  XOR U20043 ( .A(n19985), .B(n19989), .Z(n19905) );
  XNOR U20044 ( .A(n19990), .B(n19991), .Z(n19974) );
  XNOR U20045 ( .A(n19992), .B(n19972), .Z(n19991) );
  OR U20046 ( .A(n19912), .B(n19920), .Z(n19972) );
  XNOR U20047 ( .A(n19753), .B(n19921), .Z(n19920) );
  IV U20048 ( .A(n19990), .Z(n19921) );
  XOR U20049 ( .A(n19898), .B(n19973), .Z(n19912) );
  IV U20050 ( .A(n19909), .Z(n19973) );
  XOR U20051 ( .A(n19969), .B(n19993), .Z(n19909) );
  XNOR U20052 ( .A(n19988), .B(n19982), .Z(n19993) );
  XOR U20053 ( .A(n19994), .B(n19995), .Z(n19982) );
  XNOR U20054 ( .A(n19996), .B(n19424), .Z(n19995) );
  IV U20055 ( .A(n18470), .Z(n19424) );
  XNOR U20056 ( .A(n19997), .B(n19409), .Z(n18470) );
  XNOR U20057 ( .A(key[410]), .B(n19999), .Z(n19998) );
  IV U20058 ( .A(n19708), .Z(n19969) );
  XOR U20059 ( .A(n19986), .B(n20000), .Z(n19708) );
  XOR U20060 ( .A(n19985), .B(n20001), .Z(n20000) );
  NOR U20061 ( .A(n19898), .B(n19753), .Z(n19992) );
  XOR U20062 ( .A(n19986), .B(n20002), .Z(n19898) );
  XOR U20063 ( .A(n19985), .B(n20003), .Z(n20002) );
  XOR U20064 ( .A(n20004), .B(n20005), .Z(n19985) );
  XOR U20065 ( .A(n18478), .B(n19413), .Z(n20005) );
  XOR U20066 ( .A(n19405), .B(n20006), .Z(n19413) );
  XNOR U20067 ( .A(n19399), .B(n18491), .Z(n18478) );
  XNOR U20068 ( .A(n20007), .B(n20008), .Z(n18491) );
  XOR U20069 ( .A(n20009), .B(n19414), .Z(n19399) );
  XOR U20070 ( .A(n19753), .B(n20010), .Z(n20004) );
  XNOR U20071 ( .A(key[414]), .B(n20011), .Z(n20010) );
  IV U20072 ( .A(n19989), .Z(n19986) );
  XOR U20073 ( .A(n20012), .B(n20013), .Z(n19989) );
  XNOR U20074 ( .A(n20014), .B(n18485), .Z(n20013) );
  XOR U20075 ( .A(n20015), .B(n20016), .Z(n18485) );
  XOR U20076 ( .A(key[413]), .B(n20009), .Z(n20017) );
  XOR U20077 ( .A(n20018), .B(n20019), .Z(n19990) );
  XNOR U20078 ( .A(n20003), .B(n20001), .Z(n20019) );
  XNOR U20079 ( .A(n20020), .B(n20021), .Z(n20001) );
  XOR U20080 ( .A(n20022), .B(n18492), .Z(n20021) );
  XNOR U20081 ( .A(n20023), .B(n20006), .Z(n18492) );
  XNOR U20082 ( .A(key[415]), .B(n18518), .Z(n20020) );
  XNOR U20083 ( .A(n20024), .B(n20025), .Z(n20003) );
  XNOR U20084 ( .A(n18497), .B(n19390), .Z(n20025) );
  XOR U20085 ( .A(n20026), .B(n20016), .Z(n19390) );
  XOR U20086 ( .A(n19391), .B(n20027), .Z(n18497) );
  XNOR U20087 ( .A(n18496), .B(n20028), .Z(n20024) );
  XOR U20088 ( .A(key[412]), .B(n20029), .Z(n20028) );
  XNOR U20089 ( .A(n20007), .B(n18484), .Z(n18496) );
  XNOR U20090 ( .A(n19753), .B(n19984), .Z(n20018) );
  XOR U20091 ( .A(n20030), .B(n20031), .Z(n19984) );
  XOR U20092 ( .A(n19421), .B(n20032), .Z(n20031) );
  XOR U20093 ( .A(n19988), .B(n19410), .Z(n20032) );
  IV U20094 ( .A(n18505), .Z(n19410) );
  XOR U20095 ( .A(n20033), .B(n19996), .Z(n18505) );
  XOR U20096 ( .A(n20034), .B(n20035), .Z(n19988) );
  XNOR U20097 ( .A(n18471), .B(n18509), .Z(n20035) );
  XOR U20098 ( .A(n19425), .B(n20036), .Z(n18509) );
  XOR U20099 ( .A(n19997), .B(n20037), .Z(n20034) );
  XOR U20100 ( .A(key[409]), .B(n20038), .Z(n20037) );
  XNOR U20101 ( .A(n20026), .B(n20027), .Z(n19421) );
  XNOR U20102 ( .A(n18504), .B(n20039), .Z(n20030) );
  XOR U20103 ( .A(key[411]), .B(n20040), .Z(n20039) );
  XNOR U20104 ( .A(n20007), .B(n18500), .Z(n18504) );
  XNOR U20105 ( .A(n20041), .B(n20042), .Z(n19753) );
  XNOR U20106 ( .A(n20036), .B(n19430), .Z(n20042) );
  XNOR U20107 ( .A(n18508), .B(n20043), .Z(n20041) );
  XOR U20108 ( .A(key[408]), .B(n20026), .Z(n20043) );
  XOR U20109 ( .A(n16350), .B(n20044), .Z(n19882) );
  XOR U20110 ( .A(key[536]), .B(n15629), .Z(n20044) );
  XNOR U20111 ( .A(n16352), .B(n16384), .Z(n15629) );
  IV U20112 ( .A(n17366), .Z(n16384) );
  XNOR U20113 ( .A(n19763), .B(n19713), .Z(n17366) );
  XNOR U20114 ( .A(n19736), .B(n20045), .Z(n19713) );
  XNOR U20115 ( .A(n20046), .B(n19877), .Z(n20045) );
  XNOR U20116 ( .A(n19854), .B(n19717), .Z(n19852) );
  ANDN U20117 ( .B(n19854), .A(n20048), .Z(n20046) );
  XOR U20118 ( .A(n19880), .B(n20049), .Z(n19736) );
  XNOR U20119 ( .A(n20050), .B(n20051), .Z(n20049) );
  NAND U20120 ( .A(n19870), .B(n20052), .Z(n20051) );
  XNOR U20121 ( .A(n19880), .B(n20053), .Z(n19763) );
  XOR U20122 ( .A(n20054), .B(n19738), .Z(n20053) );
  OR U20123 ( .A(n20055), .B(n19864), .Z(n19738) );
  XNOR U20124 ( .A(n19741), .B(n19860), .Z(n19864) );
  ANDN U20125 ( .B(n19860), .A(n20056), .Z(n20054) );
  XNOR U20126 ( .A(n20057), .B(n20050), .Z(n19880) );
  OR U20127 ( .A(n19872), .B(n20058), .Z(n20050) );
  XNOR U20128 ( .A(n20059), .B(n19870), .Z(n19872) );
  XOR U20129 ( .A(n19860), .B(n19717), .Z(n19870) );
  XOR U20130 ( .A(n20060), .B(n20061), .Z(n19717) );
  NANDN U20131 ( .A(n20062), .B(n20063), .Z(n20061) );
  XOR U20132 ( .A(n20064), .B(n20065), .Z(n19860) );
  NANDN U20133 ( .A(n20062), .B(n20066), .Z(n20065) );
  ANDN U20134 ( .B(n20059), .A(n20067), .Z(n20057) );
  IV U20135 ( .A(n19875), .Z(n20059) );
  XNOR U20136 ( .A(n19854), .B(n19741), .Z(n19875) );
  XNOR U20137 ( .A(n20068), .B(n20064), .Z(n19741) );
  NANDN U20138 ( .A(n20069), .B(n20070), .Z(n20064) );
  XOR U20139 ( .A(n20066), .B(n20071), .Z(n20070) );
  ANDN U20140 ( .B(n20071), .A(n20072), .Z(n20068) );
  XNOR U20141 ( .A(n20073), .B(n20060), .Z(n19854) );
  NANDN U20142 ( .A(n20069), .B(n20074), .Z(n20060) );
  XOR U20143 ( .A(n20075), .B(n20063), .Z(n20074) );
  XNOR U20144 ( .A(n20076), .B(n20077), .Z(n20062) );
  XOR U20145 ( .A(n20078), .B(n20079), .Z(n20077) );
  XNOR U20146 ( .A(n20080), .B(n20081), .Z(n20076) );
  XNOR U20147 ( .A(n20082), .B(n20083), .Z(n20081) );
  ANDN U20148 ( .B(n20075), .A(n20079), .Z(n20082) );
  ANDN U20149 ( .B(n20075), .A(n20072), .Z(n20073) );
  XNOR U20150 ( .A(n20078), .B(n20084), .Z(n20072) );
  XOR U20151 ( .A(n20085), .B(n20083), .Z(n20084) );
  NAND U20152 ( .A(n20086), .B(n20087), .Z(n20083) );
  XNOR U20153 ( .A(n20080), .B(n20063), .Z(n20087) );
  IV U20154 ( .A(n20075), .Z(n20080) );
  XNOR U20155 ( .A(n20066), .B(n20079), .Z(n20086) );
  IV U20156 ( .A(n20071), .Z(n20079) );
  XOR U20157 ( .A(n20088), .B(n20089), .Z(n20071) );
  XNOR U20158 ( .A(n20090), .B(n20091), .Z(n20089) );
  XNOR U20159 ( .A(n20092), .B(n20093), .Z(n20088) );
  NOR U20160 ( .A(n19855), .B(n20048), .Z(n20092) );
  AND U20161 ( .A(n20063), .B(n20066), .Z(n20085) );
  XNOR U20162 ( .A(n20063), .B(n20066), .Z(n20078) );
  XNOR U20163 ( .A(n20094), .B(n20095), .Z(n20066) );
  XNOR U20164 ( .A(n20096), .B(n20091), .Z(n20095) );
  XOR U20165 ( .A(n20097), .B(n20098), .Z(n20094) );
  XNOR U20166 ( .A(n20099), .B(n20093), .Z(n20098) );
  OR U20167 ( .A(n19853), .B(n20047), .Z(n20093) );
  XNOR U20168 ( .A(n20048), .B(n19879), .Z(n20047) );
  XNOR U20169 ( .A(n19855), .B(n19718), .Z(n19853) );
  ANDN U20170 ( .B(n20100), .A(n19879), .Z(n20099) );
  XNOR U20171 ( .A(n20101), .B(n20102), .Z(n20063) );
  XNOR U20172 ( .A(n20091), .B(n20103), .Z(n20102) );
  XOR U20173 ( .A(n19863), .B(n20097), .Z(n20103) );
  XNOR U20174 ( .A(n20048), .B(n20104), .Z(n20091) );
  XOR U20175 ( .A(n19740), .B(n20105), .Z(n20101) );
  XNOR U20176 ( .A(n20106), .B(n20107), .Z(n20105) );
  ANDN U20177 ( .B(n20108), .A(n20056), .Z(n20106) );
  XNOR U20178 ( .A(n20109), .B(n20110), .Z(n20075) );
  XNOR U20179 ( .A(n20096), .B(n20111), .Z(n20110) );
  XNOR U20180 ( .A(n19859), .B(n20090), .Z(n20111) );
  XOR U20181 ( .A(n20097), .B(n20112), .Z(n20090) );
  XNOR U20182 ( .A(n20113), .B(n20114), .Z(n20112) );
  NAND U20183 ( .A(n20052), .B(n19869), .Z(n20114) );
  XNOR U20184 ( .A(n20115), .B(n20113), .Z(n20097) );
  NANDN U20185 ( .A(n20058), .B(n19873), .Z(n20113) );
  XOR U20186 ( .A(n19874), .B(n19869), .Z(n19873) );
  XNOR U20187 ( .A(n20108), .B(n19718), .Z(n19869) );
  XOR U20188 ( .A(n20067), .B(n20052), .Z(n20058) );
  XNOR U20189 ( .A(n20056), .B(n20116), .Z(n20052) );
  ANDN U20190 ( .B(n19874), .A(n20067), .Z(n20115) );
  XNOR U20191 ( .A(n19740), .B(n20048), .Z(n20067) );
  XOR U20192 ( .A(n20117), .B(n20118), .Z(n20048) );
  XNOR U20193 ( .A(n20119), .B(n20120), .Z(n20118) );
  XOR U20194 ( .A(n20116), .B(n20100), .Z(n20096) );
  IV U20195 ( .A(n19718), .Z(n20100) );
  XOR U20196 ( .A(n20121), .B(n20122), .Z(n19718) );
  XNOR U20197 ( .A(n20123), .B(n20120), .Z(n20122) );
  IV U20198 ( .A(n19879), .Z(n20116) );
  XOR U20199 ( .A(n20120), .B(n20124), .Z(n19879) );
  XNOR U20200 ( .A(n20125), .B(n20126), .Z(n20109) );
  XNOR U20201 ( .A(n20127), .B(n20107), .Z(n20126) );
  OR U20202 ( .A(n19865), .B(n20055), .Z(n20107) );
  XNOR U20203 ( .A(n19740), .B(n20056), .Z(n20055) );
  IV U20204 ( .A(n20125), .Z(n20056) );
  XOR U20205 ( .A(n19863), .B(n20108), .Z(n19865) );
  IV U20206 ( .A(n19859), .Z(n20108) );
  XOR U20207 ( .A(n20104), .B(n20128), .Z(n19859) );
  XNOR U20208 ( .A(n20123), .B(n20117), .Z(n20128) );
  XOR U20209 ( .A(n20129), .B(n20130), .Z(n20117) );
  XNOR U20210 ( .A(n19258), .B(n19294), .Z(n20130) );
  XNOR U20211 ( .A(key[418]), .B(n20131), .Z(n20129) );
  IV U20212 ( .A(n19855), .Z(n20104) );
  XOR U20213 ( .A(n20121), .B(n20132), .Z(n19855) );
  XOR U20214 ( .A(n20120), .B(n20133), .Z(n20132) );
  NOR U20215 ( .A(n19863), .B(n19740), .Z(n20127) );
  XOR U20216 ( .A(n20121), .B(n20134), .Z(n19863) );
  XOR U20217 ( .A(n20120), .B(n20135), .Z(n20134) );
  XOR U20218 ( .A(n20136), .B(n20137), .Z(n20120) );
  XOR U20219 ( .A(n18633), .B(n19267), .Z(n20137) );
  XNOR U20220 ( .A(n20138), .B(n20139), .Z(n19267) );
  XNOR U20221 ( .A(n20140), .B(n19281), .Z(n18633) );
  XOR U20222 ( .A(n19740), .B(n20141), .Z(n20136) );
  XNOR U20223 ( .A(key[422]), .B(n19275), .Z(n20141) );
  IV U20224 ( .A(n20124), .Z(n20121) );
  XOR U20225 ( .A(n20142), .B(n20143), .Z(n20124) );
  XNOR U20226 ( .A(n20144), .B(n19272), .Z(n20143) );
  XNOR U20227 ( .A(n20145), .B(n18613), .Z(n19272) );
  XNOR U20228 ( .A(key[421]), .B(n20146), .Z(n20142) );
  XOR U20229 ( .A(n20147), .B(n20148), .Z(n20125) );
  XNOR U20230 ( .A(n20135), .B(n20133), .Z(n20148) );
  XNOR U20231 ( .A(n20149), .B(n20150), .Z(n20133) );
  XOR U20232 ( .A(n20139), .B(n19280), .Z(n20150) );
  XNOR U20233 ( .A(n20151), .B(n18620), .Z(n19280) );
  XOR U20234 ( .A(n20152), .B(n20153), .Z(n20139) );
  XNOR U20235 ( .A(key[423]), .B(n20140), .Z(n20149) );
  XNOR U20236 ( .A(n20154), .B(n19283), .Z(n20135) );
  XOR U20237 ( .A(n20155), .B(n20156), .Z(n19283) );
  XOR U20238 ( .A(n20157), .B(n18608), .Z(n20156) );
  XNOR U20239 ( .A(n20158), .B(n20144), .Z(n20155) );
  XNOR U20240 ( .A(n18605), .B(n20159), .Z(n20154) );
  XOR U20241 ( .A(key[420]), .B(n20160), .Z(n20159) );
  XOR U20242 ( .A(n20140), .B(n19273), .Z(n18605) );
  XNOR U20243 ( .A(n19740), .B(n20119), .Z(n20147) );
  XOR U20244 ( .A(n20161), .B(n20162), .Z(n20119) );
  XOR U20245 ( .A(n19291), .B(n20163), .Z(n20162) );
  XOR U20246 ( .A(n20123), .B(n18641), .Z(n20163) );
  XOR U20247 ( .A(n18656), .B(n19286), .Z(n18641) );
  XOR U20248 ( .A(n20164), .B(n20165), .Z(n20123) );
  XOR U20249 ( .A(n20166), .B(n18627), .Z(n20165) );
  XNOR U20250 ( .A(key[417]), .B(n19297), .Z(n20164) );
  XOR U20251 ( .A(n20158), .B(n20160), .Z(n19291) );
  XOR U20252 ( .A(n19290), .B(n20167), .Z(n20161) );
  XNOR U20253 ( .A(key[419]), .B(n19260), .Z(n20167) );
  XNOR U20254 ( .A(n20168), .B(n20169), .Z(n19740) );
  XNOR U20255 ( .A(n18648), .B(n18655), .Z(n20169) );
  XNOR U20256 ( .A(n20152), .B(n19303), .Z(n18655) );
  XNOR U20257 ( .A(key[416]), .B(n20170), .Z(n20168) );
  IV U20258 ( .A(n16367), .Z(n16352) );
  XOR U20259 ( .A(n19694), .B(n19745), .Z(n16367) );
  XOR U20260 ( .A(n19831), .B(n20171), .Z(n19745) );
  XOR U20261 ( .A(n20172), .B(n19730), .Z(n20171) );
  OR U20262 ( .A(n20173), .B(n19819), .Z(n19730) );
  XNOR U20263 ( .A(n19733), .B(n19815), .Z(n19819) );
  ANDN U20264 ( .B(n19815), .A(n20174), .Z(n20172) );
  IV U20265 ( .A(n20175), .Z(n19831) );
  XNOR U20266 ( .A(n19728), .B(n20176), .Z(n19694) );
  XNOR U20267 ( .A(n20177), .B(n19833), .Z(n20176) );
  XNOR U20268 ( .A(n19810), .B(n19698), .Z(n19807) );
  ANDN U20269 ( .B(n20179), .A(n19810), .Z(n20177) );
  XOR U20270 ( .A(n20175), .B(n20180), .Z(n19728) );
  XNOR U20271 ( .A(n20181), .B(n20182), .Z(n20180) );
  NAND U20272 ( .A(n19825), .B(n20183), .Z(n20182) );
  XNOR U20273 ( .A(n20184), .B(n20181), .Z(n20175) );
  OR U20274 ( .A(n19827), .B(n20185), .Z(n20181) );
  XNOR U20275 ( .A(n20186), .B(n19825), .Z(n19827) );
  XOR U20276 ( .A(n19815), .B(n19698), .Z(n19825) );
  XOR U20277 ( .A(n20187), .B(n20188), .Z(n19698) );
  NANDN U20278 ( .A(n20189), .B(n20190), .Z(n20188) );
  XOR U20279 ( .A(n20191), .B(n20192), .Z(n19815) );
  NANDN U20280 ( .A(n20189), .B(n20193), .Z(n20192) );
  ANDN U20281 ( .B(n20186), .A(n20194), .Z(n20184) );
  IV U20282 ( .A(n19830), .Z(n20186) );
  XOR U20283 ( .A(n19810), .B(n19733), .Z(n19830) );
  XNOR U20284 ( .A(n20195), .B(n20191), .Z(n19733) );
  NANDN U20285 ( .A(n20196), .B(n20197), .Z(n20191) );
  XOR U20286 ( .A(n20193), .B(n20198), .Z(n20197) );
  ANDN U20287 ( .B(n20198), .A(n20199), .Z(n20195) );
  XOR U20288 ( .A(n20200), .B(n20187), .Z(n19810) );
  NANDN U20289 ( .A(n20196), .B(n20201), .Z(n20187) );
  XOR U20290 ( .A(n20202), .B(n20190), .Z(n20201) );
  XNOR U20291 ( .A(n20203), .B(n20204), .Z(n20189) );
  XOR U20292 ( .A(n20205), .B(n20206), .Z(n20204) );
  XNOR U20293 ( .A(n20207), .B(n20208), .Z(n20203) );
  XNOR U20294 ( .A(n20209), .B(n20210), .Z(n20208) );
  ANDN U20295 ( .B(n20202), .A(n20206), .Z(n20209) );
  ANDN U20296 ( .B(n20202), .A(n20199), .Z(n20200) );
  XNOR U20297 ( .A(n20205), .B(n20211), .Z(n20199) );
  XOR U20298 ( .A(n20212), .B(n20210), .Z(n20211) );
  NAND U20299 ( .A(n20213), .B(n20214), .Z(n20210) );
  XNOR U20300 ( .A(n20207), .B(n20190), .Z(n20214) );
  IV U20301 ( .A(n20202), .Z(n20207) );
  XNOR U20302 ( .A(n20193), .B(n20206), .Z(n20213) );
  IV U20303 ( .A(n20198), .Z(n20206) );
  XOR U20304 ( .A(n20215), .B(n20216), .Z(n20198) );
  XNOR U20305 ( .A(n20217), .B(n20218), .Z(n20216) );
  XNOR U20306 ( .A(n20219), .B(n20220), .Z(n20215) );
  ANDN U20307 ( .B(n20179), .A(n19809), .Z(n20219) );
  AND U20308 ( .A(n20190), .B(n20193), .Z(n20212) );
  XNOR U20309 ( .A(n20190), .B(n20193), .Z(n20205) );
  XNOR U20310 ( .A(n20221), .B(n20222), .Z(n20193) );
  XNOR U20311 ( .A(n20223), .B(n20218), .Z(n20222) );
  XOR U20312 ( .A(n20224), .B(n20225), .Z(n20221) );
  XNOR U20313 ( .A(n20226), .B(n20220), .Z(n20225) );
  OR U20314 ( .A(n19808), .B(n20178), .Z(n20220) );
  XNOR U20315 ( .A(n20179), .B(n20227), .Z(n20178) );
  XNOR U20316 ( .A(n19809), .B(n19699), .Z(n19808) );
  ANDN U20317 ( .B(n20228), .A(n19835), .Z(n20226) );
  XNOR U20318 ( .A(n20229), .B(n20230), .Z(n20190) );
  XNOR U20319 ( .A(n20218), .B(n20231), .Z(n20230) );
  XOR U20320 ( .A(n19818), .B(n20224), .Z(n20231) );
  XNOR U20321 ( .A(n20179), .B(n19809), .Z(n20218) );
  XOR U20322 ( .A(n19732), .B(n20232), .Z(n20229) );
  XNOR U20323 ( .A(n20233), .B(n20234), .Z(n20232) );
  ANDN U20324 ( .B(n20235), .A(n20174), .Z(n20233) );
  XNOR U20325 ( .A(n20236), .B(n20237), .Z(n20202) );
  XNOR U20326 ( .A(n20223), .B(n20238), .Z(n20237) );
  XNOR U20327 ( .A(n19814), .B(n20217), .Z(n20238) );
  XOR U20328 ( .A(n20224), .B(n20239), .Z(n20217) );
  XNOR U20329 ( .A(n20240), .B(n20241), .Z(n20239) );
  NAND U20330 ( .A(n20183), .B(n19824), .Z(n20241) );
  XNOR U20331 ( .A(n20242), .B(n20240), .Z(n20224) );
  NANDN U20332 ( .A(n20185), .B(n19828), .Z(n20240) );
  XOR U20333 ( .A(n19829), .B(n19824), .Z(n19828) );
  XNOR U20334 ( .A(n20235), .B(n19699), .Z(n19824) );
  XOR U20335 ( .A(n20194), .B(n20183), .Z(n20185) );
  XNOR U20336 ( .A(n20174), .B(n20227), .Z(n20183) );
  ANDN U20337 ( .B(n19829), .A(n20194), .Z(n20242) );
  XOR U20338 ( .A(n19732), .B(n20179), .Z(n20194) );
  XNOR U20339 ( .A(n20243), .B(n20244), .Z(n20179) );
  XNOR U20340 ( .A(n20245), .B(n20246), .Z(n20244) );
  XOR U20341 ( .A(n20227), .B(n20228), .Z(n20223) );
  IV U20342 ( .A(n19699), .Z(n20228) );
  XOR U20343 ( .A(n20247), .B(n20248), .Z(n19699) );
  XNOR U20344 ( .A(n20249), .B(n20246), .Z(n20248) );
  IV U20345 ( .A(n19835), .Z(n20227) );
  XOR U20346 ( .A(n20246), .B(n20250), .Z(n19835) );
  XNOR U20347 ( .A(n20251), .B(n20252), .Z(n20236) );
  XNOR U20348 ( .A(n20253), .B(n20234), .Z(n20252) );
  OR U20349 ( .A(n19820), .B(n20173), .Z(n20234) );
  XNOR U20350 ( .A(n19732), .B(n20174), .Z(n20173) );
  IV U20351 ( .A(n20251), .Z(n20174) );
  XOR U20352 ( .A(n19818), .B(n20235), .Z(n19820) );
  IV U20353 ( .A(n19814), .Z(n20235) );
  XNOR U20354 ( .A(n20249), .B(n20243), .Z(n20254) );
  XOR U20355 ( .A(n20255), .B(n20256), .Z(n20243) );
  XOR U20356 ( .A(n20257), .B(n18195), .Z(n20256) );
  IV U20357 ( .A(n19111), .Z(n18195) );
  XNOR U20358 ( .A(n19098), .B(n20258), .Z(n19111) );
  XNOR U20359 ( .A(key[458]), .B(n20260), .Z(n20259) );
  XOR U20360 ( .A(n20247), .B(n20261), .Z(n19809) );
  XOR U20361 ( .A(n20246), .B(n20262), .Z(n20261) );
  NOR U20362 ( .A(n19818), .B(n19732), .Z(n20253) );
  XOR U20363 ( .A(n20247), .B(n20263), .Z(n19818) );
  XOR U20364 ( .A(n20246), .B(n20264), .Z(n20263) );
  XOR U20365 ( .A(n20265), .B(n20266), .Z(n20246) );
  XNOR U20366 ( .A(n18203), .B(n19131), .Z(n20266) );
  XOR U20367 ( .A(n19120), .B(n20267), .Z(n19131) );
  XNOR U20368 ( .A(n19142), .B(n18216), .Z(n18203) );
  XNOR U20369 ( .A(n20268), .B(n20269), .Z(n18216) );
  XOR U20370 ( .A(n20270), .B(n19136), .Z(n19142) );
  XOR U20371 ( .A(n19732), .B(n20271), .Z(n20265) );
  XNOR U20372 ( .A(key[462]), .B(n20272), .Z(n20271) );
  IV U20373 ( .A(n20250), .Z(n20247) );
  XOR U20374 ( .A(n20273), .B(n20274), .Z(n20250) );
  XOR U20375 ( .A(n20275), .B(n18210), .Z(n20274) );
  XOR U20376 ( .A(n19143), .B(n20276), .Z(n18210) );
  XOR U20377 ( .A(key[461]), .B(n20270), .Z(n20277) );
  XOR U20378 ( .A(n20278), .B(n20279), .Z(n20251) );
  XNOR U20379 ( .A(n20264), .B(n20262), .Z(n20279) );
  XNOR U20380 ( .A(n20280), .B(n20281), .Z(n20262) );
  XOR U20381 ( .A(n20282), .B(n18217), .Z(n20281) );
  XOR U20382 ( .A(n20283), .B(n20267), .Z(n18217) );
  XNOR U20383 ( .A(key[463]), .B(n18243), .Z(n20280) );
  XNOR U20384 ( .A(n20284), .B(n20285), .Z(n20264) );
  XOR U20385 ( .A(n18222), .B(n19125), .Z(n20285) );
  XOR U20386 ( .A(n20286), .B(n20276), .Z(n19125) );
  XNOR U20387 ( .A(n19128), .B(n20287), .Z(n18222) );
  XNOR U20388 ( .A(n18221), .B(n20288), .Z(n20284) );
  XNOR U20389 ( .A(key[460]), .B(n20289), .Z(n20288) );
  XNOR U20390 ( .A(n20268), .B(n18209), .Z(n18221) );
  XNOR U20391 ( .A(n19732), .B(n20245), .Z(n20278) );
  XOR U20392 ( .A(n20290), .B(n20291), .Z(n20245) );
  XOR U20393 ( .A(n19108), .B(n20292), .Z(n20291) );
  XOR U20394 ( .A(n20249), .B(n18230), .Z(n20292) );
  XNOR U20395 ( .A(n19135), .B(n18223), .Z(n18230) );
  IV U20396 ( .A(n20268), .Z(n19135) );
  XOR U20397 ( .A(n20293), .B(n20294), .Z(n20249) );
  XNOR U20398 ( .A(n20258), .B(n18234), .Z(n20294) );
  XNOR U20399 ( .A(n19112), .B(n20295), .Z(n18234) );
  IV U20400 ( .A(n20296), .Z(n19112) );
  XOR U20401 ( .A(n18194), .B(n20297), .Z(n20293) );
  XOR U20402 ( .A(key[457]), .B(n20298), .Z(n20297) );
  XNOR U20403 ( .A(n20286), .B(n20287), .Z(n19108) );
  XOR U20404 ( .A(n18229), .B(n20299), .Z(n20290) );
  XOR U20405 ( .A(key[459]), .B(n20300), .Z(n20299) );
  XNOR U20406 ( .A(n20301), .B(n19107), .Z(n18229) );
  XNOR U20407 ( .A(n20302), .B(n20303), .Z(n19732) );
  XOR U20408 ( .A(n18235), .B(n19134), .Z(n20303) );
  XOR U20409 ( .A(n20295), .B(n20304), .Z(n20302) );
  XOR U20410 ( .A(key[456]), .B(n20286), .Z(n20304) );
  XOR U20411 ( .A(n19700), .B(n20305), .Z(n16350) );
  XOR U20412 ( .A(n19801), .B(n19802), .Z(n20305) );
  XOR U20413 ( .A(n19886), .B(n20307), .Z(n20306) );
  NANDN U20414 ( .A(n20308), .B(n19778), .Z(n20307) );
  NOR U20415 ( .A(n19798), .B(n20309), .Z(n19886) );
  XOR U20416 ( .A(n19800), .B(n19778), .Z(n19798) );
  XNOR U20417 ( .A(n19794), .B(n20310), .Z(n19801) );
  XNOR U20418 ( .A(n20311), .B(n20312), .Z(n20310) );
  NAND U20419 ( .A(n20313), .B(n19773), .Z(n20312) );
  XNOR U20420 ( .A(n19774), .B(n20314), .Z(n19794) );
  XNOR U20421 ( .A(n20315), .B(n20316), .Z(n20314) );
  XNOR U20422 ( .A(n19793), .B(n19881), .Z(n19700) );
  XNOR U20423 ( .A(n19888), .B(n20318), .Z(n19881) );
  XOR U20424 ( .A(n20319), .B(n19770), .Z(n20318) );
  OR U20425 ( .A(n20320), .B(n20321), .Z(n19770) );
  ANDN U20426 ( .B(n20322), .A(n20323), .Z(n20319) );
  XNOR U20427 ( .A(n20324), .B(n19890), .Z(n19888) );
  NANDN U20428 ( .A(n20325), .B(n20326), .Z(n19890) );
  AND U20429 ( .A(n20327), .B(n20328), .Z(n20324) );
  XOR U20430 ( .A(n19774), .B(n20329), .Z(n19793) );
  XNOR U20431 ( .A(n20311), .B(n20330), .Z(n20329) );
  NANDN U20432 ( .A(n20331), .B(n20322), .Z(n20330) );
  OR U20433 ( .A(n20320), .B(n20332), .Z(n20311) );
  XNOR U20434 ( .A(n19773), .B(n20322), .Z(n20320) );
  XOR U20435 ( .A(n20333), .B(n20315), .Z(n19774) );
  OR U20436 ( .A(n20334), .B(n20325), .Z(n20315) );
  XOR U20437 ( .A(n20328), .B(n19892), .Z(n20325) );
  XNOR U20438 ( .A(n20322), .B(n19778), .Z(n19892) );
  XOR U20439 ( .A(n20335), .B(n20336), .Z(n19778) );
  NANDN U20440 ( .A(n20337), .B(n20338), .Z(n20336) );
  XOR U20441 ( .A(n20339), .B(n20340), .Z(n20322) );
  NANDN U20442 ( .A(n20337), .B(n20341), .Z(n20340) );
  ANDN U20443 ( .B(n20328), .A(n20342), .Z(n20333) );
  XNOR U20444 ( .A(n19800), .B(n19773), .Z(n20328) );
  XNOR U20445 ( .A(n20343), .B(n20339), .Z(n19773) );
  NANDN U20446 ( .A(n20344), .B(n20345), .Z(n20339) );
  XOR U20447 ( .A(n20341), .B(n20346), .Z(n20345) );
  ANDN U20448 ( .B(n20346), .A(n20347), .Z(n20343) );
  NANDN U20449 ( .A(n20344), .B(n20349), .Z(n20335) );
  XOR U20450 ( .A(n20350), .B(n20338), .Z(n20349) );
  XNOR U20451 ( .A(n20351), .B(n20352), .Z(n20337) );
  XOR U20452 ( .A(n20353), .B(n20354), .Z(n20352) );
  XNOR U20453 ( .A(n20355), .B(n20356), .Z(n20351) );
  XNOR U20454 ( .A(n20357), .B(n20358), .Z(n20356) );
  ANDN U20455 ( .B(n20350), .A(n20354), .Z(n20357) );
  ANDN U20456 ( .B(n20350), .A(n20347), .Z(n20348) );
  XNOR U20457 ( .A(n20353), .B(n20359), .Z(n20347) );
  XOR U20458 ( .A(n20360), .B(n20358), .Z(n20359) );
  NAND U20459 ( .A(n20361), .B(n20362), .Z(n20358) );
  XNOR U20460 ( .A(n20355), .B(n20338), .Z(n20362) );
  IV U20461 ( .A(n20350), .Z(n20355) );
  XNOR U20462 ( .A(n20341), .B(n20354), .Z(n20361) );
  IV U20463 ( .A(n20346), .Z(n20354) );
  XOR U20464 ( .A(n20363), .B(n20364), .Z(n20346) );
  XNOR U20465 ( .A(n20365), .B(n20366), .Z(n20364) );
  XNOR U20466 ( .A(n20367), .B(n20368), .Z(n20363) );
  ANDN U20467 ( .B(n19887), .A(n19799), .Z(n20367) );
  AND U20468 ( .A(n20338), .B(n20341), .Z(n20360) );
  XNOR U20469 ( .A(n20338), .B(n20341), .Z(n20353) );
  XNOR U20470 ( .A(n20369), .B(n20370), .Z(n20341) );
  XNOR U20471 ( .A(n20371), .B(n20366), .Z(n20370) );
  XOR U20472 ( .A(n20372), .B(n20373), .Z(n20369) );
  XNOR U20473 ( .A(n20374), .B(n20368), .Z(n20373) );
  OR U20474 ( .A(n19797), .B(n20309), .Z(n20368) );
  XNOR U20475 ( .A(n19887), .B(n20414), .Z(n20309) );
  XNOR U20476 ( .A(n19799), .B(n19779), .Z(n19797) );
  ANDN U20477 ( .B(n20375), .A(n20308), .Z(n20374) );
  XNOR U20478 ( .A(n20376), .B(n20377), .Z(n20338) );
  XNOR U20479 ( .A(n20366), .B(n20378), .Z(n20377) );
  XNOR U20480 ( .A(n20313), .B(n20372), .Z(n20378) );
  XNOR U20481 ( .A(n19799), .B(n19887), .Z(n20366) );
  XOR U20482 ( .A(n19772), .B(n20379), .Z(n20376) );
  XNOR U20483 ( .A(n20380), .B(n20381), .Z(n20379) );
  ANDN U20484 ( .B(n20382), .A(n20323), .Z(n20380) );
  XNOR U20485 ( .A(n20383), .B(n20384), .Z(n20350) );
  XNOR U20486 ( .A(n20371), .B(n20385), .Z(n20384) );
  XNOR U20487 ( .A(n20386), .B(n20365), .Z(n20385) );
  XOR U20488 ( .A(n20372), .B(n20387), .Z(n20365) );
  XNOR U20489 ( .A(n20388), .B(n20389), .Z(n20387) );
  NANDN U20490 ( .A(n20317), .B(n19893), .Z(n20389) );
  XNOR U20491 ( .A(n20390), .B(n20388), .Z(n20372) );
  NANDN U20492 ( .A(n20334), .B(n20326), .Z(n20388) );
  XOR U20493 ( .A(n20327), .B(n19893), .Z(n20326) );
  XNOR U20494 ( .A(n20323), .B(n20414), .Z(n19893) );
  XOR U20495 ( .A(n20391), .B(n20317), .Z(n20334) );
  XNOR U20496 ( .A(n20375), .B(n20382), .Z(n20317) );
  IV U20497 ( .A(n19779), .Z(n20375) );
  ANDN U20498 ( .B(n20327), .A(n20342), .Z(n20390) );
  IV U20499 ( .A(n20391), .Z(n20342) );
  XOR U20500 ( .A(n20392), .B(n20313), .Z(n20391) );
  XNOR U20501 ( .A(n19772), .B(n19887), .Z(n20327) );
  XNOR U20502 ( .A(n20393), .B(n20394), .Z(n19887) );
  XNOR U20503 ( .A(n20395), .B(n20396), .Z(n20394) );
  XOR U20504 ( .A(n19779), .B(n20308), .Z(n20371) );
  XOR U20505 ( .A(n20397), .B(n20395), .Z(n20308) );
  XOR U20506 ( .A(n20398), .B(n20399), .Z(n19779) );
  XOR U20507 ( .A(n20400), .B(n20395), .Z(n20399) );
  XNOR U20508 ( .A(n20331), .B(n20401), .Z(n20383) );
  XNOR U20509 ( .A(n20402), .B(n20381), .Z(n20401) );
  OR U20510 ( .A(n20332), .B(n20321), .Z(n20381) );
  XNOR U20511 ( .A(n19772), .B(n20323), .Z(n20321) );
  IV U20512 ( .A(n20386), .Z(n20323) );
  XOR U20513 ( .A(n20403), .B(n20404), .Z(n20386) );
  XNOR U20514 ( .A(n20405), .B(n20393), .Z(n20404) );
  XOR U20515 ( .A(n20406), .B(n20407), .Z(n20393) );
  XOR U20516 ( .A(n19547), .B(n20408), .Z(n20407) );
  XNOR U20517 ( .A(n20398), .B(n18361), .Z(n20408) );
  XNOR U20518 ( .A(n18383), .B(n19515), .Z(n18361) );
  XOR U20519 ( .A(n20409), .B(n20410), .Z(n19547) );
  XNOR U20520 ( .A(n20411), .B(n20412), .Z(n20406) );
  XOR U20521 ( .A(key[499]), .B(n19555), .Z(n20412) );
  XNOR U20522 ( .A(n19772), .B(n20413), .Z(n20403) );
  XNOR U20523 ( .A(n20313), .B(n20382), .Z(n20332) );
  IV U20524 ( .A(n20331), .Z(n20382) );
  ANDN U20525 ( .B(n20313), .A(n19772), .Z(n20402) );
  XOR U20526 ( .A(n20405), .B(n20414), .Z(n20313) );
  XOR U20527 ( .A(n20415), .B(n19514), .Z(n20405) );
  XNOR U20528 ( .A(n20416), .B(n20417), .Z(n19514) );
  XNOR U20529 ( .A(n20418), .B(n18348), .Z(n20417) );
  XNOR U20530 ( .A(n20419), .B(n20420), .Z(n20416) );
  XNOR U20531 ( .A(n18345), .B(n20421), .Z(n20415) );
  XOR U20532 ( .A(n18383), .B(n19526), .Z(n18345) );
  XNOR U20533 ( .A(n20396), .B(n20422), .Z(n20331) );
  XOR U20534 ( .A(n19799), .B(n20398), .Z(n20422) );
  XNOR U20535 ( .A(n20423), .B(n20424), .Z(n20398) );
  XOR U20536 ( .A(n18376), .B(n19559), .Z(n20424) );
  XNOR U20537 ( .A(key[497]), .B(n19552), .Z(n20423) );
  IV U20538 ( .A(n20392), .Z(n19799) );
  XOR U20539 ( .A(n20413), .B(n20414), .Z(n20392) );
  XNOR U20540 ( .A(n20397), .B(n20395), .Z(n20414) );
  XOR U20541 ( .A(n20425), .B(n20426), .Z(n20395) );
  XNOR U20542 ( .A(n19772), .B(n19541), .Z(n20426) );
  XOR U20543 ( .A(n20427), .B(n20428), .Z(n19541) );
  XNOR U20544 ( .A(n20429), .B(n20430), .Z(n19772) );
  XNOR U20545 ( .A(n18365), .B(n18382), .Z(n20430) );
  XNOR U20546 ( .A(n20419), .B(n19558), .Z(n18382) );
  IV U20547 ( .A(n20409), .Z(n20419) );
  XOR U20548 ( .A(key[496]), .B(n20431), .Z(n20429) );
  XNOR U20549 ( .A(n18353), .B(n20432), .Z(n20425) );
  XNOR U20550 ( .A(key[502]), .B(n19528), .Z(n20432) );
  XNOR U20551 ( .A(n18383), .B(n19532), .Z(n18353) );
  IV U20552 ( .A(n20400), .Z(n20397) );
  XNOR U20553 ( .A(n20433), .B(n20434), .Z(n20400) );
  XNOR U20554 ( .A(n20420), .B(n19525), .Z(n20434) );
  XOR U20555 ( .A(n20435), .B(n18330), .Z(n19525) );
  XNOR U20556 ( .A(key[501]), .B(n20436), .Z(n20433) );
  XOR U20557 ( .A(n20437), .B(n20438), .Z(n20413) );
  XNOR U20558 ( .A(n20428), .B(n19531), .Z(n20438) );
  XOR U20559 ( .A(n20409), .B(n20440), .Z(n20428) );
  XNOR U20560 ( .A(key[503]), .B(n18383), .Z(n20437) );
  XOR U20561 ( .A(n20441), .B(n20442), .Z(n20396) );
  XNOR U20562 ( .A(n19536), .B(n18360), .Z(n20442) );
  XNOR U20563 ( .A(key[498]), .B(n19550), .Z(n20441) );
  XNOR U20564 ( .A(key[640]), .B(n13385), .Z(n17747) );
  XOR U20565 ( .A(n17611), .B(n17559), .Z(n13385) );
  XNOR U20566 ( .A(n17581), .B(n20443), .Z(n17559) );
  XNOR U20567 ( .A(n20444), .B(n17744), .Z(n20443) );
  XOR U20568 ( .A(n17720), .B(n17565), .Z(n17718) );
  ANDN U20569 ( .B(n17720), .A(n20446), .Z(n20444) );
  XNOR U20570 ( .A(n17742), .B(n20447), .Z(n17581) );
  XNOR U20571 ( .A(n20448), .B(n20449), .Z(n20447) );
  NANDN U20572 ( .A(n17735), .B(n20450), .Z(n20449) );
  XOR U20573 ( .A(n17742), .B(n20451), .Z(n17611) );
  XOR U20574 ( .A(n20452), .B(n17583), .Z(n20451) );
  OR U20575 ( .A(n20453), .B(n17730), .Z(n17583) );
  XNOR U20576 ( .A(n17585), .B(n17725), .Z(n17730) );
  NOR U20577 ( .A(n20454), .B(n17725), .Z(n20452) );
  XOR U20578 ( .A(n20455), .B(n20448), .Z(n17742) );
  OR U20579 ( .A(n17738), .B(n20456), .Z(n20448) );
  XOR U20580 ( .A(n20457), .B(n17735), .Z(n17738) );
  XOR U20581 ( .A(n17725), .B(n17565), .Z(n17735) );
  XOR U20582 ( .A(n20458), .B(n20459), .Z(n17565) );
  NANDN U20583 ( .A(n20460), .B(n20461), .Z(n20459) );
  XNOR U20584 ( .A(n20462), .B(n20463), .Z(n17725) );
  OR U20585 ( .A(n20460), .B(n20464), .Z(n20463) );
  ANDN U20586 ( .B(n20457), .A(n20465), .Z(n20455) );
  IV U20587 ( .A(n17741), .Z(n20457) );
  XOR U20588 ( .A(n17585), .B(n17720), .Z(n17741) );
  XNOR U20589 ( .A(n20466), .B(n20458), .Z(n17720) );
  NANDN U20590 ( .A(n20467), .B(n20468), .Z(n20458) );
  ANDN U20591 ( .B(n20469), .A(n20470), .Z(n20466) );
  NANDN U20592 ( .A(n20467), .B(n20472), .Z(n20462) );
  XOR U20593 ( .A(n20473), .B(n20460), .Z(n20467) );
  XNOR U20594 ( .A(n20474), .B(n20475), .Z(n20460) );
  XOR U20595 ( .A(n20476), .B(n20469), .Z(n20475) );
  XNOR U20596 ( .A(n20477), .B(n20478), .Z(n20474) );
  XNOR U20597 ( .A(n20479), .B(n20480), .Z(n20478) );
  ANDN U20598 ( .B(n20469), .A(n20481), .Z(n20479) );
  IV U20599 ( .A(n20482), .Z(n20469) );
  ANDN U20600 ( .B(n20473), .A(n20481), .Z(n20471) );
  IV U20601 ( .A(n20477), .Z(n20481) );
  IV U20602 ( .A(n20470), .Z(n20473) );
  XNOR U20603 ( .A(n20476), .B(n20483), .Z(n20470) );
  XOR U20604 ( .A(n20484), .B(n20480), .Z(n20483) );
  NAND U20605 ( .A(n20472), .B(n20468), .Z(n20480) );
  XNOR U20606 ( .A(n20461), .B(n20482), .Z(n20468) );
  XOR U20607 ( .A(n20485), .B(n20486), .Z(n20482) );
  XOR U20608 ( .A(n20487), .B(n20488), .Z(n20486) );
  XNOR U20609 ( .A(n17726), .B(n20489), .Z(n20488) );
  XNOR U20610 ( .A(n20490), .B(n20491), .Z(n20485) );
  XNOR U20611 ( .A(n20492), .B(n20493), .Z(n20491) );
  ANDN U20612 ( .B(n20494), .A(n17586), .Z(n20492) );
  XNOR U20613 ( .A(n20477), .B(n20464), .Z(n20472) );
  XOR U20614 ( .A(n20495), .B(n20496), .Z(n20477) );
  XNOR U20615 ( .A(n20497), .B(n20489), .Z(n20496) );
  XOR U20616 ( .A(n20498), .B(n20499), .Z(n20489) );
  XNOR U20617 ( .A(n20500), .B(n20501), .Z(n20499) );
  NAND U20618 ( .A(n20450), .B(n17736), .Z(n20501) );
  XNOR U20619 ( .A(n20502), .B(n20503), .Z(n20495) );
  ANDN U20620 ( .B(n20504), .A(n20446), .Z(n20502) );
  ANDN U20621 ( .B(n20461), .A(n20464), .Z(n20484) );
  XOR U20622 ( .A(n20464), .B(n20461), .Z(n20476) );
  XNOR U20623 ( .A(n20505), .B(n20506), .Z(n20461) );
  XNOR U20624 ( .A(n20498), .B(n20507), .Z(n20506) );
  XOR U20625 ( .A(n20497), .B(n17729), .Z(n20507) );
  XOR U20626 ( .A(n17586), .B(n20508), .Z(n20505) );
  XNOR U20627 ( .A(n20509), .B(n20493), .Z(n20508) );
  OR U20628 ( .A(n17731), .B(n20453), .Z(n20493) );
  XNOR U20629 ( .A(n17586), .B(n20454), .Z(n20453) );
  XOR U20630 ( .A(n17729), .B(n17726), .Z(n17731) );
  ANDN U20631 ( .B(n17726), .A(n20454), .Z(n20509) );
  XOR U20632 ( .A(n20510), .B(n20511), .Z(n20464) );
  XOR U20633 ( .A(n20498), .B(n20487), .Z(n20511) );
  XOR U20634 ( .A(n17746), .B(n17566), .Z(n20487) );
  XOR U20635 ( .A(n20512), .B(n20500), .Z(n20498) );
  NANDN U20636 ( .A(n20456), .B(n17739), .Z(n20500) );
  XOR U20637 ( .A(n17740), .B(n17736), .Z(n17739) );
  XNOR U20638 ( .A(n20504), .B(n20513), .Z(n17726) );
  XOR U20639 ( .A(n20514), .B(n20515), .Z(n20513) );
  XOR U20640 ( .A(n20465), .B(n20450), .Z(n20456) );
  XNOR U20641 ( .A(n20454), .B(n17746), .Z(n20450) );
  IV U20642 ( .A(n20490), .Z(n20454) );
  XOR U20643 ( .A(n20516), .B(n20517), .Z(n20490) );
  XOR U20644 ( .A(n20518), .B(n20519), .Z(n20517) );
  XNOR U20645 ( .A(n17586), .B(n20520), .Z(n20516) );
  ANDN U20646 ( .B(n17740), .A(n20465), .Z(n20512) );
  XNOR U20647 ( .A(n17586), .B(n20446), .Z(n20465) );
  XOR U20648 ( .A(n20504), .B(n20494), .Z(n17740) );
  IV U20649 ( .A(n17729), .Z(n20494) );
  XOR U20650 ( .A(n20521), .B(n20522), .Z(n17729) );
  XOR U20651 ( .A(n20523), .B(n20519), .Z(n20522) );
  XNOR U20652 ( .A(n20524), .B(n20525), .Z(n20519) );
  XNOR U20653 ( .A(n17127), .B(n17126), .Z(n20525) );
  XOR U20654 ( .A(n15338), .B(n16050), .Z(n17126) );
  XNOR U20655 ( .A(n20526), .B(n15309), .Z(n15338) );
  XNOR U20656 ( .A(n20527), .B(n16076), .Z(n17127) );
  XNOR U20657 ( .A(n20528), .B(n20529), .Z(n16076) );
  XNOR U20658 ( .A(n20530), .B(n20531), .Z(n20529) );
  XOR U20659 ( .A(n20532), .B(n20533), .Z(n20528) );
  XOR U20660 ( .A(n20534), .B(n20535), .Z(n20533) );
  ANDN U20661 ( .B(n20536), .A(n20537), .Z(n20535) );
  XNOR U20662 ( .A(n15335), .B(n20538), .Z(n20524) );
  XOR U20663 ( .A(key[588]), .B(n17113), .Z(n20538) );
  XOR U20664 ( .A(n20539), .B(n16032), .Z(n17113) );
  XOR U20665 ( .A(n15331), .B(n16074), .Z(n15335) );
  IV U20666 ( .A(n17721), .Z(n20504) );
  XOR U20667 ( .A(n20497), .B(n20540), .Z(n20510) );
  XNOR U20668 ( .A(n20541), .B(n20503), .Z(n20540) );
  OR U20669 ( .A(n17719), .B(n20445), .Z(n20503) );
  XNOR U20670 ( .A(n20542), .B(n17746), .Z(n20445) );
  XNOR U20671 ( .A(n17721), .B(n17566), .Z(n17719) );
  ANDN U20672 ( .B(n17746), .A(n17566), .Z(n20541) );
  XOR U20673 ( .A(n20521), .B(n20543), .Z(n17566) );
  XOR U20674 ( .A(n20523), .B(n20521), .Z(n17746) );
  XNOR U20675 ( .A(n20446), .B(n17721), .Z(n20497) );
  XOR U20676 ( .A(n20521), .B(n20544), .Z(n17721) );
  XNOR U20677 ( .A(n20523), .B(n20518), .Z(n20544) );
  XOR U20678 ( .A(n20545), .B(n20546), .Z(n20518) );
  XNOR U20679 ( .A(n16064), .B(n17122), .Z(n20546) );
  XOR U20680 ( .A(n16071), .B(n16054), .Z(n17122) );
  XOR U20681 ( .A(n20547), .B(n20548), .Z(n16071) );
  XNOR U20682 ( .A(n20549), .B(n20550), .Z(n20548) );
  XNOR U20683 ( .A(n20527), .B(n15331), .Z(n16064) );
  IV U20684 ( .A(n15356), .Z(n20527) );
  XNOR U20685 ( .A(key[591]), .B(n16055), .Z(n20545) );
  XOR U20686 ( .A(n20551), .B(n20552), .Z(n16055) );
  XOR U20687 ( .A(n20553), .B(n20554), .Z(n20552) );
  XNOR U20688 ( .A(n20555), .B(n20556), .Z(n20521) );
  XNOR U20689 ( .A(n16068), .B(n17140), .Z(n20556) );
  XNOR U20690 ( .A(n15324), .B(n16074), .Z(n17140) );
  XNOR U20691 ( .A(n20557), .B(n20558), .Z(n16074) );
  XOR U20692 ( .A(n20559), .B(n20560), .Z(n20558) );
  XOR U20693 ( .A(n20561), .B(n20562), .Z(n20557) );
  XNOR U20694 ( .A(n20563), .B(n20564), .Z(n20562) );
  ANDN U20695 ( .B(n20565), .A(n20566), .Z(n20563) );
  XOR U20696 ( .A(n20567), .B(n20568), .Z(n15324) );
  XNOR U20697 ( .A(n20569), .B(n20550), .Z(n20568) );
  XNOR U20698 ( .A(n20570), .B(n20571), .Z(n20550) );
  XNOR U20699 ( .A(n20572), .B(n20573), .Z(n20571) );
  OR U20700 ( .A(n20574), .B(n20575), .Z(n20573) );
  XNOR U20701 ( .A(n20526), .B(n20576), .Z(n20567) );
  XOR U20702 ( .A(n20577), .B(n20578), .Z(n20576) );
  ANDN U20703 ( .B(n20579), .A(n20580), .Z(n20578) );
  XOR U20704 ( .A(n16075), .B(n20581), .Z(n20555) );
  XNOR U20705 ( .A(key[589]), .B(n17137), .Z(n20581) );
  XNOR U20706 ( .A(n20582), .B(n20583), .Z(n17137) );
  XNOR U20707 ( .A(n20584), .B(n20585), .Z(n16075) );
  XOR U20708 ( .A(n20586), .B(n20554), .Z(n20585) );
  XNOR U20709 ( .A(n20587), .B(n20588), .Z(n20554) );
  XNOR U20710 ( .A(n20589), .B(n20590), .Z(n20588) );
  NANDN U20711 ( .A(n20591), .B(n20592), .Z(n20590) );
  XNOR U20712 ( .A(n20539), .B(n20593), .Z(n20584) );
  XOR U20713 ( .A(n20594), .B(n20595), .Z(n20593) );
  ANDN U20714 ( .B(n20596), .A(n20597), .Z(n20595) );
  IV U20715 ( .A(n20542), .Z(n20446) );
  XNOR U20716 ( .A(n20515), .B(n20598), .Z(n20542) );
  XOR U20717 ( .A(n20599), .B(n20600), .Z(n20523) );
  XNOR U20718 ( .A(n17586), .B(n17135), .Z(n20600) );
  XOR U20719 ( .A(n15323), .B(n17121), .Z(n17135) );
  XNOR U20720 ( .A(n15356), .B(n16056), .Z(n17121) );
  XNOR U20721 ( .A(n20601), .B(n20602), .Z(n16056) );
  XOR U20722 ( .A(n20603), .B(n20531), .Z(n20602) );
  XNOR U20723 ( .A(n20604), .B(n20605), .Z(n20531) );
  XNOR U20724 ( .A(n20606), .B(n20607), .Z(n20605) );
  NANDN U20725 ( .A(n20608), .B(n20609), .Z(n20607) );
  XOR U20726 ( .A(n20583), .B(n20610), .Z(n20601) );
  XNOR U20727 ( .A(n15318), .B(n16068), .Z(n15323) );
  XOR U20728 ( .A(n20611), .B(n20612), .Z(n16068) );
  IV U20729 ( .A(n16079), .Z(n15318) );
  XNOR U20730 ( .A(n20549), .B(n20613), .Z(n16079) );
  XNOR U20731 ( .A(n20614), .B(n20615), .Z(n17586) );
  XOR U20732 ( .A(n17116), .B(n20616), .Z(n20615) );
  XNOR U20733 ( .A(n20617), .B(n20618), .Z(n17116) );
  XOR U20734 ( .A(n20583), .B(n20619), .Z(n20618) );
  XOR U20735 ( .A(n16034), .B(n20622), .Z(n20614) );
  XOR U20736 ( .A(key[584]), .B(n15354), .Z(n20622) );
  IV U20737 ( .A(n16057), .Z(n15354) );
  XOR U20738 ( .A(n16067), .B(n17134), .Z(n16057) );
  IV U20739 ( .A(n16036), .Z(n17134) );
  XOR U20740 ( .A(n20623), .B(n20526), .Z(n16036) );
  XNOR U20741 ( .A(n20570), .B(n20624), .Z(n20526) );
  XOR U20742 ( .A(n20625), .B(n20626), .Z(n20624) );
  ANDN U20743 ( .B(n20627), .A(n20628), .Z(n20625) );
  XOR U20744 ( .A(n20629), .B(n20630), .Z(n20570) );
  XNOR U20745 ( .A(n20631), .B(n20632), .Z(n20630) );
  NANDN U20746 ( .A(n20633), .B(n20634), .Z(n20632) );
  XOR U20747 ( .A(n20539), .B(n20635), .Z(n16067) );
  XNOR U20748 ( .A(n20587), .B(n20636), .Z(n20539) );
  XOR U20749 ( .A(n20637), .B(n20638), .Z(n20636) );
  NOR U20750 ( .A(n20639), .B(n20640), .Z(n20637) );
  XOR U20751 ( .A(n20641), .B(n20642), .Z(n20587) );
  XNOR U20752 ( .A(n20643), .B(n20644), .Z(n20642) );
  NAND U20753 ( .A(n20645), .B(n20646), .Z(n20644) );
  XNOR U20754 ( .A(n15317), .B(n20647), .Z(n20599) );
  XOR U20755 ( .A(key[590]), .B(n16077), .Z(n20647) );
  XOR U20756 ( .A(n20648), .B(n20649), .Z(n16077) );
  XOR U20757 ( .A(n15331), .B(n16054), .Z(n15317) );
  XNOR U20758 ( .A(n20650), .B(n20651), .Z(n16054) );
  XNOR U20759 ( .A(n20652), .B(n20560), .Z(n20651) );
  XNOR U20760 ( .A(n20653), .B(n20654), .Z(n20560) );
  XNOR U20761 ( .A(n20655), .B(n20656), .Z(n20654) );
  OR U20762 ( .A(n20657), .B(n20658), .Z(n20656) );
  XNOR U20763 ( .A(n20612), .B(n20659), .Z(n20650) );
  XOR U20764 ( .A(n20660), .B(n20661), .Z(n20520) );
  XNOR U20765 ( .A(n17112), .B(n20662), .Z(n20661) );
  XOR U20766 ( .A(n15308), .B(n20514), .Z(n20662) );
  XNOR U20767 ( .A(n20663), .B(n20664), .Z(n20514) );
  XNOR U20768 ( .A(n16040), .B(n17101), .Z(n20664) );
  XOR U20769 ( .A(n17133), .B(n20665), .Z(n20663) );
  XOR U20770 ( .A(key[585]), .B(n15355), .Z(n20665) );
  XOR U20771 ( .A(n15348), .B(n16034), .Z(n15355) );
  XOR U20772 ( .A(n20652), .B(n20666), .Z(n16034) );
  XOR U20773 ( .A(n20612), .B(n20659), .Z(n20666) );
  XOR U20774 ( .A(n20667), .B(n20668), .Z(n20612) );
  IV U20775 ( .A(n16065), .Z(n15348) );
  XNOR U20776 ( .A(n20549), .B(n20669), .Z(n16065) );
  XNOR U20777 ( .A(n20670), .B(n20671), .Z(n20669) );
  XOR U20778 ( .A(n20623), .B(n20672), .Z(n20549) );
  IV U20779 ( .A(n16063), .Z(n17133) );
  XOR U20780 ( .A(n20553), .B(n20673), .Z(n16063) );
  XNOR U20781 ( .A(n20674), .B(n20675), .Z(n20673) );
  IV U20782 ( .A(n20648), .Z(n20553) );
  XOR U20783 ( .A(n20635), .B(n20676), .Z(n20648) );
  XOR U20784 ( .A(n16042), .B(n16028), .Z(n15308) );
  IV U20785 ( .A(n15349), .Z(n16042) );
  XNOR U20786 ( .A(n20547), .B(n20677), .Z(n15349) );
  XOR U20787 ( .A(n20672), .B(n20613), .Z(n20677) );
  XNOR U20788 ( .A(n20678), .B(n20679), .Z(n20613) );
  XNOR U20789 ( .A(n20680), .B(n20577), .Z(n20679) );
  ANDN U20790 ( .B(n20681), .A(n20682), .Z(n20577) );
  ANDN U20791 ( .B(n20627), .A(n20683), .Z(n20680) );
  XOR U20792 ( .A(n20569), .B(n20684), .Z(n20672) );
  XNOR U20793 ( .A(n20685), .B(n20686), .Z(n20684) );
  NANDN U20794 ( .A(n20687), .B(n20688), .Z(n20686) );
  XOR U20795 ( .A(n20670), .B(n20671), .Z(n20547) );
  XNOR U20796 ( .A(n20685), .B(n20690), .Z(n20689) );
  OR U20797 ( .A(n20574), .B(n20691), .Z(n20690) );
  OR U20798 ( .A(n20692), .B(n20693), .Z(n20685) );
  XNOR U20799 ( .A(n20569), .B(n20694), .Z(n20678) );
  XNOR U20800 ( .A(n20695), .B(n20696), .Z(n20694) );
  NANDN U20801 ( .A(n20633), .B(n20697), .Z(n20696) );
  XOR U20802 ( .A(n20698), .B(n20695), .Z(n20569) );
  NANDN U20803 ( .A(n20699), .B(n20700), .Z(n20695) );
  ANDN U20804 ( .B(n20701), .A(n20702), .Z(n20698) );
  XOR U20805 ( .A(n15356), .B(n16048), .Z(n17112) );
  XNOR U20806 ( .A(n20532), .B(n17101), .Z(n16048) );
  XNOR U20807 ( .A(n20620), .B(n20610), .Z(n17101) );
  XOR U20808 ( .A(n20620), .B(n20532), .Z(n15356) );
  XOR U20809 ( .A(n20604), .B(n20703), .Z(n20532) );
  XNOR U20810 ( .A(n20704), .B(n20705), .Z(n20703) );
  NANDN U20811 ( .A(n20706), .B(n20707), .Z(n20705) );
  XNOR U20812 ( .A(n20708), .B(n20709), .Z(n20604) );
  XNOR U20813 ( .A(n20710), .B(n20711), .Z(n20709) );
  NAND U20814 ( .A(n20712), .B(n20713), .Z(n20711) );
  XOR U20815 ( .A(n20708), .B(n20714), .Z(n20620) );
  XOR U20816 ( .A(n20715), .B(n20606), .Z(n20714) );
  OR U20817 ( .A(n20716), .B(n20717), .Z(n20606) );
  NOR U20818 ( .A(n20718), .B(n20719), .Z(n20715) );
  XNOR U20819 ( .A(n15341), .B(n20720), .Z(n20660) );
  XOR U20820 ( .A(key[587]), .B(n17103), .Z(n20720) );
  XNOR U20821 ( .A(n20551), .B(n20721), .Z(n17103) );
  XOR U20822 ( .A(n20676), .B(n20649), .Z(n20721) );
  XNOR U20823 ( .A(n20722), .B(n20723), .Z(n20649) );
  XNOR U20824 ( .A(n20724), .B(n20594), .Z(n20723) );
  ANDN U20825 ( .B(n20725), .A(n20726), .Z(n20594) );
  NOR U20826 ( .A(n20727), .B(n20640), .Z(n20724) );
  XNOR U20827 ( .A(n20586), .B(n20728), .Z(n20676) );
  XNOR U20828 ( .A(n20729), .B(n20730), .Z(n20728) );
  NANDN U20829 ( .A(n20731), .B(n20732), .Z(n20730) );
  XOR U20830 ( .A(n20674), .B(n20675), .Z(n20551) );
  XNOR U20831 ( .A(n20729), .B(n20734), .Z(n20733) );
  NANDN U20832 ( .A(n20735), .B(n20592), .Z(n20734) );
  OR U20833 ( .A(n20736), .B(n20737), .Z(n20729) );
  XOR U20834 ( .A(n20586), .B(n20738), .Z(n20722) );
  XNOR U20835 ( .A(n20739), .B(n20740), .Z(n20738) );
  NAND U20836 ( .A(n20741), .B(n20645), .Z(n20740) );
  XNOR U20837 ( .A(n20742), .B(n20739), .Z(n20586) );
  NANDN U20838 ( .A(n20743), .B(n20744), .Z(n20739) );
  ANDN U20839 ( .B(n20745), .A(n20746), .Z(n20742) );
  XNOR U20840 ( .A(n15331), .B(n16050), .Z(n15341) );
  XNOR U20841 ( .A(n16040), .B(n20559), .Z(n16050) );
  IV U20842 ( .A(n20616), .Z(n15331) );
  XOR U20843 ( .A(n20667), .B(n20559), .Z(n20616) );
  XOR U20844 ( .A(n20653), .B(n20747), .Z(n20559) );
  XOR U20845 ( .A(n20748), .B(n20749), .Z(n20747) );
  ANDN U20846 ( .B(n20750), .A(n20751), .Z(n20748) );
  XNOR U20847 ( .A(n20752), .B(n20753), .Z(n20653) );
  XNOR U20848 ( .A(n20754), .B(n20755), .Z(n20753) );
  NANDN U20849 ( .A(n20756), .B(n20757), .Z(n20755) );
  XOR U20850 ( .A(n20758), .B(n20759), .Z(n20515) );
  XOR U20851 ( .A(n16032), .B(n16028), .Z(n20759) );
  XNOR U20852 ( .A(n20760), .B(n20761), .Z(n16028) );
  XNOR U20853 ( .A(n20652), .B(n20611), .Z(n20761) );
  XNOR U20854 ( .A(n20762), .B(n20763), .Z(n20611) );
  XNOR U20855 ( .A(n20564), .B(n20764), .Z(n20763) );
  NANDN U20856 ( .A(n20765), .B(n20750), .Z(n20764) );
  NANDN U20857 ( .A(n20766), .B(n20767), .Z(n20564) );
  XNOR U20858 ( .A(n20769), .B(n20770), .Z(n20768) );
  OR U20859 ( .A(n20657), .B(n20771), .Z(n20770) );
  XOR U20860 ( .A(n20561), .B(n20772), .Z(n20762) );
  XNOR U20861 ( .A(n20773), .B(n20774), .Z(n20772) );
  NANDN U20862 ( .A(n20756), .B(n20775), .Z(n20774) );
  XNOR U20863 ( .A(n20668), .B(n20659), .Z(n20760) );
  XOR U20864 ( .A(n20777), .B(n20769), .Z(n20776) );
  OR U20865 ( .A(n20778), .B(n20779), .Z(n20769) );
  AND U20866 ( .A(n20780), .B(n20781), .Z(n20777) );
  XNOR U20867 ( .A(n20782), .B(n20773), .Z(n20561) );
  NANDN U20868 ( .A(n20783), .B(n20784), .Z(n20773) );
  ANDN U20869 ( .B(n20785), .A(n20786), .Z(n20782) );
  XOR U20870 ( .A(n20635), .B(n20674), .Z(n16032) );
  XNOR U20871 ( .A(n20641), .B(n20787), .Z(n20674) );
  XNOR U20872 ( .A(n20638), .B(n20788), .Z(n20787) );
  NANDN U20873 ( .A(n20789), .B(n20596), .Z(n20788) );
  XNOR U20874 ( .A(n20640), .B(n20596), .Z(n20725) );
  XOR U20875 ( .A(n20792), .B(n20589), .Z(n20791) );
  OR U20876 ( .A(n20736), .B(n20793), .Z(n20589) );
  XNOR U20877 ( .A(n20592), .B(n20732), .Z(n20736) );
  ANDN U20878 ( .B(n20732), .A(n20794), .Z(n20792) );
  XNOR U20879 ( .A(n20795), .B(n20643), .Z(n20641) );
  OR U20880 ( .A(n20743), .B(n20796), .Z(n20643) );
  XNOR U20881 ( .A(n20797), .B(n20645), .Z(n20743) );
  XOR U20882 ( .A(n20732), .B(n20596), .Z(n20645) );
  XOR U20883 ( .A(n20798), .B(n20799), .Z(n20596) );
  NANDN U20884 ( .A(n20800), .B(n20801), .Z(n20799) );
  XOR U20885 ( .A(n20802), .B(n20803), .Z(n20732) );
  NANDN U20886 ( .A(n20800), .B(n20804), .Z(n20803) );
  ANDN U20887 ( .B(n20797), .A(n20805), .Z(n20795) );
  IV U20888 ( .A(n20746), .Z(n20797) );
  XOR U20889 ( .A(n20640), .B(n20592), .Z(n20746) );
  XNOR U20890 ( .A(n20806), .B(n20802), .Z(n20592) );
  NANDN U20891 ( .A(n20807), .B(n20808), .Z(n20802) );
  XOR U20892 ( .A(n20804), .B(n20809), .Z(n20808) );
  ANDN U20893 ( .B(n20809), .A(n20810), .Z(n20806) );
  XOR U20894 ( .A(n20811), .B(n20798), .Z(n20640) );
  NANDN U20895 ( .A(n20807), .B(n20812), .Z(n20798) );
  XOR U20896 ( .A(n20813), .B(n20801), .Z(n20812) );
  XNOR U20897 ( .A(n20814), .B(n20815), .Z(n20800) );
  XOR U20898 ( .A(n20816), .B(n20817), .Z(n20815) );
  XNOR U20899 ( .A(n20818), .B(n20819), .Z(n20814) );
  XNOR U20900 ( .A(n20820), .B(n20821), .Z(n20819) );
  ANDN U20901 ( .B(n20813), .A(n20817), .Z(n20820) );
  ANDN U20902 ( .B(n20813), .A(n20810), .Z(n20811) );
  XNOR U20903 ( .A(n20816), .B(n20822), .Z(n20810) );
  XOR U20904 ( .A(n20823), .B(n20821), .Z(n20822) );
  NAND U20905 ( .A(n20824), .B(n20825), .Z(n20821) );
  XNOR U20906 ( .A(n20818), .B(n20801), .Z(n20825) );
  IV U20907 ( .A(n20813), .Z(n20818) );
  XNOR U20908 ( .A(n20804), .B(n20817), .Z(n20824) );
  IV U20909 ( .A(n20809), .Z(n20817) );
  XOR U20910 ( .A(n20826), .B(n20827), .Z(n20809) );
  XNOR U20911 ( .A(n20828), .B(n20829), .Z(n20827) );
  XNOR U20912 ( .A(n20830), .B(n20831), .Z(n20826) );
  NOR U20913 ( .A(n20727), .B(n20639), .Z(n20830) );
  AND U20914 ( .A(n20801), .B(n20804), .Z(n20823) );
  XNOR U20915 ( .A(n20801), .B(n20804), .Z(n20816) );
  XNOR U20916 ( .A(n20832), .B(n20833), .Z(n20804) );
  XNOR U20917 ( .A(n20834), .B(n20829), .Z(n20833) );
  XOR U20918 ( .A(n20835), .B(n20836), .Z(n20832) );
  XNOR U20919 ( .A(n20837), .B(n20831), .Z(n20836) );
  OR U20920 ( .A(n20726), .B(n20790), .Z(n20831) );
  XNOR U20921 ( .A(n20639), .B(n20789), .Z(n20790) );
  XNOR U20922 ( .A(n20727), .B(n20597), .Z(n20726) );
  ANDN U20923 ( .B(n20838), .A(n20789), .Z(n20837) );
  XNOR U20924 ( .A(n20839), .B(n20840), .Z(n20801) );
  XNOR U20925 ( .A(n20829), .B(n20841), .Z(n20840) );
  XOR U20926 ( .A(n20735), .B(n20835), .Z(n20841) );
  XNOR U20927 ( .A(n20639), .B(n20842), .Z(n20829) );
  XOR U20928 ( .A(n20591), .B(n20843), .Z(n20839) );
  XNOR U20929 ( .A(n20844), .B(n20845), .Z(n20843) );
  ANDN U20930 ( .B(n20846), .A(n20794), .Z(n20844) );
  XNOR U20931 ( .A(n20847), .B(n20848), .Z(n20813) );
  XNOR U20932 ( .A(n20834), .B(n20849), .Z(n20848) );
  XNOR U20933 ( .A(n20731), .B(n20828), .Z(n20849) );
  XOR U20934 ( .A(n20835), .B(n20850), .Z(n20828) );
  XNOR U20935 ( .A(n20851), .B(n20852), .Z(n20850) );
  NAND U20936 ( .A(n20646), .B(n20741), .Z(n20852) );
  XNOR U20937 ( .A(n20853), .B(n20851), .Z(n20835) );
  NANDN U20938 ( .A(n20796), .B(n20744), .Z(n20851) );
  XOR U20939 ( .A(n20745), .B(n20741), .Z(n20744) );
  XNOR U20940 ( .A(n20846), .B(n20597), .Z(n20741) );
  XOR U20941 ( .A(n20805), .B(n20646), .Z(n20796) );
  XNOR U20942 ( .A(n20794), .B(n20854), .Z(n20646) );
  ANDN U20943 ( .B(n20745), .A(n20805), .Z(n20853) );
  XNOR U20944 ( .A(n20591), .B(n20639), .Z(n20805) );
  XOR U20945 ( .A(n20855), .B(n20856), .Z(n20639) );
  XNOR U20946 ( .A(n20857), .B(n20858), .Z(n20856) );
  XOR U20947 ( .A(n20854), .B(n20838), .Z(n20834) );
  IV U20948 ( .A(n20597), .Z(n20838) );
  XOR U20949 ( .A(n20859), .B(n20860), .Z(n20597) );
  XNOR U20950 ( .A(n20861), .B(n20858), .Z(n20860) );
  IV U20951 ( .A(n20789), .Z(n20854) );
  XOR U20952 ( .A(n20858), .B(n20862), .Z(n20789) );
  XNOR U20953 ( .A(n20863), .B(n20864), .Z(n20847) );
  XNOR U20954 ( .A(n20865), .B(n20845), .Z(n20864) );
  OR U20955 ( .A(n20737), .B(n20793), .Z(n20845) );
  XNOR U20956 ( .A(n20591), .B(n20794), .Z(n20793) );
  IV U20957 ( .A(n20863), .Z(n20794) );
  XOR U20958 ( .A(n20735), .B(n20846), .Z(n20737) );
  IV U20959 ( .A(n20731), .Z(n20846) );
  XOR U20960 ( .A(n20842), .B(n20866), .Z(n20731) );
  XNOR U20961 ( .A(n20861), .B(n20855), .Z(n20866) );
  XOR U20962 ( .A(n20867), .B(n20868), .Z(n20855) );
  XOR U20963 ( .A(n18627), .B(n19290), .Z(n20868) );
  XNOR U20964 ( .A(n20869), .B(n18640), .Z(n19290) );
  XNOR U20965 ( .A(n20870), .B(n20871), .Z(n18640) );
  XOR U20966 ( .A(n20872), .B(n20873), .Z(n20871) );
  XNOR U20967 ( .A(n20874), .B(n20875), .Z(n20870) );
  XNOR U20968 ( .A(n20876), .B(n18645), .Z(n18627) );
  XNOR U20969 ( .A(key[434]), .B(n18644), .Z(n20867) );
  IV U20970 ( .A(n20727), .Z(n20842) );
  XOR U20971 ( .A(n20859), .B(n20877), .Z(n20727) );
  XOR U20972 ( .A(n20858), .B(n20878), .Z(n20877) );
  NOR U20973 ( .A(n20735), .B(n20591), .Z(n20865) );
  XOR U20974 ( .A(n20859), .B(n20879), .Z(n20735) );
  XOR U20975 ( .A(n20858), .B(n20880), .Z(n20879) );
  XOR U20976 ( .A(n20881), .B(n20882), .Z(n20858) );
  XOR U20977 ( .A(n18615), .B(n19268), .Z(n20882) );
  XNOR U20978 ( .A(n19303), .B(n18620), .Z(n19268) );
  XNOR U20979 ( .A(n20883), .B(n20884), .Z(n18620) );
  XOR U20980 ( .A(n20885), .B(n20886), .Z(n20884) );
  XOR U20981 ( .A(n20887), .B(n20875), .Z(n20883) );
  XNOR U20982 ( .A(n18636), .B(n20888), .Z(n20881) );
  XOR U20983 ( .A(key[438]), .B(n20591), .Z(n20888) );
  XNOR U20984 ( .A(n20146), .B(n20889), .Z(n18636) );
  XNOR U20985 ( .A(n18617), .B(n19275), .Z(n20146) );
  XNOR U20986 ( .A(n20890), .B(n20891), .Z(n19275) );
  IV U20987 ( .A(n20862), .Z(n20859) );
  XOR U20988 ( .A(n20894), .B(n20895), .Z(n20862) );
  XOR U20989 ( .A(n18614), .B(n20138), .Z(n20895) );
  XOR U20990 ( .A(n18615), .B(n18634), .Z(n20138) );
  XNOR U20991 ( .A(n20896), .B(n20873), .Z(n18634) );
  XNOR U20992 ( .A(n20897), .B(n20898), .Z(n20873) );
  XOR U20993 ( .A(n20899), .B(n20900), .Z(n20898) );
  ANDN U20994 ( .B(n20901), .A(n20902), .Z(n20899) );
  XNOR U20995 ( .A(n20903), .B(n20904), .Z(n18615) );
  XNOR U20996 ( .A(n19273), .B(n20144), .Z(n18614) );
  XNOR U20997 ( .A(n20905), .B(n20906), .Z(n20144) );
  XNOR U20998 ( .A(n20907), .B(n20908), .Z(n20906) );
  XNOR U20999 ( .A(n20909), .B(n20910), .Z(n20905) );
  XOR U21000 ( .A(n20911), .B(n20912), .Z(n20910) );
  ANDN U21001 ( .B(n20913), .A(n20914), .Z(n20912) );
  XNOR U21002 ( .A(n20915), .B(n20916), .Z(n19273) );
  XOR U21003 ( .A(n20917), .B(n20918), .Z(n20916) );
  XNOR U21004 ( .A(n20919), .B(n20920), .Z(n20915) );
  XOR U21005 ( .A(n20921), .B(n20922), .Z(n20920) );
  ANDN U21006 ( .B(n20923), .A(n20924), .Z(n20922) );
  XNOR U21007 ( .A(key[437]), .B(n20145), .Z(n20894) );
  XOR U21008 ( .A(n20925), .B(n20926), .Z(n20863) );
  XNOR U21009 ( .A(n20880), .B(n20878), .Z(n20926) );
  XNOR U21010 ( .A(n20927), .B(n20928), .Z(n20878) );
  XOR U21011 ( .A(n20889), .B(n18621), .Z(n20928) );
  XNOR U21012 ( .A(n20153), .B(n19281), .Z(n18621) );
  XOR U21013 ( .A(n20929), .B(n20930), .Z(n19281) );
  XOR U21014 ( .A(n20893), .B(n20918), .Z(n20930) );
  XNOR U21015 ( .A(n20931), .B(n20932), .Z(n20918) );
  XNOR U21016 ( .A(n20933), .B(n20934), .Z(n20932) );
  NANDN U21017 ( .A(n20935), .B(n20936), .Z(n20934) );
  XNOR U21018 ( .A(n20937), .B(n20938), .Z(n20929) );
  XNOR U21019 ( .A(n20939), .B(n20940), .Z(n20153) );
  XOR U21020 ( .A(n20941), .B(n20908), .Z(n20940) );
  XNOR U21021 ( .A(n20942), .B(n20943), .Z(n20908) );
  XNOR U21022 ( .A(n20944), .B(n20945), .Z(n20943) );
  NANDN U21023 ( .A(n20946), .B(n20947), .Z(n20945) );
  XNOR U21024 ( .A(n20948), .B(n20949), .Z(n20939) );
  XNOR U21025 ( .A(n20170), .B(n20151), .Z(n20889) );
  XOR U21026 ( .A(n20950), .B(n20951), .Z(n20151) );
  XNOR U21027 ( .A(n20903), .B(n20952), .Z(n20951) );
  XNOR U21028 ( .A(key[439]), .B(n19303), .Z(n20927) );
  XNOR U21029 ( .A(n20953), .B(n20954), .Z(n20880) );
  XNOR U21030 ( .A(n18604), .B(n19284), .Z(n20954) );
  XNOR U21031 ( .A(n20955), .B(n18613), .Z(n19284) );
  XNOR U21032 ( .A(n20956), .B(n20957), .Z(n18613) );
  XOR U21033 ( .A(n20958), .B(n20886), .Z(n20957) );
  XNOR U21034 ( .A(n20959), .B(n20960), .Z(n20886) );
  XNOR U21035 ( .A(n20961), .B(n20962), .Z(n20960) );
  OR U21036 ( .A(n20963), .B(n20964), .Z(n20962) );
  XNOR U21037 ( .A(n20965), .B(n20966), .Z(n20956) );
  XNOR U21038 ( .A(n20900), .B(n20967), .Z(n20966) );
  ANDN U21039 ( .B(n20968), .A(n20969), .Z(n20967) );
  NANDN U21040 ( .A(n20970), .B(n20971), .Z(n20900) );
  XNOR U21041 ( .A(n20160), .B(n19286), .Z(n18604) );
  XOR U21042 ( .A(n20919), .B(n18645), .Z(n19286) );
  XOR U21043 ( .A(n20909), .B(n20876), .Z(n20160) );
  IV U21044 ( .A(n19294), .Z(n20876) );
  XNOR U21045 ( .A(n20973), .B(n20948), .Z(n19294) );
  XNOR U21046 ( .A(n18606), .B(n20974), .Z(n20953) );
  XOR U21047 ( .A(key[436]), .B(n20157), .Z(n20974) );
  XNOR U21048 ( .A(n20170), .B(n20145), .Z(n18606) );
  XOR U21049 ( .A(n20975), .B(n20976), .Z(n20145) );
  XNOR U21050 ( .A(n20977), .B(n20952), .Z(n20976) );
  XNOR U21051 ( .A(n20978), .B(n20979), .Z(n20952) );
  XNOR U21052 ( .A(n20980), .B(n20981), .Z(n20979) );
  OR U21053 ( .A(n20982), .B(n20983), .Z(n20981) );
  XNOR U21054 ( .A(n20984), .B(n20985), .Z(n20975) );
  XOR U21055 ( .A(n20986), .B(n20987), .Z(n20985) );
  ANDN U21056 ( .B(n20988), .A(n20989), .Z(n20987) );
  XNOR U21057 ( .A(n20591), .B(n20857), .Z(n20925) );
  XOR U21058 ( .A(n20990), .B(n20991), .Z(n20857) );
  XNOR U21059 ( .A(n19298), .B(n20992), .Z(n20991) );
  XNOR U21060 ( .A(n20861), .B(n18649), .Z(n20992) );
  XOR U21061 ( .A(n20170), .B(n20157), .Z(n18649) );
  XOR U21062 ( .A(n20977), .B(n18644), .Z(n20157) );
  IV U21063 ( .A(n20993), .Z(n18644) );
  XOR U21064 ( .A(n20994), .B(n20995), .Z(n20861) );
  XOR U21065 ( .A(n18648), .B(n19258), .Z(n20995) );
  XOR U21066 ( .A(n20993), .B(n18626), .Z(n19258) );
  XOR U21067 ( .A(n20996), .B(n20997), .Z(n20993) );
  XNOR U21068 ( .A(n20166), .B(n18654), .Z(n18648) );
  IV U21069 ( .A(n19295), .Z(n18654) );
  XOR U21070 ( .A(n20893), .B(n20998), .Z(n19295) );
  XOR U21071 ( .A(n20937), .B(n20938), .Z(n20998) );
  IV U21072 ( .A(n20999), .Z(n20938) );
  XOR U21073 ( .A(n20972), .B(n21000), .Z(n20893) );
  IV U21074 ( .A(n19302), .Z(n20166) );
  XOR U21075 ( .A(n20941), .B(n21001), .Z(n19302) );
  XOR U21076 ( .A(n20948), .B(n20949), .Z(n21001) );
  IV U21077 ( .A(n21002), .Z(n20949) );
  IV U21078 ( .A(n20891), .Z(n20941) );
  XOR U21079 ( .A(n20973), .B(n21003), .Z(n20891) );
  XNOR U21080 ( .A(key[433]), .B(n18658), .Z(n20994) );
  XOR U21081 ( .A(n19303), .B(n18608), .Z(n19298) );
  XOR U21082 ( .A(n18626), .B(n20958), .Z(n18608) );
  XOR U21083 ( .A(n20887), .B(n21004), .Z(n18626) );
  IV U21084 ( .A(n20955), .Z(n19303) );
  XOR U21085 ( .A(n21004), .B(n20958), .Z(n20955) );
  XOR U21086 ( .A(n20959), .B(n21005), .Z(n20958) );
  XOR U21087 ( .A(n21006), .B(n21007), .Z(n21005) );
  ANDN U21088 ( .B(n20901), .A(n21008), .Z(n21006) );
  XNOR U21089 ( .A(n21009), .B(n21010), .Z(n20959) );
  XNOR U21090 ( .A(n21011), .B(n21012), .Z(n21010) );
  NANDN U21091 ( .A(n21013), .B(n21014), .Z(n21012) );
  IV U21092 ( .A(n21015), .Z(n21004) );
  XNOR U21093 ( .A(n20869), .B(n21016), .Z(n20990) );
  XNOR U21094 ( .A(key[435]), .B(n20131), .Z(n21016) );
  IV U21095 ( .A(n18651), .Z(n20131) );
  XOR U21096 ( .A(n18630), .B(n19260), .Z(n18651) );
  XOR U21097 ( .A(n21017), .B(n21018), .Z(n19260) );
  XNOR U21098 ( .A(n20948), .B(n21002), .Z(n21018) );
  XOR U21099 ( .A(n21019), .B(n21020), .Z(n21002) );
  XNOR U21100 ( .A(n21021), .B(n21022), .Z(n21020) );
  NANDN U21101 ( .A(n21023), .B(n20947), .Z(n21022) );
  XNOR U21102 ( .A(n21024), .B(n21025), .Z(n20948) );
  XOR U21103 ( .A(n21026), .B(n21027), .Z(n21025) );
  NANDN U21104 ( .A(n21028), .B(n20913), .Z(n21027) );
  XNOR U21105 ( .A(n21003), .B(n20890), .Z(n21017) );
  XNOR U21106 ( .A(n21019), .B(n21029), .Z(n20890) );
  XNOR U21107 ( .A(n21030), .B(n20911), .Z(n21029) );
  ANDN U21108 ( .B(n21031), .A(n21032), .Z(n20911) );
  NOR U21109 ( .A(n21033), .B(n21034), .Z(n21030) );
  XNOR U21110 ( .A(n20907), .B(n21035), .Z(n21019) );
  XNOR U21111 ( .A(n21036), .B(n21037), .Z(n21035) );
  NAND U21112 ( .A(n21038), .B(n21039), .Z(n21037) );
  XOR U21113 ( .A(n20907), .B(n21040), .Z(n21003) );
  XNOR U21114 ( .A(n21021), .B(n21041), .Z(n21040) );
  NANDN U21115 ( .A(n21042), .B(n21043), .Z(n21041) );
  OR U21116 ( .A(n21044), .B(n21045), .Z(n21021) );
  XOR U21117 ( .A(n21046), .B(n21036), .Z(n20907) );
  NANDN U21118 ( .A(n21047), .B(n21048), .Z(n21036) );
  ANDN U21119 ( .B(n21049), .A(n21050), .Z(n21046) );
  XOR U21120 ( .A(n21051), .B(n21052), .Z(n18630) );
  XNOR U21121 ( .A(n20937), .B(n20999), .Z(n21052) );
  XNOR U21122 ( .A(n21053), .B(n21054), .Z(n20999) );
  XNOR U21123 ( .A(n21055), .B(n21056), .Z(n21054) );
  NANDN U21124 ( .A(n21057), .B(n20936), .Z(n21056) );
  XNOR U21125 ( .A(n21058), .B(n21059), .Z(n20937) );
  XOR U21126 ( .A(n21060), .B(n21061), .Z(n21059) );
  NANDN U21127 ( .A(n21062), .B(n20923), .Z(n21061) );
  XOR U21128 ( .A(n20892), .B(n21000), .Z(n21051) );
  XNOR U21129 ( .A(n20917), .B(n21063), .Z(n21000) );
  XNOR U21130 ( .A(n21055), .B(n21064), .Z(n21063) );
  NANDN U21131 ( .A(n21065), .B(n21066), .Z(n21064) );
  OR U21132 ( .A(n21067), .B(n21068), .Z(n21055) );
  XNOR U21133 ( .A(n21053), .B(n21069), .Z(n20892) );
  XNOR U21134 ( .A(n21070), .B(n20921), .Z(n21069) );
  ANDN U21135 ( .B(n21071), .A(n21072), .Z(n20921) );
  NOR U21136 ( .A(n21073), .B(n21074), .Z(n21070) );
  XNOR U21137 ( .A(n20917), .B(n21075), .Z(n21053) );
  XNOR U21138 ( .A(n21076), .B(n21077), .Z(n21075) );
  NAND U21139 ( .A(n21078), .B(n21079), .Z(n21077) );
  XNOR U21140 ( .A(n21080), .B(n21076), .Z(n20917) );
  NANDN U21141 ( .A(n21081), .B(n21082), .Z(n21076) );
  ANDN U21142 ( .B(n21083), .A(n21084), .Z(n21080) );
  IV U21143 ( .A(n18628), .Z(n20869) );
  XNOR U21144 ( .A(n20950), .B(n21085), .Z(n18628) );
  XOR U21145 ( .A(n21086), .B(n20904), .Z(n21085) );
  XNOR U21146 ( .A(n21087), .B(n21088), .Z(n20904) );
  XNOR U21147 ( .A(n21089), .B(n20986), .Z(n21088) );
  ANDN U21148 ( .B(n21090), .A(n21091), .Z(n20986) );
  ANDN U21149 ( .B(n21092), .A(n21093), .Z(n21089) );
  XNOR U21150 ( .A(n20996), .B(n21094), .Z(n20950) );
  XNOR U21151 ( .A(n21095), .B(n21096), .Z(n20591) );
  XOR U21152 ( .A(n19297), .B(n18622), .Z(n21096) );
  IV U21153 ( .A(n19304), .Z(n18622) );
  XOR U21154 ( .A(n18656), .B(n20170), .Z(n19304) );
  XOR U21155 ( .A(n21097), .B(n20977), .Z(n20170) );
  XNOR U21156 ( .A(n20978), .B(n21098), .Z(n20977) );
  XOR U21157 ( .A(n21099), .B(n21100), .Z(n21098) );
  ANDN U21158 ( .B(n21092), .A(n21101), .Z(n21099) );
  XNOR U21159 ( .A(n21102), .B(n21103), .Z(n20978) );
  XNOR U21160 ( .A(n21104), .B(n21105), .Z(n21103) );
  NANDN U21161 ( .A(n21106), .B(n21107), .Z(n21105) );
  IV U21162 ( .A(n20140), .Z(n18656) );
  XOR U21163 ( .A(n20919), .B(n20972), .Z(n20140) );
  XOR U21164 ( .A(n21109), .B(n20933), .Z(n21108) );
  OR U21165 ( .A(n21110), .B(n21067), .Z(n20933) );
  XNOR U21166 ( .A(n20936), .B(n21066), .Z(n21067) );
  ANDN U21167 ( .B(n21066), .A(n21111), .Z(n21109) );
  XNOR U21168 ( .A(n20931), .B(n21112), .Z(n20919) );
  XNOR U21169 ( .A(n21113), .B(n21060), .Z(n21112) );
  XNOR U21170 ( .A(n21074), .B(n20923), .Z(n21071) );
  ANDN U21171 ( .B(n21115), .A(n21074), .Z(n21113) );
  XOR U21172 ( .A(n21058), .B(n21116), .Z(n20931) );
  XNOR U21173 ( .A(n21117), .B(n21118), .Z(n21116) );
  NAND U21174 ( .A(n21079), .B(n21119), .Z(n21118) );
  XNOR U21175 ( .A(n21120), .B(n21117), .Z(n21058) );
  OR U21176 ( .A(n21081), .B(n21121), .Z(n21117) );
  XNOR U21177 ( .A(n21122), .B(n21079), .Z(n21081) );
  XOR U21178 ( .A(n21066), .B(n20923), .Z(n21079) );
  XOR U21179 ( .A(n21123), .B(n21124), .Z(n20923) );
  NANDN U21180 ( .A(n21125), .B(n21126), .Z(n21124) );
  XOR U21181 ( .A(n21127), .B(n21128), .Z(n21066) );
  NANDN U21182 ( .A(n21125), .B(n21129), .Z(n21128) );
  ANDN U21183 ( .B(n21122), .A(n21130), .Z(n21120) );
  IV U21184 ( .A(n21084), .Z(n21122) );
  XOR U21185 ( .A(n21074), .B(n20936), .Z(n21084) );
  XNOR U21186 ( .A(n21131), .B(n21127), .Z(n20936) );
  NANDN U21187 ( .A(n21132), .B(n21133), .Z(n21127) );
  XOR U21188 ( .A(n21129), .B(n21134), .Z(n21133) );
  ANDN U21189 ( .B(n21134), .A(n21135), .Z(n21131) );
  XOR U21190 ( .A(n21136), .B(n21123), .Z(n21074) );
  NANDN U21191 ( .A(n21132), .B(n21137), .Z(n21123) );
  XOR U21192 ( .A(n21138), .B(n21126), .Z(n21137) );
  XNOR U21193 ( .A(n21139), .B(n21140), .Z(n21125) );
  XOR U21194 ( .A(n21141), .B(n21142), .Z(n21140) );
  XNOR U21195 ( .A(n21143), .B(n21144), .Z(n21139) );
  XNOR U21196 ( .A(n21145), .B(n21146), .Z(n21144) );
  ANDN U21197 ( .B(n21138), .A(n21142), .Z(n21145) );
  ANDN U21198 ( .B(n21138), .A(n21135), .Z(n21136) );
  XNOR U21199 ( .A(n21141), .B(n21147), .Z(n21135) );
  XOR U21200 ( .A(n21148), .B(n21146), .Z(n21147) );
  NAND U21201 ( .A(n21149), .B(n21150), .Z(n21146) );
  XNOR U21202 ( .A(n21143), .B(n21126), .Z(n21150) );
  IV U21203 ( .A(n21138), .Z(n21143) );
  XNOR U21204 ( .A(n21129), .B(n21142), .Z(n21149) );
  IV U21205 ( .A(n21134), .Z(n21142) );
  XOR U21206 ( .A(n21151), .B(n21152), .Z(n21134) );
  XNOR U21207 ( .A(n21153), .B(n21154), .Z(n21152) );
  XNOR U21208 ( .A(n21155), .B(n21156), .Z(n21151) );
  ANDN U21209 ( .B(n21115), .A(n21073), .Z(n21155) );
  AND U21210 ( .A(n21126), .B(n21129), .Z(n21148) );
  XNOR U21211 ( .A(n21126), .B(n21129), .Z(n21141) );
  XNOR U21212 ( .A(n21157), .B(n21158), .Z(n21129) );
  XNOR U21213 ( .A(n21159), .B(n21154), .Z(n21158) );
  XOR U21214 ( .A(n21160), .B(n21161), .Z(n21157) );
  XNOR U21215 ( .A(n21162), .B(n21156), .Z(n21161) );
  OR U21216 ( .A(n21072), .B(n21114), .Z(n21156) );
  XNOR U21217 ( .A(n21115), .B(n21163), .Z(n21114) );
  XNOR U21218 ( .A(n21073), .B(n20924), .Z(n21072) );
  ANDN U21219 ( .B(n21164), .A(n21062), .Z(n21162) );
  XNOR U21220 ( .A(n21165), .B(n21166), .Z(n21126) );
  XNOR U21221 ( .A(n21154), .B(n21167), .Z(n21166) );
  XOR U21222 ( .A(n21057), .B(n21160), .Z(n21167) );
  XNOR U21223 ( .A(n21115), .B(n21073), .Z(n21154) );
  XOR U21224 ( .A(n20935), .B(n21168), .Z(n21165) );
  XNOR U21225 ( .A(n21169), .B(n21170), .Z(n21168) );
  ANDN U21226 ( .B(n21171), .A(n21111), .Z(n21169) );
  XNOR U21227 ( .A(n21172), .B(n21173), .Z(n21138) );
  XNOR U21228 ( .A(n21159), .B(n21174), .Z(n21173) );
  XNOR U21229 ( .A(n21065), .B(n21153), .Z(n21174) );
  XOR U21230 ( .A(n21160), .B(n21175), .Z(n21153) );
  XNOR U21231 ( .A(n21176), .B(n21177), .Z(n21175) );
  NAND U21232 ( .A(n21119), .B(n21078), .Z(n21177) );
  XNOR U21233 ( .A(n21178), .B(n21176), .Z(n21160) );
  NANDN U21234 ( .A(n21121), .B(n21082), .Z(n21176) );
  XOR U21235 ( .A(n21083), .B(n21078), .Z(n21082) );
  XNOR U21236 ( .A(n21171), .B(n20924), .Z(n21078) );
  XOR U21237 ( .A(n21130), .B(n21119), .Z(n21121) );
  XNOR U21238 ( .A(n21111), .B(n21163), .Z(n21119) );
  ANDN U21239 ( .B(n21083), .A(n21130), .Z(n21178) );
  XOR U21240 ( .A(n20935), .B(n21115), .Z(n21130) );
  XNOR U21241 ( .A(n21179), .B(n21180), .Z(n21115) );
  XNOR U21242 ( .A(n21181), .B(n21182), .Z(n21180) );
  XOR U21243 ( .A(n21163), .B(n21164), .Z(n21159) );
  IV U21244 ( .A(n20924), .Z(n21164) );
  XOR U21245 ( .A(n21183), .B(n21184), .Z(n20924) );
  XOR U21246 ( .A(n21185), .B(n21182), .Z(n21184) );
  IV U21247 ( .A(n21062), .Z(n21163) );
  XOR U21248 ( .A(n21182), .B(n21186), .Z(n21062) );
  XNOR U21249 ( .A(n21187), .B(n21188), .Z(n21172) );
  XNOR U21250 ( .A(n21189), .B(n21170), .Z(n21188) );
  OR U21251 ( .A(n21068), .B(n21110), .Z(n21170) );
  XNOR U21252 ( .A(n20935), .B(n21111), .Z(n21110) );
  IV U21253 ( .A(n21187), .Z(n21111) );
  XOR U21254 ( .A(n21057), .B(n21171), .Z(n21068) );
  IV U21255 ( .A(n21065), .Z(n21171) );
  XNOR U21256 ( .A(n21191), .B(n21179), .Z(n21190) );
  XOR U21257 ( .A(n21192), .B(n21193), .Z(n21179) );
  XOR U21258 ( .A(n21194), .B(n21195), .Z(n21193) );
  XNOR U21259 ( .A(key[322]), .B(n21196), .Z(n21192) );
  XOR U21260 ( .A(n21183), .B(n21197), .Z(n21073) );
  XOR U21261 ( .A(n21182), .B(n21198), .Z(n21197) );
  NOR U21262 ( .A(n21057), .B(n20935), .Z(n21189) );
  XOR U21263 ( .A(n21183), .B(n21199), .Z(n21057) );
  XOR U21264 ( .A(n21182), .B(n21200), .Z(n21199) );
  XOR U21265 ( .A(n21201), .B(n21202), .Z(n21182) );
  XNOR U21266 ( .A(n20935), .B(n21203), .Z(n21202) );
  XNOR U21267 ( .A(n21204), .B(n21205), .Z(n21201) );
  XNOR U21268 ( .A(key[326]), .B(n21206), .Z(n21205) );
  IV U21269 ( .A(n21186), .Z(n21183) );
  XOR U21270 ( .A(n21207), .B(n21208), .Z(n21186) );
  XNOR U21271 ( .A(n21209), .B(n21210), .Z(n21208) );
  XNOR U21272 ( .A(key[325]), .B(n21211), .Z(n21207) );
  XOR U21273 ( .A(n21212), .B(n21213), .Z(n21187) );
  XNOR U21274 ( .A(n21200), .B(n21198), .Z(n21213) );
  XNOR U21275 ( .A(n21214), .B(n21215), .Z(n21198) );
  XOR U21276 ( .A(n21216), .B(n21217), .Z(n21215) );
  XNOR U21277 ( .A(key[327]), .B(n21218), .Z(n21214) );
  XNOR U21278 ( .A(n21219), .B(n21220), .Z(n21200) );
  XOR U21279 ( .A(n21221), .B(n21222), .Z(n21220) );
  XNOR U21280 ( .A(n21223), .B(n21224), .Z(n21219) );
  XNOR U21281 ( .A(key[324]), .B(n21225), .Z(n21224) );
  XNOR U21282 ( .A(n20935), .B(n21181), .Z(n21212) );
  XOR U21283 ( .A(n21226), .B(n21227), .Z(n21181) );
  XNOR U21284 ( .A(n21228), .B(n21229), .Z(n21227) );
  XOR U21285 ( .A(n21230), .B(n21191), .Z(n21229) );
  IV U21286 ( .A(n21185), .Z(n21191) );
  XNOR U21287 ( .A(n21231), .B(n21232), .Z(n21185) );
  XOR U21288 ( .A(n21233), .B(n21234), .Z(n21232) );
  XOR U21289 ( .A(key[321]), .B(n21235), .Z(n21231) );
  XNOR U21290 ( .A(n21236), .B(n21237), .Z(n21226) );
  XNOR U21291 ( .A(key[323]), .B(n21238), .Z(n21237) );
  XNOR U21292 ( .A(n21239), .B(n21240), .Z(n20935) );
  XOR U21293 ( .A(key[320]), .B(n21243), .Z(n21239) );
  XOR U21294 ( .A(n18647), .B(n18658), .Z(n19297) );
  XNOR U21295 ( .A(n20903), .B(n21244), .Z(n18658) );
  XOR U21296 ( .A(n20996), .B(n21094), .Z(n21244) );
  XOR U21297 ( .A(n21087), .B(n21245), .Z(n21094) );
  XNOR U21298 ( .A(n21246), .B(n21247), .Z(n21245) );
  OR U21299 ( .A(n20982), .B(n21248), .Z(n21247) );
  XNOR U21300 ( .A(n20984), .B(n21249), .Z(n21087) );
  XNOR U21301 ( .A(n21250), .B(n21251), .Z(n21249) );
  NANDN U21302 ( .A(n21106), .B(n21252), .Z(n21251) );
  XNOR U21303 ( .A(n21102), .B(n21253), .Z(n20996) );
  XNOR U21304 ( .A(n21100), .B(n21254), .Z(n21253) );
  NAND U21305 ( .A(n21255), .B(n20988), .Z(n21254) );
  XOR U21306 ( .A(n21092), .B(n20988), .Z(n21090) );
  XNOR U21307 ( .A(n21097), .B(n21086), .Z(n20903) );
  XOR U21308 ( .A(n20984), .B(n21257), .Z(n21086) );
  XNOR U21309 ( .A(n21246), .B(n21258), .Z(n21257) );
  NANDN U21310 ( .A(n21259), .B(n21260), .Z(n21258) );
  OR U21311 ( .A(n21261), .B(n21262), .Z(n21246) );
  XOR U21312 ( .A(n21263), .B(n21250), .Z(n20984) );
  NANDN U21313 ( .A(n21264), .B(n21265), .Z(n21250) );
  ANDN U21314 ( .B(n21266), .A(n21267), .Z(n21263) );
  IV U21315 ( .A(n20997), .Z(n21097) );
  XNOR U21316 ( .A(n21102), .B(n21268), .Z(n20997) );
  XOR U21317 ( .A(n21269), .B(n20980), .Z(n21268) );
  OR U21318 ( .A(n21270), .B(n21261), .Z(n20980) );
  XNOR U21319 ( .A(n20982), .B(n21259), .Z(n21261) );
  NOR U21320 ( .A(n21271), .B(n21259), .Z(n21269) );
  XOR U21321 ( .A(n21272), .B(n21104), .Z(n21102) );
  OR U21322 ( .A(n21264), .B(n21273), .Z(n21104) );
  XOR U21323 ( .A(n21274), .B(n21106), .Z(n21264) );
  XOR U21324 ( .A(n21259), .B(n20988), .Z(n21106) );
  XOR U21325 ( .A(n21275), .B(n21276), .Z(n20988) );
  NANDN U21326 ( .A(n21277), .B(n21278), .Z(n21276) );
  XNOR U21327 ( .A(n21279), .B(n21280), .Z(n21259) );
  OR U21328 ( .A(n21277), .B(n21281), .Z(n21280) );
  ANDN U21329 ( .B(n21274), .A(n21282), .Z(n21272) );
  IV U21330 ( .A(n21267), .Z(n21274) );
  XOR U21331 ( .A(n20982), .B(n21092), .Z(n21267) );
  XNOR U21332 ( .A(n21283), .B(n21275), .Z(n21092) );
  NANDN U21333 ( .A(n21284), .B(n21285), .Z(n21275) );
  ANDN U21334 ( .B(n21286), .A(n21287), .Z(n21283) );
  NANDN U21335 ( .A(n21284), .B(n21289), .Z(n21279) );
  XOR U21336 ( .A(n21290), .B(n21277), .Z(n21284) );
  XNOR U21337 ( .A(n21291), .B(n21292), .Z(n21277) );
  XOR U21338 ( .A(n21293), .B(n21286), .Z(n21292) );
  XNOR U21339 ( .A(n21294), .B(n21295), .Z(n21291) );
  XNOR U21340 ( .A(n21296), .B(n21297), .Z(n21295) );
  ANDN U21341 ( .B(n21286), .A(n21298), .Z(n21296) );
  IV U21342 ( .A(n21299), .Z(n21286) );
  ANDN U21343 ( .B(n21290), .A(n21298), .Z(n21288) );
  IV U21344 ( .A(n21294), .Z(n21298) );
  IV U21345 ( .A(n21287), .Z(n21290) );
  XNOR U21346 ( .A(n21293), .B(n21300), .Z(n21287) );
  XOR U21347 ( .A(n21301), .B(n21297), .Z(n21300) );
  NAND U21348 ( .A(n21289), .B(n21285), .Z(n21297) );
  XNOR U21349 ( .A(n21278), .B(n21299), .Z(n21285) );
  XOR U21350 ( .A(n21302), .B(n21303), .Z(n21299) );
  XOR U21351 ( .A(n21304), .B(n21305), .Z(n21303) );
  XNOR U21352 ( .A(n21260), .B(n21306), .Z(n21305) );
  XNOR U21353 ( .A(n21307), .B(n21308), .Z(n21302) );
  XNOR U21354 ( .A(n21309), .B(n21310), .Z(n21308) );
  ANDN U21355 ( .B(n21311), .A(n20983), .Z(n21309) );
  XNOR U21356 ( .A(n21294), .B(n21281), .Z(n21289) );
  XOR U21357 ( .A(n21312), .B(n21313), .Z(n21294) );
  XNOR U21358 ( .A(n21314), .B(n21306), .Z(n21313) );
  XOR U21359 ( .A(n21315), .B(n21316), .Z(n21306) );
  XNOR U21360 ( .A(n21317), .B(n21318), .Z(n21316) );
  NAND U21361 ( .A(n21107), .B(n21252), .Z(n21318) );
  XNOR U21362 ( .A(n21319), .B(n21320), .Z(n21312) );
  ANDN U21363 ( .B(n21321), .A(n21101), .Z(n21319) );
  ANDN U21364 ( .B(n21278), .A(n21281), .Z(n21301) );
  XOR U21365 ( .A(n21281), .B(n21278), .Z(n21293) );
  XNOR U21366 ( .A(n21322), .B(n21323), .Z(n21278) );
  XNOR U21367 ( .A(n21315), .B(n21324), .Z(n21323) );
  XOR U21368 ( .A(n21314), .B(n21248), .Z(n21324) );
  XOR U21369 ( .A(n20983), .B(n21325), .Z(n21322) );
  XNOR U21370 ( .A(n21326), .B(n21310), .Z(n21325) );
  OR U21371 ( .A(n21262), .B(n21270), .Z(n21310) );
  XNOR U21372 ( .A(n20983), .B(n21271), .Z(n21270) );
  XOR U21373 ( .A(n21248), .B(n21260), .Z(n21262) );
  ANDN U21374 ( .B(n21260), .A(n21271), .Z(n21326) );
  XOR U21375 ( .A(n21327), .B(n21328), .Z(n21281) );
  XOR U21376 ( .A(n21315), .B(n21304), .Z(n21328) );
  XOR U21377 ( .A(n21255), .B(n20989), .Z(n21304) );
  XOR U21378 ( .A(n21329), .B(n21317), .Z(n21315) );
  NANDN U21379 ( .A(n21273), .B(n21265), .Z(n21317) );
  XOR U21380 ( .A(n21266), .B(n21252), .Z(n21265) );
  XNOR U21381 ( .A(n21321), .B(n21330), .Z(n21260) );
  XOR U21382 ( .A(n21331), .B(n21332), .Z(n21330) );
  XOR U21383 ( .A(n21282), .B(n21107), .Z(n21273) );
  XNOR U21384 ( .A(n21271), .B(n21255), .Z(n21107) );
  IV U21385 ( .A(n21307), .Z(n21271) );
  XOR U21386 ( .A(n21333), .B(n21334), .Z(n21307) );
  XOR U21387 ( .A(n21335), .B(n21336), .Z(n21334) );
  XNOR U21388 ( .A(n20983), .B(n21337), .Z(n21333) );
  ANDN U21389 ( .B(n21266), .A(n21282), .Z(n21329) );
  XNOR U21390 ( .A(n20983), .B(n21101), .Z(n21282) );
  XOR U21391 ( .A(n21321), .B(n21311), .Z(n21266) );
  IV U21392 ( .A(n21248), .Z(n21311) );
  XOR U21393 ( .A(n21338), .B(n21339), .Z(n21248) );
  XOR U21394 ( .A(n21340), .B(n21336), .Z(n21339) );
  XNOR U21395 ( .A(n21341), .B(n21342), .Z(n21336) );
  XNOR U21396 ( .A(n21343), .B(n21344), .Z(n21342) );
  XNOR U21397 ( .A(n21345), .B(n21346), .Z(n21341) );
  XNOR U21398 ( .A(key[364]), .B(n21347), .Z(n21346) );
  IV U21399 ( .A(n21093), .Z(n21321) );
  XOR U21400 ( .A(n21314), .B(n21348), .Z(n21327) );
  XNOR U21401 ( .A(n21349), .B(n21320), .Z(n21348) );
  OR U21402 ( .A(n21091), .B(n21256), .Z(n21320) );
  XNOR U21403 ( .A(n21350), .B(n21255), .Z(n21256) );
  XNOR U21404 ( .A(n21093), .B(n20989), .Z(n21091) );
  ANDN U21405 ( .B(n21255), .A(n20989), .Z(n21349) );
  XOR U21406 ( .A(n21338), .B(n21351), .Z(n20989) );
  XNOR U21407 ( .A(n21352), .B(n21340), .Z(n21351) );
  XOR U21408 ( .A(n21340), .B(n21338), .Z(n21255) );
  XNOR U21409 ( .A(n21101), .B(n21093), .Z(n21314) );
  XOR U21410 ( .A(n21338), .B(n21353), .Z(n21093) );
  XNOR U21411 ( .A(n21340), .B(n21335), .Z(n21353) );
  XOR U21412 ( .A(n21354), .B(n21355), .Z(n21335) );
  XOR U21413 ( .A(n21356), .B(n21357), .Z(n21355) );
  XNOR U21414 ( .A(key[367]), .B(n21358), .Z(n21354) );
  XNOR U21415 ( .A(n21359), .B(n21360), .Z(n21338) );
  XNOR U21416 ( .A(n21361), .B(n21362), .Z(n21360) );
  XOR U21417 ( .A(n21363), .B(n21364), .Z(n21359) );
  XOR U21418 ( .A(key[365]), .B(n21365), .Z(n21364) );
  IV U21419 ( .A(n21350), .Z(n21101) );
  XNOR U21420 ( .A(n21332), .B(n21366), .Z(n21350) );
  XOR U21421 ( .A(n21367), .B(n21368), .Z(n21340) );
  XOR U21422 ( .A(n20983), .B(n21369), .Z(n21368) );
  XNOR U21423 ( .A(n21370), .B(n21371), .Z(n20983) );
  XOR U21424 ( .A(n21372), .B(n21373), .Z(n21371) );
  XNOR U21425 ( .A(n21374), .B(n21375), .Z(n21370) );
  XOR U21426 ( .A(key[360]), .B(n21376), .Z(n21375) );
  XOR U21427 ( .A(n21377), .B(n21378), .Z(n21367) );
  XNOR U21428 ( .A(key[366]), .B(n21379), .Z(n21378) );
  XOR U21429 ( .A(n21380), .B(n21381), .Z(n21337) );
  XNOR U21430 ( .A(n21382), .B(n21383), .Z(n21381) );
  XNOR U21431 ( .A(n21384), .B(n21352), .Z(n21383) );
  IV U21432 ( .A(n21331), .Z(n21352) );
  XNOR U21433 ( .A(n21385), .B(n21386), .Z(n21331) );
  XOR U21434 ( .A(n21387), .B(n21388), .Z(n21386) );
  XNOR U21435 ( .A(n21389), .B(n21390), .Z(n21385) );
  XOR U21436 ( .A(key[361]), .B(n21391), .Z(n21390) );
  XNOR U21437 ( .A(n21392), .B(n21393), .Z(n21380) );
  XNOR U21438 ( .A(key[363]), .B(n21394), .Z(n21393) );
  XOR U21439 ( .A(n21395), .B(n21396), .Z(n21332) );
  XOR U21440 ( .A(n21397), .B(n21398), .Z(n21396) );
  XOR U21441 ( .A(n21399), .B(n21400), .Z(n21395) );
  XNOR U21442 ( .A(key[362]), .B(n21401), .Z(n21400) );
  IV U21443 ( .A(n19306), .Z(n18647) );
  XOR U21444 ( .A(n20885), .B(n21402), .Z(n19306) );
  XOR U21445 ( .A(n20874), .B(n20875), .Z(n21402) );
  XOR U21446 ( .A(n20897), .B(n21403), .Z(n20875) );
  XNOR U21447 ( .A(n21404), .B(n21405), .Z(n21403) );
  OR U21448 ( .A(n20963), .B(n21406), .Z(n21405) );
  XNOR U21449 ( .A(n20965), .B(n21407), .Z(n20897) );
  XNOR U21450 ( .A(n21408), .B(n21409), .Z(n21407) );
  NANDN U21451 ( .A(n21013), .B(n21410), .Z(n21409) );
  IV U21452 ( .A(n20887), .Z(n20874) );
  XOR U21453 ( .A(n21009), .B(n21411), .Z(n20887) );
  XNOR U21454 ( .A(n21007), .B(n21412), .Z(n21411) );
  NAND U21455 ( .A(n21413), .B(n20968), .Z(n21412) );
  NANDN U21456 ( .A(n21414), .B(n20971), .Z(n21007) );
  XOR U21457 ( .A(n20901), .B(n20968), .Z(n20971) );
  IV U21458 ( .A(n20896), .Z(n20885) );
  XOR U21459 ( .A(n20872), .B(n21015), .Z(n20896) );
  XNOR U21460 ( .A(n21009), .B(n21415), .Z(n21015) );
  XOR U21461 ( .A(n21416), .B(n20961), .Z(n21415) );
  OR U21462 ( .A(n21417), .B(n21418), .Z(n20961) );
  NOR U21463 ( .A(n21419), .B(n21420), .Z(n21416) );
  XOR U21464 ( .A(n21421), .B(n21011), .Z(n21009) );
  OR U21465 ( .A(n21422), .B(n21423), .Z(n21011) );
  ANDN U21466 ( .B(n21424), .A(n21425), .Z(n21421) );
  XOR U21467 ( .A(n20965), .B(n21426), .Z(n20872) );
  XNOR U21468 ( .A(n21404), .B(n21427), .Z(n21426) );
  NANDN U21469 ( .A(n21420), .B(n21428), .Z(n21427) );
  OR U21470 ( .A(n21417), .B(n21429), .Z(n21404) );
  XNOR U21471 ( .A(n20963), .B(n21420), .Z(n21417) );
  XOR U21472 ( .A(n21430), .B(n21408), .Z(n20965) );
  NANDN U21473 ( .A(n21422), .B(n21431), .Z(n21408) );
  XOR U21474 ( .A(n21424), .B(n21013), .Z(n21422) );
  XOR U21475 ( .A(n21420), .B(n20968), .Z(n21013) );
  XOR U21476 ( .A(n21432), .B(n21433), .Z(n20968) );
  NANDN U21477 ( .A(n21434), .B(n21435), .Z(n21433) );
  XNOR U21478 ( .A(n21436), .B(n21437), .Z(n21420) );
  OR U21479 ( .A(n21434), .B(n21438), .Z(n21437) );
  IV U21480 ( .A(n21439), .Z(n21424) );
  ANDN U21481 ( .B(n21440), .A(n21439), .Z(n21430) );
  XOR U21482 ( .A(n20963), .B(n20901), .Z(n21439) );
  XNOR U21483 ( .A(n21441), .B(n21432), .Z(n20901) );
  NANDN U21484 ( .A(n21442), .B(n21443), .Z(n21432) );
  ANDN U21485 ( .B(n21444), .A(n21445), .Z(n21441) );
  NANDN U21486 ( .A(n21442), .B(n21447), .Z(n21436) );
  XOR U21487 ( .A(n21448), .B(n21434), .Z(n21442) );
  XNOR U21488 ( .A(n21449), .B(n21450), .Z(n21434) );
  XOR U21489 ( .A(n21451), .B(n21444), .Z(n21450) );
  XNOR U21490 ( .A(n21452), .B(n21453), .Z(n21449) );
  XNOR U21491 ( .A(n21454), .B(n21455), .Z(n21453) );
  ANDN U21492 ( .B(n21444), .A(n21456), .Z(n21454) );
  IV U21493 ( .A(n21457), .Z(n21444) );
  ANDN U21494 ( .B(n21448), .A(n21456), .Z(n21446) );
  IV U21495 ( .A(n21452), .Z(n21456) );
  IV U21496 ( .A(n21445), .Z(n21448) );
  XNOR U21497 ( .A(n21451), .B(n21458), .Z(n21445) );
  XOR U21498 ( .A(n21459), .B(n21455), .Z(n21458) );
  NAND U21499 ( .A(n21447), .B(n21443), .Z(n21455) );
  XNOR U21500 ( .A(n21435), .B(n21457), .Z(n21443) );
  XOR U21501 ( .A(n21460), .B(n21461), .Z(n21457) );
  XOR U21502 ( .A(n21462), .B(n21463), .Z(n21461) );
  XNOR U21503 ( .A(n21428), .B(n21464), .Z(n21463) );
  XNOR U21504 ( .A(n21465), .B(n21466), .Z(n21460) );
  XNOR U21505 ( .A(n21467), .B(n21468), .Z(n21466) );
  ANDN U21506 ( .B(n21469), .A(n20964), .Z(n21467) );
  XNOR U21507 ( .A(n21452), .B(n21438), .Z(n21447) );
  XOR U21508 ( .A(n21470), .B(n21471), .Z(n21452) );
  XNOR U21509 ( .A(n21472), .B(n21464), .Z(n21471) );
  XOR U21510 ( .A(n21473), .B(n21474), .Z(n21464) );
  XNOR U21511 ( .A(n21475), .B(n21476), .Z(n21474) );
  NAND U21512 ( .A(n21014), .B(n21410), .Z(n21476) );
  XNOR U21513 ( .A(n21477), .B(n21478), .Z(n21470) );
  ANDN U21514 ( .B(n21479), .A(n21008), .Z(n21477) );
  ANDN U21515 ( .B(n21435), .A(n21438), .Z(n21459) );
  XOR U21516 ( .A(n21438), .B(n21435), .Z(n21451) );
  XNOR U21517 ( .A(n21480), .B(n21481), .Z(n21435) );
  XNOR U21518 ( .A(n21473), .B(n21482), .Z(n21481) );
  XOR U21519 ( .A(n21472), .B(n21406), .Z(n21482) );
  XOR U21520 ( .A(n20964), .B(n21483), .Z(n21480) );
  XNOR U21521 ( .A(n21484), .B(n21468), .Z(n21483) );
  OR U21522 ( .A(n21429), .B(n21418), .Z(n21468) );
  XNOR U21523 ( .A(n20964), .B(n21419), .Z(n21418) );
  XOR U21524 ( .A(n21406), .B(n21428), .Z(n21429) );
  ANDN U21525 ( .B(n21428), .A(n21419), .Z(n21484) );
  XOR U21526 ( .A(n21485), .B(n21486), .Z(n21438) );
  XOR U21527 ( .A(n21473), .B(n21462), .Z(n21486) );
  XOR U21528 ( .A(n21413), .B(n20969), .Z(n21462) );
  XOR U21529 ( .A(n21487), .B(n21475), .Z(n21473) );
  NANDN U21530 ( .A(n21423), .B(n21431), .Z(n21475) );
  XOR U21531 ( .A(n21440), .B(n21410), .Z(n21431) );
  XNOR U21532 ( .A(n21479), .B(n21488), .Z(n21428) );
  XOR U21533 ( .A(n21489), .B(n21490), .Z(n21488) );
  XOR U21534 ( .A(n21425), .B(n21014), .Z(n21423) );
  XNOR U21535 ( .A(n21419), .B(n21413), .Z(n21014) );
  IV U21536 ( .A(n21465), .Z(n21419) );
  XOR U21537 ( .A(n21491), .B(n21492), .Z(n21465) );
  XOR U21538 ( .A(n21493), .B(n21494), .Z(n21492) );
  XNOR U21539 ( .A(n20964), .B(n21495), .Z(n21491) );
  ANDN U21540 ( .B(n21440), .A(n21425), .Z(n21487) );
  XNOR U21541 ( .A(n20964), .B(n21008), .Z(n21425) );
  XOR U21542 ( .A(n21472), .B(n21496), .Z(n21485) );
  XNOR U21543 ( .A(n21497), .B(n21478), .Z(n21496) );
  OR U21544 ( .A(n20970), .B(n21414), .Z(n21478) );
  XNOR U21545 ( .A(n21498), .B(n21413), .Z(n21414) );
  XNOR U21546 ( .A(n20902), .B(n20969), .Z(n20970) );
  ANDN U21547 ( .B(n21413), .A(n20969), .Z(n21497) );
  XOR U21548 ( .A(n21499), .B(n21500), .Z(n20969) );
  XNOR U21549 ( .A(n21501), .B(n21502), .Z(n21500) );
  XOR U21550 ( .A(n21502), .B(n21499), .Z(n21413) );
  XNOR U21551 ( .A(n21008), .B(n20902), .Z(n21472) );
  IV U21552 ( .A(n21498), .Z(n21008) );
  XNOR U21553 ( .A(n21490), .B(n21503), .Z(n21498) );
  XOR U21554 ( .A(n21504), .B(n21505), .Z(n21495) );
  XNOR U21555 ( .A(n21506), .B(n21507), .Z(n21505) );
  XOR U21556 ( .A(n21508), .B(n21501), .Z(n21507) );
  IV U21557 ( .A(n21489), .Z(n21501) );
  XNOR U21558 ( .A(n21509), .B(n21510), .Z(n21489) );
  XOR U21559 ( .A(n21511), .B(n21512), .Z(n21510) );
  XOR U21560 ( .A(key[273]), .B(n21513), .Z(n21509) );
  XNOR U21561 ( .A(n21514), .B(n21515), .Z(n21504) );
  XNOR U21562 ( .A(key[275]), .B(n21516), .Z(n21515) );
  XOR U21563 ( .A(n21517), .B(n21518), .Z(n21490) );
  XOR U21564 ( .A(n21519), .B(n21520), .Z(n21518) );
  XNOR U21565 ( .A(key[274]), .B(n21521), .Z(n21517) );
  XOR U21566 ( .A(n21479), .B(n21469), .Z(n21440) );
  IV U21567 ( .A(n21406), .Z(n21469) );
  XOR U21568 ( .A(n21499), .B(n21522), .Z(n21406) );
  XOR U21569 ( .A(n21502), .B(n21494), .Z(n21522) );
  XNOR U21570 ( .A(n21523), .B(n21524), .Z(n21494) );
  XOR U21571 ( .A(n21525), .B(n21526), .Z(n21524) );
  IV U21572 ( .A(n20902), .Z(n21479) );
  XOR U21573 ( .A(n21499), .B(n21528), .Z(n20902) );
  XNOR U21574 ( .A(n21502), .B(n21493), .Z(n21528) );
  XOR U21575 ( .A(n21529), .B(n21530), .Z(n21493) );
  XOR U21576 ( .A(n21531), .B(n21532), .Z(n21530) );
  XNOR U21577 ( .A(key[279]), .B(n21533), .Z(n21529) );
  XOR U21578 ( .A(n21534), .B(n21535), .Z(n21502) );
  XNOR U21579 ( .A(n20964), .B(n21536), .Z(n21535) );
  XNOR U21580 ( .A(n21537), .B(n21538), .Z(n20964) );
  XNOR U21581 ( .A(n21539), .B(n21540), .Z(n21538) );
  XNOR U21582 ( .A(n21542), .B(n21543), .Z(n21534) );
  XOR U21583 ( .A(key[278]), .B(n21544), .Z(n21543) );
  XNOR U21584 ( .A(n21545), .B(n21546), .Z(n21499) );
  XNOR U21585 ( .A(n21547), .B(n21548), .Z(n21546) );
  XNOR U21586 ( .A(key[277]), .B(n21549), .Z(n21545) );
  XNOR U21587 ( .A(key[432]), .B(n20152), .Z(n21095) );
  IV U21588 ( .A(n20158), .Z(n20152) );
  XOR U21589 ( .A(n20909), .B(n20973), .Z(n20158) );
  XOR U21590 ( .A(n21551), .B(n20944), .Z(n21550) );
  OR U21591 ( .A(n21552), .B(n21044), .Z(n20944) );
  XNOR U21592 ( .A(n20947), .B(n21043), .Z(n21044) );
  ANDN U21593 ( .B(n21043), .A(n21553), .Z(n21551) );
  XNOR U21594 ( .A(n20942), .B(n21554), .Z(n20909) );
  XNOR U21595 ( .A(n21555), .B(n21026), .Z(n21554) );
  XNOR U21596 ( .A(n21034), .B(n20913), .Z(n21031) );
  ANDN U21597 ( .B(n21557), .A(n21034), .Z(n21555) );
  XOR U21598 ( .A(n21024), .B(n21558), .Z(n20942) );
  XNOR U21599 ( .A(n21559), .B(n21560), .Z(n21558) );
  NAND U21600 ( .A(n21039), .B(n21561), .Z(n21560) );
  XNOR U21601 ( .A(n21562), .B(n21559), .Z(n21024) );
  OR U21602 ( .A(n21047), .B(n21563), .Z(n21559) );
  XNOR U21603 ( .A(n21564), .B(n21039), .Z(n21047) );
  XOR U21604 ( .A(n21043), .B(n20913), .Z(n21039) );
  XOR U21605 ( .A(n21565), .B(n21566), .Z(n20913) );
  NANDN U21606 ( .A(n21567), .B(n21568), .Z(n21566) );
  XOR U21607 ( .A(n21569), .B(n21570), .Z(n21043) );
  NANDN U21608 ( .A(n21567), .B(n21571), .Z(n21570) );
  ANDN U21609 ( .B(n21564), .A(n21572), .Z(n21562) );
  IV U21610 ( .A(n21050), .Z(n21564) );
  XOR U21611 ( .A(n21034), .B(n20947), .Z(n21050) );
  XNOR U21612 ( .A(n21573), .B(n21569), .Z(n20947) );
  NANDN U21613 ( .A(n21574), .B(n21575), .Z(n21569) );
  XOR U21614 ( .A(n21571), .B(n21576), .Z(n21575) );
  ANDN U21615 ( .B(n21576), .A(n21577), .Z(n21573) );
  XOR U21616 ( .A(n21578), .B(n21565), .Z(n21034) );
  NANDN U21617 ( .A(n21574), .B(n21579), .Z(n21565) );
  XOR U21618 ( .A(n21580), .B(n21568), .Z(n21579) );
  XNOR U21619 ( .A(n21581), .B(n21582), .Z(n21567) );
  XOR U21620 ( .A(n21583), .B(n21584), .Z(n21582) );
  XNOR U21621 ( .A(n21585), .B(n21586), .Z(n21581) );
  XNOR U21622 ( .A(n21587), .B(n21588), .Z(n21586) );
  ANDN U21623 ( .B(n21580), .A(n21584), .Z(n21587) );
  ANDN U21624 ( .B(n21580), .A(n21577), .Z(n21578) );
  XNOR U21625 ( .A(n21583), .B(n21589), .Z(n21577) );
  XOR U21626 ( .A(n21590), .B(n21588), .Z(n21589) );
  NAND U21627 ( .A(n21591), .B(n21592), .Z(n21588) );
  XNOR U21628 ( .A(n21585), .B(n21568), .Z(n21592) );
  IV U21629 ( .A(n21580), .Z(n21585) );
  XNOR U21630 ( .A(n21571), .B(n21584), .Z(n21591) );
  IV U21631 ( .A(n21576), .Z(n21584) );
  XOR U21632 ( .A(n21593), .B(n21594), .Z(n21576) );
  XNOR U21633 ( .A(n21595), .B(n21596), .Z(n21594) );
  XNOR U21634 ( .A(n21597), .B(n21598), .Z(n21593) );
  ANDN U21635 ( .B(n21557), .A(n21033), .Z(n21597) );
  AND U21636 ( .A(n21568), .B(n21571), .Z(n21590) );
  XNOR U21637 ( .A(n21568), .B(n21571), .Z(n21583) );
  XNOR U21638 ( .A(n21599), .B(n21600), .Z(n21571) );
  XNOR U21639 ( .A(n21601), .B(n21596), .Z(n21600) );
  XOR U21640 ( .A(n21602), .B(n21603), .Z(n21599) );
  XNOR U21641 ( .A(n21604), .B(n21598), .Z(n21603) );
  OR U21642 ( .A(n21032), .B(n21556), .Z(n21598) );
  XNOR U21643 ( .A(n21557), .B(n21605), .Z(n21556) );
  XNOR U21644 ( .A(n21033), .B(n20914), .Z(n21032) );
  ANDN U21645 ( .B(n21606), .A(n21028), .Z(n21604) );
  XNOR U21646 ( .A(n21607), .B(n21608), .Z(n21568) );
  XNOR U21647 ( .A(n21596), .B(n21609), .Z(n21608) );
  XOR U21648 ( .A(n21023), .B(n21602), .Z(n21609) );
  XNOR U21649 ( .A(n21557), .B(n21033), .Z(n21596) );
  XOR U21650 ( .A(n20946), .B(n21610), .Z(n21607) );
  XNOR U21651 ( .A(n21611), .B(n21612), .Z(n21610) );
  ANDN U21652 ( .B(n21613), .A(n21553), .Z(n21611) );
  XNOR U21653 ( .A(n21614), .B(n21615), .Z(n21580) );
  XNOR U21654 ( .A(n21601), .B(n21616), .Z(n21615) );
  XNOR U21655 ( .A(n21042), .B(n21595), .Z(n21616) );
  XOR U21656 ( .A(n21602), .B(n21617), .Z(n21595) );
  XNOR U21657 ( .A(n21618), .B(n21619), .Z(n21617) );
  NAND U21658 ( .A(n21561), .B(n21038), .Z(n21619) );
  XNOR U21659 ( .A(n21620), .B(n21618), .Z(n21602) );
  NANDN U21660 ( .A(n21563), .B(n21048), .Z(n21618) );
  XOR U21661 ( .A(n21049), .B(n21038), .Z(n21048) );
  XNOR U21662 ( .A(n21613), .B(n20914), .Z(n21038) );
  XOR U21663 ( .A(n21572), .B(n21561), .Z(n21563) );
  XNOR U21664 ( .A(n21553), .B(n21605), .Z(n21561) );
  ANDN U21665 ( .B(n21049), .A(n21572), .Z(n21620) );
  XOR U21666 ( .A(n20946), .B(n21557), .Z(n21572) );
  XNOR U21667 ( .A(n21621), .B(n21622), .Z(n21557) );
  XNOR U21668 ( .A(n21623), .B(n21624), .Z(n21622) );
  XOR U21669 ( .A(n21605), .B(n21606), .Z(n21601) );
  IV U21670 ( .A(n20914), .Z(n21606) );
  XOR U21671 ( .A(n21625), .B(n21626), .Z(n20914) );
  XOR U21672 ( .A(n21627), .B(n21624), .Z(n21626) );
  IV U21673 ( .A(n21028), .Z(n21605) );
  XOR U21674 ( .A(n21624), .B(n21628), .Z(n21028) );
  XNOR U21675 ( .A(n21629), .B(n21630), .Z(n21614) );
  XNOR U21676 ( .A(n21631), .B(n21612), .Z(n21630) );
  OR U21677 ( .A(n21045), .B(n21552), .Z(n21612) );
  XNOR U21678 ( .A(n20946), .B(n21553), .Z(n21552) );
  IV U21679 ( .A(n21629), .Z(n21553) );
  XOR U21680 ( .A(n21023), .B(n21613), .Z(n21045) );
  IV U21681 ( .A(n21042), .Z(n21613) );
  XNOR U21682 ( .A(n21633), .B(n21621), .Z(n21632) );
  XOR U21683 ( .A(n21634), .B(n21635), .Z(n21621) );
  XNOR U21684 ( .A(n21636), .B(n21637), .Z(n21635) );
  XOR U21685 ( .A(n21638), .B(n21639), .Z(n21634) );
  XNOR U21686 ( .A(key[314]), .B(n21640), .Z(n21639) );
  XOR U21687 ( .A(n21625), .B(n21641), .Z(n21033) );
  XOR U21688 ( .A(n21624), .B(n21642), .Z(n21641) );
  NOR U21689 ( .A(n21023), .B(n20946), .Z(n21631) );
  XOR U21690 ( .A(n21625), .B(n21643), .Z(n21023) );
  XOR U21691 ( .A(n21624), .B(n21644), .Z(n21643) );
  XOR U21692 ( .A(n21645), .B(n21646), .Z(n21624) );
  XOR U21693 ( .A(n20946), .B(n21647), .Z(n21646) );
  XOR U21694 ( .A(n21648), .B(n21649), .Z(n21645) );
  XNOR U21695 ( .A(key[318]), .B(n21650), .Z(n21649) );
  IV U21696 ( .A(n21628), .Z(n21625) );
  XOR U21697 ( .A(n21651), .B(n21652), .Z(n21628) );
  XNOR U21698 ( .A(n21653), .B(n21654), .Z(n21652) );
  XOR U21699 ( .A(n21655), .B(n21656), .Z(n21651) );
  XOR U21700 ( .A(key[317]), .B(n21657), .Z(n21656) );
  XOR U21701 ( .A(n21658), .B(n21659), .Z(n21629) );
  XNOR U21702 ( .A(n21644), .B(n21642), .Z(n21659) );
  XNOR U21703 ( .A(n21660), .B(n21661), .Z(n21642) );
  XOR U21704 ( .A(n21662), .B(n21663), .Z(n21661) );
  XNOR U21705 ( .A(key[319]), .B(n21664), .Z(n21660) );
  XNOR U21706 ( .A(n21665), .B(n21666), .Z(n21644) );
  XNOR U21707 ( .A(n21667), .B(n21668), .Z(n21666) );
  XNOR U21708 ( .A(n21669), .B(n21670), .Z(n21665) );
  XNOR U21709 ( .A(key[316]), .B(n21671), .Z(n21670) );
  XNOR U21710 ( .A(n20946), .B(n21623), .Z(n21658) );
  XOR U21711 ( .A(n21672), .B(n21673), .Z(n21623) );
  XNOR U21712 ( .A(n21674), .B(n21675), .Z(n21673) );
  XNOR U21713 ( .A(n21676), .B(n21633), .Z(n21675) );
  IV U21714 ( .A(n21627), .Z(n21633) );
  XNOR U21715 ( .A(n21677), .B(n21678), .Z(n21627) );
  XOR U21716 ( .A(n21679), .B(n21680), .Z(n21678) );
  XNOR U21717 ( .A(n21681), .B(n21682), .Z(n21677) );
  XOR U21718 ( .A(key[313]), .B(n21683), .Z(n21682) );
  XNOR U21719 ( .A(n21684), .B(n21685), .Z(n21672) );
  XNOR U21720 ( .A(key[315]), .B(n21686), .Z(n21685) );
  XNOR U21721 ( .A(n21687), .B(n21688), .Z(n20946) );
  XOR U21722 ( .A(n21689), .B(n21690), .Z(n21688) );
  XNOR U21723 ( .A(n21691), .B(n21692), .Z(n21687) );
  XOR U21724 ( .A(key[312]), .B(n21693), .Z(n21692) );
  XNOR U21725 ( .A(n17102), .B(n21694), .Z(n20758) );
  XOR U21726 ( .A(key[586]), .B(n15347), .Z(n21694) );
  XNOR U21727 ( .A(n15309), .B(n16040), .Z(n15347) );
  XOR U21728 ( .A(n20667), .B(n20659), .Z(n16040) );
  XOR U21729 ( .A(n20752), .B(n21695), .Z(n20659) );
  XNOR U21730 ( .A(n20749), .B(n21696), .Z(n21695) );
  NAND U21731 ( .A(n21697), .B(n20565), .Z(n21696) );
  NANDN U21732 ( .A(n21698), .B(n20767), .Z(n20749) );
  XOR U21733 ( .A(n20750), .B(n20565), .Z(n20767) );
  XOR U21734 ( .A(n20752), .B(n21699), .Z(n20667) );
  XOR U21735 ( .A(n21700), .B(n20655), .Z(n21699) );
  OR U21736 ( .A(n21701), .B(n20778), .Z(n20655) );
  XOR U21737 ( .A(n20657), .B(n20781), .Z(n20778) );
  ANDN U21738 ( .B(n20781), .A(n21702), .Z(n21700) );
  XOR U21739 ( .A(n21703), .B(n20754), .Z(n20752) );
  OR U21740 ( .A(n20783), .B(n21704), .Z(n20754) );
  XOR U21741 ( .A(n21705), .B(n20756), .Z(n20783) );
  XNOR U21742 ( .A(n20781), .B(n20565), .Z(n20756) );
  XOR U21743 ( .A(n21706), .B(n21707), .Z(n20565) );
  NANDN U21744 ( .A(n21708), .B(n21709), .Z(n21707) );
  XOR U21745 ( .A(n21710), .B(n21711), .Z(n20781) );
  OR U21746 ( .A(n21708), .B(n21712), .Z(n21711) );
  ANDN U21747 ( .B(n21705), .A(n21713), .Z(n21703) );
  IV U21748 ( .A(n20786), .Z(n21705) );
  XOR U21749 ( .A(n20657), .B(n20750), .Z(n20786) );
  XNOR U21750 ( .A(n21714), .B(n21706), .Z(n20750) );
  NANDN U21751 ( .A(n21715), .B(n21716), .Z(n21706) );
  ANDN U21752 ( .B(n21717), .A(n21718), .Z(n21714) );
  NANDN U21753 ( .A(n21715), .B(n21720), .Z(n21710) );
  XOR U21754 ( .A(n21721), .B(n21708), .Z(n21715) );
  XNOR U21755 ( .A(n21722), .B(n21723), .Z(n21708) );
  XOR U21756 ( .A(n21724), .B(n21717), .Z(n21723) );
  XNOR U21757 ( .A(n21725), .B(n21726), .Z(n21722) );
  XNOR U21758 ( .A(n21727), .B(n21728), .Z(n21726) );
  ANDN U21759 ( .B(n21717), .A(n21729), .Z(n21727) );
  IV U21760 ( .A(n21730), .Z(n21717) );
  ANDN U21761 ( .B(n21721), .A(n21729), .Z(n21719) );
  IV U21762 ( .A(n21725), .Z(n21729) );
  IV U21763 ( .A(n21718), .Z(n21721) );
  XNOR U21764 ( .A(n21724), .B(n21731), .Z(n21718) );
  XOR U21765 ( .A(n21732), .B(n21728), .Z(n21731) );
  NAND U21766 ( .A(n21720), .B(n21716), .Z(n21728) );
  XNOR U21767 ( .A(n21709), .B(n21730), .Z(n21716) );
  XOR U21768 ( .A(n21733), .B(n21734), .Z(n21730) );
  XOR U21769 ( .A(n21735), .B(n21736), .Z(n21734) );
  XNOR U21770 ( .A(n20780), .B(n21737), .Z(n21736) );
  XNOR U21771 ( .A(n21738), .B(n21739), .Z(n21733) );
  XNOR U21772 ( .A(n21740), .B(n21741), .Z(n21739) );
  ANDN U21773 ( .B(n21742), .A(n20658), .Z(n21740) );
  XNOR U21774 ( .A(n21725), .B(n21712), .Z(n21720) );
  XOR U21775 ( .A(n21743), .B(n21744), .Z(n21725) );
  XNOR U21776 ( .A(n21745), .B(n21737), .Z(n21744) );
  XOR U21777 ( .A(n21746), .B(n21747), .Z(n21737) );
  XNOR U21778 ( .A(n21748), .B(n21749), .Z(n21747) );
  NAND U21779 ( .A(n20757), .B(n20775), .Z(n21749) );
  XNOR U21780 ( .A(n21750), .B(n21751), .Z(n21743) );
  ANDN U21781 ( .B(n21752), .A(n20751), .Z(n21750) );
  ANDN U21782 ( .B(n21709), .A(n21712), .Z(n21732) );
  XOR U21783 ( .A(n21712), .B(n21709), .Z(n21724) );
  XNOR U21784 ( .A(n21753), .B(n21754), .Z(n21709) );
  XNOR U21785 ( .A(n21746), .B(n21755), .Z(n21754) );
  XOR U21786 ( .A(n21745), .B(n20771), .Z(n21755) );
  XOR U21787 ( .A(n20658), .B(n21756), .Z(n21753) );
  XNOR U21788 ( .A(n21757), .B(n21741), .Z(n21756) );
  OR U21789 ( .A(n20779), .B(n21701), .Z(n21741) );
  XNOR U21790 ( .A(n20658), .B(n21702), .Z(n21701) );
  XOR U21791 ( .A(n20771), .B(n20780), .Z(n20779) );
  ANDN U21792 ( .B(n20780), .A(n21702), .Z(n21757) );
  XOR U21793 ( .A(n21758), .B(n21759), .Z(n21712) );
  XOR U21794 ( .A(n21746), .B(n21735), .Z(n21759) );
  XOR U21795 ( .A(n21697), .B(n20566), .Z(n21735) );
  XOR U21796 ( .A(n21760), .B(n21748), .Z(n21746) );
  NANDN U21797 ( .A(n21704), .B(n20784), .Z(n21748) );
  XOR U21798 ( .A(n20785), .B(n20775), .Z(n20784) );
  XNOR U21799 ( .A(n21752), .B(n21761), .Z(n20780) );
  XOR U21800 ( .A(n21762), .B(n21763), .Z(n21761) );
  XOR U21801 ( .A(n21713), .B(n20757), .Z(n21704) );
  XNOR U21802 ( .A(n21702), .B(n21697), .Z(n20757) );
  IV U21803 ( .A(n21738), .Z(n21702) );
  XOR U21804 ( .A(n21764), .B(n21765), .Z(n21738) );
  XOR U21805 ( .A(n21766), .B(n21767), .Z(n21765) );
  XNOR U21806 ( .A(n20658), .B(n21768), .Z(n21764) );
  ANDN U21807 ( .B(n20785), .A(n21713), .Z(n21760) );
  XNOR U21808 ( .A(n20658), .B(n20751), .Z(n21713) );
  XOR U21809 ( .A(n21752), .B(n21742), .Z(n20785) );
  IV U21810 ( .A(n20771), .Z(n21742) );
  XOR U21811 ( .A(n21769), .B(n21770), .Z(n20771) );
  XOR U21812 ( .A(n21771), .B(n21767), .Z(n21770) );
  XNOR U21813 ( .A(n21772), .B(n21773), .Z(n21767) );
  XOR U21814 ( .A(n19517), .B(n18344), .Z(n21773) );
  XOR U21815 ( .A(n20410), .B(n19515), .Z(n18344) );
  XNOR U21816 ( .A(n21774), .B(n18364), .Z(n19515) );
  XOR U21817 ( .A(n21775), .B(n19550), .Z(n20410) );
  IV U21818 ( .A(n21776), .Z(n19550) );
  XOR U21819 ( .A(n19558), .B(n18330), .Z(n19517) );
  XNOR U21820 ( .A(n21777), .B(n21778), .Z(n18330) );
  XNOR U21821 ( .A(n21779), .B(n21780), .Z(n21778) );
  XNOR U21822 ( .A(n21781), .B(n21782), .Z(n21777) );
  XOR U21823 ( .A(n21783), .B(n21784), .Z(n21782) );
  ANDN U21824 ( .B(n21785), .A(n21786), .Z(n21784) );
  XNOR U21825 ( .A(n18346), .B(n21787), .Z(n21772) );
  XOR U21826 ( .A(key[484]), .B(n20418), .Z(n21787) );
  XOR U21827 ( .A(n21788), .B(n20435), .Z(n18346) );
  IV U21828 ( .A(n20765), .Z(n21752) );
  XOR U21829 ( .A(n21745), .B(n21789), .Z(n21758) );
  XNOR U21830 ( .A(n21790), .B(n21751), .Z(n21789) );
  OR U21831 ( .A(n20766), .B(n21698), .Z(n21751) );
  XNOR U21832 ( .A(n21791), .B(n21697), .Z(n21698) );
  XNOR U21833 ( .A(n20765), .B(n20566), .Z(n20766) );
  ANDN U21834 ( .B(n21697), .A(n20566), .Z(n21790) );
  XOR U21835 ( .A(n21769), .B(n21792), .Z(n20566) );
  XNOR U21836 ( .A(n21793), .B(n21771), .Z(n21792) );
  XOR U21837 ( .A(n21771), .B(n21769), .Z(n21697) );
  XNOR U21838 ( .A(n20751), .B(n20765), .Z(n21745) );
  XOR U21839 ( .A(n21769), .B(n21794), .Z(n20765) );
  XNOR U21840 ( .A(n21771), .B(n21766), .Z(n21794) );
  XOR U21841 ( .A(n21795), .B(n21796), .Z(n21766) );
  XOR U21842 ( .A(n21797), .B(n18340), .Z(n21796) );
  XNOR U21843 ( .A(n20440), .B(n19532), .Z(n18340) );
  XOR U21844 ( .A(n21798), .B(n21799), .Z(n19532) );
  XNOR U21845 ( .A(n21800), .B(n21801), .Z(n21799) );
  XNOR U21846 ( .A(n21802), .B(n21803), .Z(n21798) );
  XNOR U21847 ( .A(n21804), .B(n21805), .Z(n20440) );
  XOR U21848 ( .A(n21806), .B(n21807), .Z(n21805) );
  XOR U21849 ( .A(n21808), .B(n21809), .Z(n21804) );
  XNOR U21850 ( .A(key[487]), .B(n19558), .Z(n21795) );
  XNOR U21851 ( .A(n21810), .B(n21811), .Z(n21769) );
  XOR U21852 ( .A(n18331), .B(n20427), .Z(n21811) );
  XOR U21853 ( .A(n18332), .B(n19524), .Z(n20427) );
  IV U21854 ( .A(n18354), .Z(n19524) );
  XOR U21855 ( .A(n21812), .B(n21813), .Z(n18354) );
  XNOR U21856 ( .A(n19526), .B(n20420), .Z(n18331) );
  XNOR U21857 ( .A(n21814), .B(n21815), .Z(n20420) );
  XNOR U21858 ( .A(n21816), .B(n21807), .Z(n21815) );
  XNOR U21859 ( .A(n21817), .B(n21818), .Z(n21807) );
  XNOR U21860 ( .A(n21819), .B(n21820), .Z(n21818) );
  NANDN U21861 ( .A(n21821), .B(n21822), .Z(n21820) );
  XNOR U21862 ( .A(n21775), .B(n21823), .Z(n21814) );
  XOR U21863 ( .A(n21824), .B(n21825), .Z(n21823) );
  ANDN U21864 ( .B(n21826), .A(n21827), .Z(n21825) );
  XNOR U21865 ( .A(n21828), .B(n21829), .Z(n19526) );
  XNOR U21866 ( .A(n21830), .B(n21801), .Z(n21829) );
  XNOR U21867 ( .A(n21831), .B(n21832), .Z(n21801) );
  XNOR U21868 ( .A(n21833), .B(n21834), .Z(n21832) );
  NANDN U21869 ( .A(n21835), .B(n21836), .Z(n21834) );
  XNOR U21870 ( .A(n21774), .B(n21837), .Z(n21828) );
  XOR U21871 ( .A(n21838), .B(n21839), .Z(n21837) );
  ANDN U21872 ( .B(n21840), .A(n21841), .Z(n21839) );
  XOR U21873 ( .A(key[485]), .B(n20435), .Z(n21810) );
  XNOR U21874 ( .A(n21842), .B(n21843), .Z(n20435) );
  XNOR U21875 ( .A(n21844), .B(n21845), .Z(n21843) );
  XOR U21876 ( .A(n21846), .B(n21847), .Z(n21842) );
  XOR U21877 ( .A(n21848), .B(n21849), .Z(n21847) );
  ANDN U21878 ( .B(n21850), .A(n21851), .Z(n21849) );
  IV U21879 ( .A(n21791), .Z(n20751) );
  XNOR U21880 ( .A(n21762), .B(n21768), .Z(n21852) );
  XOR U21881 ( .A(n21853), .B(n21854), .Z(n21768) );
  XOR U21882 ( .A(n18360), .B(n21855), .Z(n21854) );
  XOR U21883 ( .A(n19553), .B(n21763), .Z(n21855) );
  IV U21884 ( .A(n21793), .Z(n21763) );
  XOR U21885 ( .A(n21856), .B(n21857), .Z(n21793) );
  XOR U21886 ( .A(n19536), .B(n18365), .Z(n21857) );
  XOR U21887 ( .A(n19559), .B(n18381), .Z(n18365) );
  XOR U21888 ( .A(n21800), .B(n21858), .Z(n18381) );
  XNOR U21889 ( .A(n21859), .B(n21803), .Z(n21858) );
  XOR U21890 ( .A(n21806), .B(n21860), .Z(n19559) );
  XNOR U21891 ( .A(n21808), .B(n21809), .Z(n21860) );
  XOR U21892 ( .A(n18366), .B(n18374), .Z(n19536) );
  XNOR U21893 ( .A(key[481]), .B(n18385), .Z(n21856) );
  XNOR U21894 ( .A(n19558), .B(n18348), .Z(n19553) );
  XOR U21895 ( .A(n21779), .B(n18374), .Z(n18348) );
  XOR U21896 ( .A(n21861), .B(n21862), .Z(n18374) );
  XOR U21897 ( .A(n19537), .B(n18375), .Z(n18360) );
  XNOR U21898 ( .A(n21863), .B(n21864), .Z(n18375) );
  XOR U21899 ( .A(n21800), .B(n21865), .Z(n21864) );
  XNOR U21900 ( .A(n21866), .B(n21867), .Z(n21800) );
  XNOR U21901 ( .A(n21868), .B(n21869), .Z(n21867) );
  NANDN U21902 ( .A(n21870), .B(n21836), .Z(n21869) );
  XNOR U21903 ( .A(n21859), .B(n21871), .Z(n21863) );
  IV U21904 ( .A(n20411), .Z(n19537) );
  XOR U21905 ( .A(n21872), .B(n21873), .Z(n20411) );
  XNOR U21906 ( .A(n21874), .B(n21875), .Z(n21873) );
  XOR U21907 ( .A(n21876), .B(n21877), .Z(n21809) );
  XNOR U21908 ( .A(n21878), .B(n21879), .Z(n21877) );
  NANDN U21909 ( .A(n21880), .B(n21822), .Z(n21879) );
  XNOR U21910 ( .A(n18369), .B(n21881), .Z(n21853) );
  XNOR U21911 ( .A(key[483]), .B(n18378), .Z(n21881) );
  XNOR U21912 ( .A(n20431), .B(n20418), .Z(n18369) );
  XNOR U21913 ( .A(n21844), .B(n18366), .Z(n20418) );
  XOR U21914 ( .A(n21882), .B(n21883), .Z(n21762) );
  XNOR U21915 ( .A(n19555), .B(n18376), .Z(n21883) );
  XOR U21916 ( .A(n21776), .B(n18364), .Z(n18376) );
  XOR U21917 ( .A(n21884), .B(n21859), .Z(n18364) );
  IV U21918 ( .A(n21802), .Z(n21859) );
  XOR U21919 ( .A(n21886), .B(n21887), .Z(n21885) );
  NANDN U21920 ( .A(n21888), .B(n21840), .Z(n21887) );
  XOR U21921 ( .A(n21890), .B(n21808), .Z(n21776) );
  XOR U21922 ( .A(n21891), .B(n21892), .Z(n21808) );
  XOR U21923 ( .A(n21893), .B(n21894), .Z(n21892) );
  NANDN U21924 ( .A(n21895), .B(n21826), .Z(n21894) );
  XOR U21925 ( .A(n18378), .B(n18371), .Z(n19555) );
  XOR U21926 ( .A(n21896), .B(n21897), .Z(n18371) );
  XNOR U21927 ( .A(n21898), .B(n21813), .Z(n21897) );
  XNOR U21928 ( .A(n21899), .B(n21900), .Z(n21813) );
  XNOR U21929 ( .A(n21901), .B(n21783), .Z(n21900) );
  ANDN U21930 ( .B(n21902), .A(n21903), .Z(n21783) );
  NOR U21931 ( .A(n21904), .B(n21905), .Z(n21901) );
  XOR U21932 ( .A(n21861), .B(n21906), .Z(n21896) );
  XOR U21933 ( .A(n21907), .B(n21908), .Z(n18378) );
  XOR U21934 ( .A(n21909), .B(n21910), .Z(n21908) );
  XNOR U21935 ( .A(n21911), .B(n21912), .Z(n21907) );
  XOR U21936 ( .A(key[482]), .B(n18366), .Z(n21882) );
  XOR U21937 ( .A(n21913), .B(n21912), .Z(n18366) );
  XOR U21938 ( .A(n21914), .B(n21915), .Z(n21771) );
  XOR U21939 ( .A(n18356), .B(n18332), .Z(n21915) );
  XNOR U21940 ( .A(n21916), .B(n21910), .Z(n18332) );
  XNOR U21941 ( .A(n21917), .B(n21918), .Z(n21910) );
  XNOR U21942 ( .A(n21919), .B(n21848), .Z(n21918) );
  ANDN U21943 ( .B(n21920), .A(n21921), .Z(n21848) );
  NOR U21944 ( .A(n21922), .B(n21923), .Z(n21919) );
  XOR U21945 ( .A(n21797), .B(n20436), .Z(n18356) );
  XNOR U21946 ( .A(n18334), .B(n19528), .Z(n20436) );
  XNOR U21947 ( .A(n21806), .B(n21875), .Z(n19528) );
  XOR U21948 ( .A(n21876), .B(n21924), .Z(n21875) );
  XNOR U21949 ( .A(n21925), .B(n21824), .Z(n21924) );
  ANDN U21950 ( .B(n21926), .A(n21927), .Z(n21824) );
  NOR U21951 ( .A(n21928), .B(n21929), .Z(n21925) );
  XNOR U21952 ( .A(n21816), .B(n21930), .Z(n21876) );
  XNOR U21953 ( .A(n21931), .B(n21932), .Z(n21930) );
  NAND U21954 ( .A(n21933), .B(n21934), .Z(n21932) );
  XOR U21955 ( .A(n21890), .B(n21874), .Z(n21806) );
  XOR U21956 ( .A(n21816), .B(n21935), .Z(n21874) );
  XNOR U21957 ( .A(n21878), .B(n21936), .Z(n21935) );
  NANDN U21958 ( .A(n21937), .B(n21938), .Z(n21936) );
  OR U21959 ( .A(n21939), .B(n21940), .Z(n21878) );
  XOR U21960 ( .A(n21941), .B(n21931), .Z(n21816) );
  NANDN U21961 ( .A(n21942), .B(n21943), .Z(n21931) );
  ANDN U21962 ( .B(n21944), .A(n21945), .Z(n21941) );
  XOR U21963 ( .A(n21803), .B(n21865), .Z(n18334) );
  XOR U21964 ( .A(n21866), .B(n21946), .Z(n21865) );
  XNOR U21965 ( .A(n21947), .B(n21838), .Z(n21946) );
  ANDN U21966 ( .B(n21948), .A(n21949), .Z(n21838) );
  NOR U21967 ( .A(n21950), .B(n21951), .Z(n21947) );
  XNOR U21968 ( .A(n21830), .B(n21952), .Z(n21866) );
  XNOR U21969 ( .A(n21953), .B(n21954), .Z(n21952) );
  NAND U21970 ( .A(n21955), .B(n21956), .Z(n21954) );
  XNOR U21971 ( .A(n21957), .B(n21871), .Z(n21803) );
  XOR U21972 ( .A(n21830), .B(n21958), .Z(n21871) );
  XNOR U21973 ( .A(n21868), .B(n21959), .Z(n21958) );
  NANDN U21974 ( .A(n21960), .B(n21961), .Z(n21959) );
  OR U21975 ( .A(n21962), .B(n21963), .Z(n21868) );
  XOR U21976 ( .A(n21964), .B(n21953), .Z(n21830) );
  NANDN U21977 ( .A(n21965), .B(n21966), .Z(n21953) );
  ANDN U21978 ( .B(n21967), .A(n21968), .Z(n21964) );
  XOR U21979 ( .A(n21788), .B(n20439), .Z(n21797) );
  XNOR U21980 ( .A(n21969), .B(n21970), .Z(n20439) );
  XNOR U21981 ( .A(n21909), .B(n21845), .Z(n21970) );
  XNOR U21982 ( .A(n21971), .B(n21972), .Z(n21845) );
  XNOR U21983 ( .A(n21973), .B(n21974), .Z(n21972) );
  NANDN U21984 ( .A(n21975), .B(n21976), .Z(n21974) );
  XOR U21985 ( .A(n21916), .B(n21912), .Z(n21969) );
  IV U21986 ( .A(n20431), .Z(n21788) );
  XNOR U21987 ( .A(n19543), .B(n21977), .Z(n21914) );
  XOR U21988 ( .A(key[486]), .B(n20658), .Z(n21977) );
  XNOR U21989 ( .A(n21978), .B(n21979), .Z(n20658) );
  XOR U21990 ( .A(n18341), .B(n20409), .Z(n21979) );
  XNOR U21991 ( .A(n21890), .B(n21775), .Z(n20409) );
  XNOR U21992 ( .A(n21817), .B(n21980), .Z(n21775) );
  XNOR U21993 ( .A(n21981), .B(n21893), .Z(n21980) );
  XNOR U21994 ( .A(n21929), .B(n21826), .Z(n21926) );
  ANDN U21995 ( .B(n21983), .A(n21929), .Z(n21981) );
  XNOR U21996 ( .A(n21891), .B(n21984), .Z(n21817) );
  XNOR U21997 ( .A(n21985), .B(n21986), .Z(n21984) );
  NAND U21998 ( .A(n21934), .B(n21987), .Z(n21986) );
  XOR U21999 ( .A(n21891), .B(n21988), .Z(n21890) );
  XOR U22000 ( .A(n21989), .B(n21819), .Z(n21988) );
  OR U22001 ( .A(n21990), .B(n21939), .Z(n21819) );
  XNOR U22002 ( .A(n21822), .B(n21938), .Z(n21939) );
  ANDN U22003 ( .B(n21991), .A(n21992), .Z(n21989) );
  XOR U22004 ( .A(n21993), .B(n21985), .Z(n21891) );
  OR U22005 ( .A(n21942), .B(n21994), .Z(n21985) );
  XNOR U22006 ( .A(n21995), .B(n21934), .Z(n21942) );
  XOR U22007 ( .A(n21938), .B(n21826), .Z(n21934) );
  XOR U22008 ( .A(n21996), .B(n21997), .Z(n21826) );
  NANDN U22009 ( .A(n21998), .B(n21999), .Z(n21997) );
  IV U22010 ( .A(n21992), .Z(n21938) );
  XNOR U22011 ( .A(n22000), .B(n22001), .Z(n21992) );
  NANDN U22012 ( .A(n21998), .B(n22002), .Z(n22001) );
  ANDN U22013 ( .B(n21995), .A(n22003), .Z(n21993) );
  IV U22014 ( .A(n21945), .Z(n21995) );
  XOR U22015 ( .A(n21929), .B(n21822), .Z(n21945) );
  XNOR U22016 ( .A(n22004), .B(n22000), .Z(n21822) );
  NANDN U22017 ( .A(n22005), .B(n22006), .Z(n22000) );
  XOR U22018 ( .A(n22002), .B(n22007), .Z(n22006) );
  ANDN U22019 ( .B(n22007), .A(n22008), .Z(n22004) );
  XOR U22020 ( .A(n22009), .B(n21996), .Z(n21929) );
  NANDN U22021 ( .A(n22005), .B(n22010), .Z(n21996) );
  XOR U22022 ( .A(n22011), .B(n21999), .Z(n22010) );
  XNOR U22023 ( .A(n22012), .B(n22013), .Z(n21998) );
  XOR U22024 ( .A(n22014), .B(n22015), .Z(n22013) );
  XNOR U22025 ( .A(n22016), .B(n22017), .Z(n22012) );
  XNOR U22026 ( .A(n22018), .B(n22019), .Z(n22017) );
  ANDN U22027 ( .B(n22011), .A(n22015), .Z(n22018) );
  ANDN U22028 ( .B(n22011), .A(n22008), .Z(n22009) );
  XNOR U22029 ( .A(n22014), .B(n22020), .Z(n22008) );
  XOR U22030 ( .A(n22021), .B(n22019), .Z(n22020) );
  NAND U22031 ( .A(n22022), .B(n22023), .Z(n22019) );
  XNOR U22032 ( .A(n22016), .B(n21999), .Z(n22023) );
  IV U22033 ( .A(n22011), .Z(n22016) );
  XNOR U22034 ( .A(n22002), .B(n22015), .Z(n22022) );
  IV U22035 ( .A(n22007), .Z(n22015) );
  XOR U22036 ( .A(n22024), .B(n22025), .Z(n22007) );
  XNOR U22037 ( .A(n22026), .B(n22027), .Z(n22025) );
  XNOR U22038 ( .A(n22028), .B(n22029), .Z(n22024) );
  ANDN U22039 ( .B(n21983), .A(n21928), .Z(n22028) );
  AND U22040 ( .A(n21999), .B(n22002), .Z(n22021) );
  XNOR U22041 ( .A(n21999), .B(n22002), .Z(n22014) );
  XNOR U22042 ( .A(n22030), .B(n22031), .Z(n22002) );
  XNOR U22043 ( .A(n22032), .B(n22027), .Z(n22031) );
  XOR U22044 ( .A(n22033), .B(n22034), .Z(n22030) );
  XNOR U22045 ( .A(n22035), .B(n22029), .Z(n22034) );
  OR U22046 ( .A(n21927), .B(n21982), .Z(n22029) );
  XNOR U22047 ( .A(n21983), .B(n22036), .Z(n21982) );
  XNOR U22048 ( .A(n21928), .B(n21827), .Z(n21927) );
  ANDN U22049 ( .B(n22037), .A(n21895), .Z(n22035) );
  XNOR U22050 ( .A(n22038), .B(n22039), .Z(n21999) );
  XNOR U22051 ( .A(n22027), .B(n22040), .Z(n22039) );
  XOR U22052 ( .A(n21880), .B(n22033), .Z(n22040) );
  XNOR U22053 ( .A(n21983), .B(n21928), .Z(n22027) );
  XNOR U22054 ( .A(n22041), .B(n22042), .Z(n22038) );
  XNOR U22055 ( .A(n22043), .B(n22044), .Z(n22042) );
  ANDN U22056 ( .B(n21991), .A(n21937), .Z(n22043) );
  XNOR U22057 ( .A(n22045), .B(n22046), .Z(n22011) );
  XNOR U22058 ( .A(n22032), .B(n22047), .Z(n22046) );
  XNOR U22059 ( .A(n21937), .B(n22026), .Z(n22047) );
  XOR U22060 ( .A(n22033), .B(n22048), .Z(n22026) );
  XNOR U22061 ( .A(n22049), .B(n22050), .Z(n22048) );
  NAND U22062 ( .A(n21987), .B(n21933), .Z(n22050) );
  XNOR U22063 ( .A(n22051), .B(n22049), .Z(n22033) );
  NANDN U22064 ( .A(n21994), .B(n21943), .Z(n22049) );
  XOR U22065 ( .A(n21944), .B(n21933), .Z(n21943) );
  XNOR U22066 ( .A(n22052), .B(n21827), .Z(n21933) );
  XOR U22067 ( .A(n22003), .B(n21987), .Z(n21994) );
  XOR U22068 ( .A(n21991), .B(n22036), .Z(n21987) );
  ANDN U22069 ( .B(n21944), .A(n22003), .Z(n22051) );
  XNOR U22070 ( .A(n22041), .B(n21983), .Z(n22003) );
  XNOR U22071 ( .A(n22053), .B(n22054), .Z(n21983) );
  XNOR U22072 ( .A(n22055), .B(n22056), .Z(n22054) );
  XOR U22073 ( .A(n22057), .B(n22058), .Z(n21944) );
  XOR U22074 ( .A(n22036), .B(n22037), .Z(n22032) );
  IV U22075 ( .A(n21827), .Z(n22037) );
  XOR U22076 ( .A(n22059), .B(n22060), .Z(n21827) );
  XNOR U22077 ( .A(n22061), .B(n22056), .Z(n22060) );
  IV U22078 ( .A(n21895), .Z(n22036) );
  XOR U22079 ( .A(n22056), .B(n22062), .Z(n21895) );
  XNOR U22080 ( .A(n21991), .B(n22063), .Z(n22045) );
  XNOR U22081 ( .A(n22064), .B(n22044), .Z(n22063) );
  OR U22082 ( .A(n21940), .B(n21990), .Z(n22044) );
  XNOR U22083 ( .A(n22041), .B(n21991), .Z(n21990) );
  XOR U22084 ( .A(n21880), .B(n22052), .Z(n21940) );
  IV U22085 ( .A(n21937), .Z(n22052) );
  XOR U22086 ( .A(n22058), .B(n22065), .Z(n21937) );
  XNOR U22087 ( .A(n22061), .B(n22053), .Z(n22065) );
  XOR U22088 ( .A(n22066), .B(n22067), .Z(n22053) );
  XNOR U22089 ( .A(n21676), .B(n21680), .Z(n22067) );
  XNOR U22090 ( .A(n22068), .B(n22069), .Z(n22066) );
  XNOR U22091 ( .A(key[298]), .B(n22070), .Z(n22069) );
  IV U22092 ( .A(n21928), .Z(n22058) );
  XOR U22093 ( .A(n22059), .B(n22071), .Z(n21928) );
  XOR U22094 ( .A(n22056), .B(n22072), .Z(n22071) );
  ANDN U22095 ( .B(n22057), .A(n21821), .Z(n22064) );
  IV U22096 ( .A(n21880), .Z(n22057) );
  XOR U22097 ( .A(n22059), .B(n22073), .Z(n21880) );
  XOR U22098 ( .A(n22056), .B(n22074), .Z(n22073) );
  XOR U22099 ( .A(n22075), .B(n22076), .Z(n22056) );
  XNOR U22100 ( .A(n22077), .B(n21821), .Z(n22076) );
  IV U22101 ( .A(n22041), .Z(n21821) );
  XOR U22102 ( .A(n21655), .B(n22078), .Z(n22075) );
  XNOR U22103 ( .A(key[302]), .B(n22079), .Z(n22078) );
  IV U22104 ( .A(n22062), .Z(n22059) );
  XOR U22105 ( .A(n22080), .B(n22081), .Z(n22062) );
  XNOR U22106 ( .A(n22082), .B(n22083), .Z(n22081) );
  XOR U22107 ( .A(n21648), .B(n22084), .Z(n22080) );
  XOR U22108 ( .A(key[301]), .B(n22085), .Z(n22084) );
  XOR U22109 ( .A(n22086), .B(n22087), .Z(n21991) );
  XNOR U22110 ( .A(n22074), .B(n22072), .Z(n22087) );
  XNOR U22111 ( .A(n22088), .B(n22089), .Z(n22072) );
  XNOR U22112 ( .A(n21690), .B(n22090), .Z(n22089) );
  XOR U22113 ( .A(key[303]), .B(n22091), .Z(n22088) );
  XNOR U22114 ( .A(n22092), .B(n22093), .Z(n22074) );
  XNOR U22115 ( .A(n22094), .B(n22095), .Z(n22092) );
  XNOR U22116 ( .A(key[300]), .B(n22096), .Z(n22095) );
  XOR U22117 ( .A(n22041), .B(n22055), .Z(n22086) );
  XOR U22118 ( .A(n22097), .B(n22098), .Z(n22055) );
  XNOR U22119 ( .A(n22061), .B(n22099), .Z(n22098) );
  XNOR U22120 ( .A(n22100), .B(n22101), .Z(n22099) );
  XOR U22121 ( .A(n22102), .B(n22103), .Z(n22061) );
  XNOR U22122 ( .A(n21689), .B(n22104), .Z(n22103) );
  XOR U22123 ( .A(n21638), .B(n22105), .Z(n22102) );
  XOR U22124 ( .A(key[297]), .B(n22106), .Z(n22105) );
  XOR U22125 ( .A(n21636), .B(n22107), .Z(n22097) );
  XNOR U22126 ( .A(key[299]), .B(n22108), .Z(n22107) );
  XOR U22127 ( .A(n22109), .B(n22110), .Z(n22041) );
  XOR U22128 ( .A(n22111), .B(n22112), .Z(n22110) );
  XOR U22129 ( .A(n21683), .B(n22113), .Z(n22109) );
  XNOR U22130 ( .A(key[296]), .B(n21664), .Z(n22113) );
  XOR U22131 ( .A(n20431), .B(n18383), .Z(n18341) );
  XOR U22132 ( .A(n21957), .B(n21774), .Z(n18383) );
  XNOR U22133 ( .A(n21831), .B(n22114), .Z(n21774) );
  XNOR U22134 ( .A(n22115), .B(n21886), .Z(n22114) );
  XNOR U22135 ( .A(n21951), .B(n21840), .Z(n21948) );
  ANDN U22136 ( .B(n22117), .A(n21951), .Z(n22115) );
  XOR U22137 ( .A(n21889), .B(n22118), .Z(n21831) );
  XNOR U22138 ( .A(n22119), .B(n22120), .Z(n22118) );
  NAND U22139 ( .A(n21956), .B(n22121), .Z(n22120) );
  IV U22140 ( .A(n21884), .Z(n21957) );
  XOR U22141 ( .A(n21889), .B(n22122), .Z(n21884) );
  XOR U22142 ( .A(n22123), .B(n21833), .Z(n22122) );
  OR U22143 ( .A(n22124), .B(n21962), .Z(n21833) );
  XNOR U22144 ( .A(n21836), .B(n21961), .Z(n21962) );
  ANDN U22145 ( .B(n22125), .A(n22126), .Z(n22123) );
  XNOR U22146 ( .A(n22127), .B(n22119), .Z(n21889) );
  OR U22147 ( .A(n21965), .B(n22128), .Z(n22119) );
  XNOR U22148 ( .A(n22129), .B(n21956), .Z(n21965) );
  XOR U22149 ( .A(n21961), .B(n21840), .Z(n21956) );
  XOR U22150 ( .A(n22130), .B(n22131), .Z(n21840) );
  NANDN U22151 ( .A(n22132), .B(n22133), .Z(n22131) );
  IV U22152 ( .A(n22126), .Z(n21961) );
  XNOR U22153 ( .A(n22134), .B(n22135), .Z(n22126) );
  NANDN U22154 ( .A(n22132), .B(n22136), .Z(n22135) );
  ANDN U22155 ( .B(n22129), .A(n22137), .Z(n22127) );
  IV U22156 ( .A(n21968), .Z(n22129) );
  XOR U22157 ( .A(n21951), .B(n21836), .Z(n21968) );
  XNOR U22158 ( .A(n22138), .B(n22134), .Z(n21836) );
  NANDN U22159 ( .A(n22139), .B(n22140), .Z(n22134) );
  XOR U22160 ( .A(n22136), .B(n22141), .Z(n22140) );
  ANDN U22161 ( .B(n22141), .A(n22142), .Z(n22138) );
  XOR U22162 ( .A(n22143), .B(n22130), .Z(n21951) );
  NANDN U22163 ( .A(n22139), .B(n22144), .Z(n22130) );
  XOR U22164 ( .A(n22145), .B(n22133), .Z(n22144) );
  XNOR U22165 ( .A(n22146), .B(n22147), .Z(n22132) );
  XOR U22166 ( .A(n22148), .B(n22149), .Z(n22147) );
  XNOR U22167 ( .A(n22150), .B(n22151), .Z(n22146) );
  XNOR U22168 ( .A(n22152), .B(n22153), .Z(n22151) );
  ANDN U22169 ( .B(n22145), .A(n22149), .Z(n22152) );
  ANDN U22170 ( .B(n22145), .A(n22142), .Z(n22143) );
  XNOR U22171 ( .A(n22148), .B(n22154), .Z(n22142) );
  XOR U22172 ( .A(n22155), .B(n22153), .Z(n22154) );
  NAND U22173 ( .A(n22156), .B(n22157), .Z(n22153) );
  XNOR U22174 ( .A(n22150), .B(n22133), .Z(n22157) );
  IV U22175 ( .A(n22145), .Z(n22150) );
  XNOR U22176 ( .A(n22136), .B(n22149), .Z(n22156) );
  IV U22177 ( .A(n22141), .Z(n22149) );
  XOR U22178 ( .A(n22158), .B(n22159), .Z(n22141) );
  XNOR U22179 ( .A(n22160), .B(n22161), .Z(n22159) );
  XNOR U22180 ( .A(n22162), .B(n22163), .Z(n22158) );
  ANDN U22181 ( .B(n22117), .A(n21950), .Z(n22162) );
  AND U22182 ( .A(n22133), .B(n22136), .Z(n22155) );
  XNOR U22183 ( .A(n22133), .B(n22136), .Z(n22148) );
  XNOR U22184 ( .A(n22164), .B(n22165), .Z(n22136) );
  XNOR U22185 ( .A(n22166), .B(n22161), .Z(n22165) );
  XOR U22186 ( .A(n22167), .B(n22168), .Z(n22164) );
  XNOR U22187 ( .A(n22169), .B(n22163), .Z(n22168) );
  OR U22188 ( .A(n21949), .B(n22116), .Z(n22163) );
  XNOR U22189 ( .A(n22117), .B(n22170), .Z(n22116) );
  XNOR U22190 ( .A(n21950), .B(n21841), .Z(n21949) );
  ANDN U22191 ( .B(n22171), .A(n21888), .Z(n22169) );
  XNOR U22192 ( .A(n22172), .B(n22173), .Z(n22133) );
  XNOR U22193 ( .A(n22161), .B(n22174), .Z(n22173) );
  XOR U22194 ( .A(n21870), .B(n22167), .Z(n22174) );
  XNOR U22195 ( .A(n22117), .B(n21950), .Z(n22161) );
  XNOR U22196 ( .A(n22175), .B(n22176), .Z(n22172) );
  XNOR U22197 ( .A(n22177), .B(n22178), .Z(n22176) );
  ANDN U22198 ( .B(n22125), .A(n21960), .Z(n22177) );
  XNOR U22199 ( .A(n22179), .B(n22180), .Z(n22145) );
  XNOR U22200 ( .A(n22166), .B(n22181), .Z(n22180) );
  XNOR U22201 ( .A(n21960), .B(n22160), .Z(n22181) );
  XOR U22202 ( .A(n22167), .B(n22182), .Z(n22160) );
  XNOR U22203 ( .A(n22183), .B(n22184), .Z(n22182) );
  NAND U22204 ( .A(n22121), .B(n21955), .Z(n22184) );
  XNOR U22205 ( .A(n22185), .B(n22183), .Z(n22167) );
  NANDN U22206 ( .A(n22128), .B(n21966), .Z(n22183) );
  XOR U22207 ( .A(n21967), .B(n21955), .Z(n21966) );
  XNOR U22208 ( .A(n22186), .B(n21841), .Z(n21955) );
  XOR U22209 ( .A(n22137), .B(n22121), .Z(n22128) );
  XOR U22210 ( .A(n22125), .B(n22170), .Z(n22121) );
  ANDN U22211 ( .B(n21967), .A(n22137), .Z(n22185) );
  XNOR U22212 ( .A(n22175), .B(n22117), .Z(n22137) );
  XNOR U22213 ( .A(n22187), .B(n22188), .Z(n22117) );
  XNOR U22214 ( .A(n22189), .B(n22190), .Z(n22188) );
  XOR U22215 ( .A(n22191), .B(n22192), .Z(n21967) );
  XOR U22216 ( .A(n22170), .B(n22171), .Z(n22166) );
  IV U22217 ( .A(n21841), .Z(n22171) );
  XOR U22218 ( .A(n22193), .B(n22194), .Z(n21841) );
  XNOR U22219 ( .A(n22195), .B(n22190), .Z(n22194) );
  IV U22220 ( .A(n21888), .Z(n22170) );
  XOR U22221 ( .A(n22190), .B(n22196), .Z(n21888) );
  XNOR U22222 ( .A(n22125), .B(n22197), .Z(n22179) );
  XNOR U22223 ( .A(n22198), .B(n22178), .Z(n22197) );
  OR U22224 ( .A(n21963), .B(n22124), .Z(n22178) );
  XNOR U22225 ( .A(n22175), .B(n22125), .Z(n22124) );
  XOR U22226 ( .A(n21870), .B(n22186), .Z(n21963) );
  IV U22227 ( .A(n21960), .Z(n22186) );
  XOR U22228 ( .A(n22192), .B(n22199), .Z(n21960) );
  XNOR U22229 ( .A(n22195), .B(n22187), .Z(n22199) );
  XOR U22230 ( .A(n22200), .B(n22201), .Z(n22187) );
  XOR U22231 ( .A(n21233), .B(n21230), .Z(n22201) );
  XNOR U22232 ( .A(key[338]), .B(n22202), .Z(n22200) );
  IV U22233 ( .A(n21950), .Z(n22192) );
  XOR U22234 ( .A(n22193), .B(n22203), .Z(n21950) );
  XOR U22235 ( .A(n22190), .B(n22204), .Z(n22203) );
  ANDN U22236 ( .B(n22191), .A(n21835), .Z(n22198) );
  IV U22237 ( .A(n21870), .Z(n22191) );
  XOR U22238 ( .A(n22193), .B(n22205), .Z(n21870) );
  XOR U22239 ( .A(n22190), .B(n22206), .Z(n22205) );
  XOR U22240 ( .A(n22207), .B(n22208), .Z(n22190) );
  XOR U22241 ( .A(n22209), .B(n21835), .Z(n22208) );
  IV U22242 ( .A(n22175), .Z(n21835) );
  XNOR U22243 ( .A(n22210), .B(n22211), .Z(n22207) );
  XNOR U22244 ( .A(key[342]), .B(n22212), .Z(n22211) );
  IV U22245 ( .A(n22196), .Z(n22193) );
  XOR U22246 ( .A(n22213), .B(n22214), .Z(n22196) );
  XOR U22247 ( .A(n22215), .B(n22216), .Z(n22214) );
  XNOR U22248 ( .A(key[341]), .B(n22217), .Z(n22213) );
  XOR U22249 ( .A(n22218), .B(n22219), .Z(n22125) );
  XNOR U22250 ( .A(n22206), .B(n22204), .Z(n22219) );
  XNOR U22251 ( .A(n22220), .B(n22221), .Z(n22204) );
  XNOR U22252 ( .A(n22222), .B(n22223), .Z(n22221) );
  XNOR U22253 ( .A(key[343]), .B(n22224), .Z(n22220) );
  XNOR U22254 ( .A(n22225), .B(n22226), .Z(n22206) );
  XNOR U22255 ( .A(n22227), .B(n22228), .Z(n22226) );
  XNOR U22256 ( .A(n22229), .B(n22230), .Z(n22225) );
  XNOR U22257 ( .A(key[340]), .B(n22231), .Z(n22230) );
  XOR U22258 ( .A(n22175), .B(n22189), .Z(n22218) );
  XOR U22259 ( .A(n22232), .B(n22233), .Z(n22189) );
  XNOR U22260 ( .A(n22195), .B(n22234), .Z(n22233) );
  XNOR U22261 ( .A(n22235), .B(n22236), .Z(n22234) );
  XOR U22262 ( .A(n22237), .B(n22238), .Z(n22195) );
  XNOR U22263 ( .A(n21241), .B(n21195), .Z(n22238) );
  XNOR U22264 ( .A(key[337]), .B(n22239), .Z(n22237) );
  XNOR U22265 ( .A(n22240), .B(n22241), .Z(n22232) );
  XNOR U22266 ( .A(key[339]), .B(n21196), .Z(n22241) );
  IV U22267 ( .A(n22242), .Z(n21196) );
  XOR U22268 ( .A(n22243), .B(n22244), .Z(n22175) );
  XNOR U22269 ( .A(n22245), .B(n21234), .Z(n22244) );
  XNOR U22270 ( .A(key[336]), .B(n22246), .Z(n22243) );
  XNOR U22271 ( .A(n21913), .B(n21844), .Z(n20431) );
  XNOR U22272 ( .A(n21971), .B(n22247), .Z(n21844) );
  XOR U22273 ( .A(n22248), .B(n22249), .Z(n22247) );
  ANDN U22274 ( .B(n22250), .A(n21923), .Z(n22248) );
  XNOR U22275 ( .A(n22251), .B(n22252), .Z(n21971) );
  XNOR U22276 ( .A(n22253), .B(n22254), .Z(n22252) );
  NAND U22277 ( .A(n22255), .B(n22256), .Z(n22254) );
  XNOR U22278 ( .A(key[480]), .B(n19552), .Z(n21978) );
  XOR U22279 ( .A(n18368), .B(n18385), .Z(n19552) );
  XNOR U22280 ( .A(n21909), .B(n22257), .Z(n18385) );
  XNOR U22281 ( .A(n21916), .B(n21912), .Z(n22257) );
  XOR U22282 ( .A(n22251), .B(n22258), .Z(n21912) );
  XNOR U22283 ( .A(n22249), .B(n22259), .Z(n22258) );
  NANDN U22284 ( .A(n22260), .B(n21850), .Z(n22259) );
  XNOR U22285 ( .A(n21923), .B(n21850), .Z(n21920) );
  XNOR U22286 ( .A(n21913), .B(n21911), .Z(n21916) );
  XNOR U22287 ( .A(n22262), .B(n22263), .Z(n21911) );
  XNOR U22288 ( .A(n22264), .B(n22265), .Z(n22263) );
  NANDN U22289 ( .A(n22266), .B(n22267), .Z(n22265) );
  XOR U22290 ( .A(n22251), .B(n22268), .Z(n21913) );
  XOR U22291 ( .A(n22269), .B(n21973), .Z(n22268) );
  OR U22292 ( .A(n22270), .B(n22271), .Z(n21973) );
  ANDN U22293 ( .B(n22272), .A(n22273), .Z(n22269) );
  XOR U22294 ( .A(n22274), .B(n22253), .Z(n22251) );
  OR U22295 ( .A(n22275), .B(n22276), .Z(n22253) );
  ANDN U22296 ( .B(n22277), .A(n22278), .Z(n22274) );
  XOR U22297 ( .A(n21917), .B(n22279), .Z(n21909) );
  XNOR U22298 ( .A(n22264), .B(n22280), .Z(n22279) );
  NANDN U22299 ( .A(n22281), .B(n21976), .Z(n22280) );
  OR U22300 ( .A(n22270), .B(n22282), .Z(n22264) );
  XNOR U22301 ( .A(n21976), .B(n22267), .Z(n22270) );
  XOR U22302 ( .A(n22262), .B(n22283), .Z(n21917) );
  XNOR U22303 ( .A(n22284), .B(n22285), .Z(n22283) );
  NAND U22304 ( .A(n22286), .B(n22255), .Z(n22285) );
  IV U22305 ( .A(n21846), .Z(n22262) );
  XNOR U22306 ( .A(n22287), .B(n22284), .Z(n21846) );
  NANDN U22307 ( .A(n22275), .B(n22288), .Z(n22284) );
  XNOR U22308 ( .A(n22277), .B(n22255), .Z(n22275) );
  XOR U22309 ( .A(n22267), .B(n21850), .Z(n22255) );
  XOR U22310 ( .A(n22289), .B(n22290), .Z(n21850) );
  NANDN U22311 ( .A(n22291), .B(n22292), .Z(n22290) );
  IV U22312 ( .A(n22273), .Z(n22267) );
  XNOR U22313 ( .A(n22293), .B(n22294), .Z(n22273) );
  NANDN U22314 ( .A(n22291), .B(n22295), .Z(n22294) );
  IV U22315 ( .A(n22296), .Z(n22277) );
  ANDN U22316 ( .B(n22297), .A(n22296), .Z(n22287) );
  XOR U22317 ( .A(n21923), .B(n21976), .Z(n22296) );
  XNOR U22318 ( .A(n22298), .B(n22293), .Z(n21976) );
  NANDN U22319 ( .A(n22299), .B(n22300), .Z(n22293) );
  XOR U22320 ( .A(n22295), .B(n22301), .Z(n22300) );
  ANDN U22321 ( .B(n22301), .A(n22302), .Z(n22298) );
  XOR U22322 ( .A(n22303), .B(n22289), .Z(n21923) );
  NANDN U22323 ( .A(n22299), .B(n22304), .Z(n22289) );
  XOR U22324 ( .A(n22305), .B(n22292), .Z(n22304) );
  XNOR U22325 ( .A(n22306), .B(n22307), .Z(n22291) );
  XOR U22326 ( .A(n22308), .B(n22309), .Z(n22307) );
  XNOR U22327 ( .A(n22310), .B(n22311), .Z(n22306) );
  XNOR U22328 ( .A(n22312), .B(n22313), .Z(n22311) );
  ANDN U22329 ( .B(n22305), .A(n22309), .Z(n22312) );
  ANDN U22330 ( .B(n22305), .A(n22302), .Z(n22303) );
  XNOR U22331 ( .A(n22308), .B(n22314), .Z(n22302) );
  XOR U22332 ( .A(n22315), .B(n22313), .Z(n22314) );
  NAND U22333 ( .A(n22316), .B(n22317), .Z(n22313) );
  XNOR U22334 ( .A(n22310), .B(n22292), .Z(n22317) );
  IV U22335 ( .A(n22305), .Z(n22310) );
  XNOR U22336 ( .A(n22295), .B(n22309), .Z(n22316) );
  IV U22337 ( .A(n22301), .Z(n22309) );
  XOR U22338 ( .A(n22318), .B(n22319), .Z(n22301) );
  XNOR U22339 ( .A(n22320), .B(n22321), .Z(n22319) );
  XNOR U22340 ( .A(n22322), .B(n22323), .Z(n22318) );
  ANDN U22341 ( .B(n22250), .A(n21922), .Z(n22322) );
  AND U22342 ( .A(n22292), .B(n22295), .Z(n22315) );
  XNOR U22343 ( .A(n22292), .B(n22295), .Z(n22308) );
  XNOR U22344 ( .A(n22324), .B(n22325), .Z(n22295) );
  XNOR U22345 ( .A(n22326), .B(n22321), .Z(n22325) );
  XOR U22346 ( .A(n22327), .B(n22328), .Z(n22324) );
  XNOR U22347 ( .A(n22329), .B(n22323), .Z(n22328) );
  OR U22348 ( .A(n21921), .B(n22261), .Z(n22323) );
  XNOR U22349 ( .A(n22250), .B(n22330), .Z(n22261) );
  XNOR U22350 ( .A(n21922), .B(n21851), .Z(n21921) );
  ANDN U22351 ( .B(n22331), .A(n22260), .Z(n22329) );
  XNOR U22352 ( .A(n22332), .B(n22333), .Z(n22292) );
  XNOR U22353 ( .A(n22321), .B(n22334), .Z(n22333) );
  XOR U22354 ( .A(n22281), .B(n22327), .Z(n22334) );
  XNOR U22355 ( .A(n22250), .B(n21922), .Z(n22321) );
  XNOR U22356 ( .A(n22335), .B(n22336), .Z(n22332) );
  XNOR U22357 ( .A(n22337), .B(n22338), .Z(n22336) );
  ANDN U22358 ( .B(n22272), .A(n22266), .Z(n22337) );
  XNOR U22359 ( .A(n22339), .B(n22340), .Z(n22305) );
  XNOR U22360 ( .A(n22326), .B(n22341), .Z(n22340) );
  XNOR U22361 ( .A(n22266), .B(n22320), .Z(n22341) );
  XOR U22362 ( .A(n22327), .B(n22342), .Z(n22320) );
  XNOR U22363 ( .A(n22343), .B(n22344), .Z(n22342) );
  NAND U22364 ( .A(n22256), .B(n22286), .Z(n22344) );
  XNOR U22365 ( .A(n22345), .B(n22343), .Z(n22327) );
  NANDN U22366 ( .A(n22276), .B(n22288), .Z(n22343) );
  XOR U22367 ( .A(n22297), .B(n22286), .Z(n22288) );
  XNOR U22368 ( .A(n22346), .B(n21851), .Z(n22286) );
  XOR U22369 ( .A(n22278), .B(n22256), .Z(n22276) );
  XOR U22370 ( .A(n22272), .B(n22330), .Z(n22256) );
  ANDN U22371 ( .B(n22297), .A(n22278), .Z(n22345) );
  XNOR U22372 ( .A(n22335), .B(n22250), .Z(n22278) );
  XNOR U22373 ( .A(n22347), .B(n22348), .Z(n22250) );
  XNOR U22374 ( .A(n22349), .B(n22350), .Z(n22348) );
  XOR U22375 ( .A(n22330), .B(n22331), .Z(n22326) );
  IV U22376 ( .A(n21851), .Z(n22331) );
  XOR U22377 ( .A(n22351), .B(n22352), .Z(n21851) );
  XNOR U22378 ( .A(n22353), .B(n22350), .Z(n22352) );
  IV U22379 ( .A(n22260), .Z(n22330) );
  XOR U22380 ( .A(n22350), .B(n22354), .Z(n22260) );
  XNOR U22381 ( .A(n22272), .B(n22355), .Z(n22339) );
  XNOR U22382 ( .A(n22356), .B(n22338), .Z(n22355) );
  OR U22383 ( .A(n22282), .B(n22271), .Z(n22338) );
  XNOR U22384 ( .A(n22335), .B(n22272), .Z(n22271) );
  XOR U22385 ( .A(n22281), .B(n22346), .Z(n22282) );
  IV U22386 ( .A(n22266), .Z(n22346) );
  XOR U22387 ( .A(n22357), .B(n22358), .Z(n22266) );
  XNOR U22388 ( .A(n22353), .B(n22347), .Z(n22358) );
  XOR U22389 ( .A(n22359), .B(n22360), .Z(n22347) );
  XNOR U22390 ( .A(n21384), .B(n21388), .Z(n22360) );
  XNOR U22391 ( .A(n22361), .B(n22362), .Z(n22359) );
  XOR U22392 ( .A(key[378]), .B(n22363), .Z(n22362) );
  ANDN U22393 ( .B(n22364), .A(n21975), .Z(n22356) );
  XOR U22394 ( .A(n22365), .B(n22366), .Z(n22272) );
  XNOR U22395 ( .A(n22367), .B(n22368), .Z(n22366) );
  XOR U22396 ( .A(n22335), .B(n22349), .Z(n22365) );
  XOR U22397 ( .A(n22369), .B(n22370), .Z(n22349) );
  XNOR U22398 ( .A(n22353), .B(n22371), .Z(n22370) );
  XNOR U22399 ( .A(n22372), .B(n22373), .Z(n22371) );
  XOR U22400 ( .A(n22374), .B(n22375), .Z(n22353) );
  XNOR U22401 ( .A(n21372), .B(n22376), .Z(n22375) );
  XOR U22402 ( .A(n21399), .B(n22377), .Z(n22374) );
  XOR U22403 ( .A(key[377]), .B(n22378), .Z(n22377) );
  XOR U22404 ( .A(n21397), .B(n22379), .Z(n22369) );
  XNOR U22405 ( .A(key[379]), .B(n22380), .Z(n22379) );
  XOR U22406 ( .A(n22364), .B(n22357), .Z(n22297) );
  IV U22407 ( .A(n21922), .Z(n22357) );
  XOR U22408 ( .A(n22351), .B(n22381), .Z(n21922) );
  XOR U22409 ( .A(n22350), .B(n22368), .Z(n22381) );
  XNOR U22410 ( .A(n22382), .B(n22383), .Z(n22368) );
  XNOR U22411 ( .A(n21373), .B(n22384), .Z(n22383) );
  XNOR U22412 ( .A(key[383]), .B(n22385), .Z(n22382) );
  IV U22413 ( .A(n22281), .Z(n22364) );
  XOR U22414 ( .A(n22351), .B(n22386), .Z(n22281) );
  XOR U22415 ( .A(n22350), .B(n22367), .Z(n22386) );
  XNOR U22416 ( .A(n22387), .B(n22388), .Z(n22367) );
  XNOR U22417 ( .A(n22389), .B(n22390), .Z(n22387) );
  XNOR U22418 ( .A(key[380]), .B(n22391), .Z(n22390) );
  XOR U22419 ( .A(n22392), .B(n22393), .Z(n22350) );
  XNOR U22420 ( .A(n22394), .B(n21975), .Z(n22393) );
  IV U22421 ( .A(n22335), .Z(n21975) );
  XOR U22422 ( .A(n22395), .B(n22396), .Z(n22335) );
  XOR U22423 ( .A(n22397), .B(n22398), .Z(n22396) );
  XOR U22424 ( .A(n21391), .B(n22399), .Z(n22395) );
  XNOR U22425 ( .A(key[376]), .B(n21358), .Z(n22399) );
  XOR U22426 ( .A(n21363), .B(n22400), .Z(n22392) );
  XNOR U22427 ( .A(key[382]), .B(n22401), .Z(n22400) );
  IV U22428 ( .A(n22354), .Z(n22351) );
  XOR U22429 ( .A(n22402), .B(n22403), .Z(n22354) );
  XOR U22430 ( .A(n22404), .B(n22405), .Z(n22403) );
  XOR U22431 ( .A(n21377), .B(n22406), .Z(n22402) );
  XNOR U22432 ( .A(key[381]), .B(n22407), .Z(n22406) );
  IV U22433 ( .A(n19561), .Z(n18368) );
  XOR U22434 ( .A(n22408), .B(n22409), .Z(n19561) );
  XOR U22435 ( .A(n22410), .B(n21906), .Z(n22409) );
  XOR U22436 ( .A(n19558), .B(n18339), .Z(n19543) );
  XNOR U22437 ( .A(n22411), .B(n22412), .Z(n18339) );
  XNOR U22438 ( .A(n21812), .B(n21780), .Z(n22412) );
  XNOR U22439 ( .A(n22413), .B(n22414), .Z(n21780) );
  XNOR U22440 ( .A(n22415), .B(n22416), .Z(n22414) );
  NANDN U22441 ( .A(n22417), .B(n22418), .Z(n22416) );
  IV U22442 ( .A(n22408), .Z(n21812) );
  XNOR U22443 ( .A(n21862), .B(n21898), .Z(n22408) );
  XNOR U22444 ( .A(n21781), .B(n22419), .Z(n21898) );
  XNOR U22445 ( .A(n22420), .B(n22421), .Z(n22419) );
  NANDN U22446 ( .A(n22422), .B(n22423), .Z(n22421) );
  XNOR U22447 ( .A(n22410), .B(n21906), .Z(n22411) );
  XNOR U22448 ( .A(n22420), .B(n22425), .Z(n22424) );
  NANDN U22449 ( .A(n22426), .B(n22418), .Z(n22425) );
  OR U22450 ( .A(n22427), .B(n22428), .Z(n22420) );
  XNOR U22451 ( .A(n21781), .B(n22429), .Z(n21899) );
  XNOR U22452 ( .A(n22430), .B(n22431), .Z(n22429) );
  NAND U22453 ( .A(n22432), .B(n22433), .Z(n22431) );
  XOR U22454 ( .A(n22434), .B(n22430), .Z(n21781) );
  NANDN U22455 ( .A(n22435), .B(n22436), .Z(n22430) );
  ANDN U22456 ( .B(n22437), .A(n22438), .Z(n22434) );
  IV U22457 ( .A(n21861), .Z(n22410) );
  XOR U22458 ( .A(n22440), .B(n22441), .Z(n22439) );
  NANDN U22459 ( .A(n22442), .B(n21785), .Z(n22441) );
  XOR U22460 ( .A(n21862), .B(n21779), .Z(n19558) );
  XNOR U22461 ( .A(n22413), .B(n22444), .Z(n21779) );
  XNOR U22462 ( .A(n22445), .B(n22440), .Z(n22444) );
  XNOR U22463 ( .A(n21905), .B(n21785), .Z(n21902) );
  ANDN U22464 ( .B(n22447), .A(n21905), .Z(n22445) );
  XOR U22465 ( .A(n22443), .B(n22448), .Z(n22413) );
  XNOR U22466 ( .A(n22449), .B(n22450), .Z(n22448) );
  NAND U22467 ( .A(n22433), .B(n22451), .Z(n22450) );
  XNOR U22468 ( .A(n22443), .B(n22452), .Z(n21862) );
  XOR U22469 ( .A(n22453), .B(n22415), .Z(n22452) );
  OR U22470 ( .A(n22454), .B(n22427), .Z(n22415) );
  XNOR U22471 ( .A(n22418), .B(n22423), .Z(n22427) );
  ANDN U22472 ( .B(n22455), .A(n22456), .Z(n22453) );
  XNOR U22473 ( .A(n22457), .B(n22449), .Z(n22443) );
  OR U22474 ( .A(n22435), .B(n22458), .Z(n22449) );
  XNOR U22475 ( .A(n22459), .B(n22433), .Z(n22435) );
  XOR U22476 ( .A(n22423), .B(n21785), .Z(n22433) );
  XOR U22477 ( .A(n22460), .B(n22461), .Z(n21785) );
  NANDN U22478 ( .A(n22462), .B(n22463), .Z(n22461) );
  IV U22479 ( .A(n22456), .Z(n22423) );
  XNOR U22480 ( .A(n22464), .B(n22465), .Z(n22456) );
  NANDN U22481 ( .A(n22462), .B(n22466), .Z(n22465) );
  ANDN U22482 ( .B(n22459), .A(n22467), .Z(n22457) );
  IV U22483 ( .A(n22438), .Z(n22459) );
  XOR U22484 ( .A(n21905), .B(n22418), .Z(n22438) );
  XNOR U22485 ( .A(n22468), .B(n22464), .Z(n22418) );
  NANDN U22486 ( .A(n22469), .B(n22470), .Z(n22464) );
  XOR U22487 ( .A(n22466), .B(n22471), .Z(n22470) );
  ANDN U22488 ( .B(n22471), .A(n22472), .Z(n22468) );
  XOR U22489 ( .A(n22473), .B(n22460), .Z(n21905) );
  NANDN U22490 ( .A(n22469), .B(n22474), .Z(n22460) );
  XOR U22491 ( .A(n22475), .B(n22463), .Z(n22474) );
  XNOR U22492 ( .A(n22476), .B(n22477), .Z(n22462) );
  XOR U22493 ( .A(n22478), .B(n22479), .Z(n22477) );
  XNOR U22494 ( .A(n22480), .B(n22481), .Z(n22476) );
  XNOR U22495 ( .A(n22482), .B(n22483), .Z(n22481) );
  ANDN U22496 ( .B(n22475), .A(n22479), .Z(n22482) );
  ANDN U22497 ( .B(n22475), .A(n22472), .Z(n22473) );
  XNOR U22498 ( .A(n22478), .B(n22484), .Z(n22472) );
  XOR U22499 ( .A(n22485), .B(n22483), .Z(n22484) );
  NAND U22500 ( .A(n22486), .B(n22487), .Z(n22483) );
  XNOR U22501 ( .A(n22480), .B(n22463), .Z(n22487) );
  IV U22502 ( .A(n22475), .Z(n22480) );
  XNOR U22503 ( .A(n22466), .B(n22479), .Z(n22486) );
  IV U22504 ( .A(n22471), .Z(n22479) );
  XOR U22505 ( .A(n22488), .B(n22489), .Z(n22471) );
  XNOR U22506 ( .A(n22490), .B(n22491), .Z(n22489) );
  XNOR U22507 ( .A(n22492), .B(n22493), .Z(n22488) );
  ANDN U22508 ( .B(n22447), .A(n21904), .Z(n22492) );
  AND U22509 ( .A(n22463), .B(n22466), .Z(n22485) );
  XNOR U22510 ( .A(n22463), .B(n22466), .Z(n22478) );
  XNOR U22511 ( .A(n22494), .B(n22495), .Z(n22466) );
  XNOR U22512 ( .A(n22496), .B(n22491), .Z(n22495) );
  XOR U22513 ( .A(n22497), .B(n22498), .Z(n22494) );
  XNOR U22514 ( .A(n22499), .B(n22493), .Z(n22498) );
  OR U22515 ( .A(n21903), .B(n22446), .Z(n22493) );
  XNOR U22516 ( .A(n22447), .B(n22500), .Z(n22446) );
  XNOR U22517 ( .A(n21904), .B(n21786), .Z(n21903) );
  ANDN U22518 ( .B(n22501), .A(n22442), .Z(n22499) );
  XNOR U22519 ( .A(n22502), .B(n22503), .Z(n22463) );
  XNOR U22520 ( .A(n22491), .B(n22504), .Z(n22503) );
  XOR U22521 ( .A(n22426), .B(n22497), .Z(n22504) );
  XNOR U22522 ( .A(n22447), .B(n21904), .Z(n22491) );
  XNOR U22523 ( .A(n22505), .B(n22506), .Z(n22502) );
  XNOR U22524 ( .A(n22507), .B(n22508), .Z(n22506) );
  ANDN U22525 ( .B(n22455), .A(n22422), .Z(n22507) );
  XNOR U22526 ( .A(n22509), .B(n22510), .Z(n22475) );
  XNOR U22527 ( .A(n22496), .B(n22511), .Z(n22510) );
  XNOR U22528 ( .A(n22422), .B(n22490), .Z(n22511) );
  XOR U22529 ( .A(n22497), .B(n22512), .Z(n22490) );
  XNOR U22530 ( .A(n22513), .B(n22514), .Z(n22512) );
  NAND U22531 ( .A(n22451), .B(n22432), .Z(n22514) );
  XNOR U22532 ( .A(n22515), .B(n22513), .Z(n22497) );
  NANDN U22533 ( .A(n22458), .B(n22436), .Z(n22513) );
  XOR U22534 ( .A(n22437), .B(n22432), .Z(n22436) );
  XNOR U22535 ( .A(n22516), .B(n21786), .Z(n22432) );
  XOR U22536 ( .A(n22467), .B(n22451), .Z(n22458) );
  XOR U22537 ( .A(n22455), .B(n22500), .Z(n22451) );
  ANDN U22538 ( .B(n22437), .A(n22467), .Z(n22515) );
  XNOR U22539 ( .A(n22505), .B(n22447), .Z(n22467) );
  XNOR U22540 ( .A(n22517), .B(n22518), .Z(n22447) );
  XNOR U22541 ( .A(n22519), .B(n22520), .Z(n22518) );
  XOR U22542 ( .A(n22521), .B(n22522), .Z(n22437) );
  XOR U22543 ( .A(n22500), .B(n22501), .Z(n22496) );
  IV U22544 ( .A(n21786), .Z(n22501) );
  XOR U22545 ( .A(n22523), .B(n22524), .Z(n21786) );
  XNOR U22546 ( .A(n22525), .B(n22520), .Z(n22524) );
  IV U22547 ( .A(n22442), .Z(n22500) );
  XOR U22548 ( .A(n22520), .B(n22526), .Z(n22442) );
  XNOR U22549 ( .A(n22455), .B(n22527), .Z(n22509) );
  XNOR U22550 ( .A(n22528), .B(n22508), .Z(n22527) );
  OR U22551 ( .A(n22428), .B(n22454), .Z(n22508) );
  XNOR U22552 ( .A(n22505), .B(n22455), .Z(n22454) );
  XOR U22553 ( .A(n22426), .B(n22516), .Z(n22428) );
  IV U22554 ( .A(n22422), .Z(n22516) );
  XOR U22555 ( .A(n22522), .B(n22529), .Z(n22422) );
  XNOR U22556 ( .A(n22525), .B(n22517), .Z(n22529) );
  XOR U22557 ( .A(n22530), .B(n22531), .Z(n22517) );
  XOR U22558 ( .A(n21511), .B(n21508), .Z(n22531) );
  XNOR U22559 ( .A(key[258]), .B(n22532), .Z(n22530) );
  IV U22560 ( .A(n21904), .Z(n22522) );
  XOR U22561 ( .A(n22523), .B(n22533), .Z(n21904) );
  XOR U22562 ( .A(n22520), .B(n22534), .Z(n22533) );
  ANDN U22563 ( .B(n22521), .A(n22417), .Z(n22528) );
  IV U22564 ( .A(n22426), .Z(n22521) );
  XOR U22565 ( .A(n22523), .B(n22535), .Z(n22426) );
  XOR U22566 ( .A(n22520), .B(n22536), .Z(n22535) );
  XOR U22567 ( .A(n22537), .B(n22538), .Z(n22520) );
  XOR U22568 ( .A(n22539), .B(n22417), .Z(n22538) );
  IV U22569 ( .A(n22505), .Z(n22417) );
  XNOR U22570 ( .A(n22540), .B(n22541), .Z(n22537) );
  XNOR U22571 ( .A(key[262]), .B(n22542), .Z(n22541) );
  IV U22572 ( .A(n22526), .Z(n22523) );
  XOR U22573 ( .A(n22543), .B(n22544), .Z(n22526) );
  XOR U22574 ( .A(n22545), .B(n22546), .Z(n22544) );
  XNOR U22575 ( .A(key[261]), .B(n22547), .Z(n22543) );
  XOR U22576 ( .A(n22548), .B(n22549), .Z(n22455) );
  XNOR U22577 ( .A(n22536), .B(n22534), .Z(n22549) );
  XNOR U22578 ( .A(n22550), .B(n22551), .Z(n22534) );
  XNOR U22579 ( .A(n22552), .B(n22553), .Z(n22551) );
  XOR U22580 ( .A(key[263]), .B(n22554), .Z(n22550) );
  XNOR U22581 ( .A(n22555), .B(n22556), .Z(n22536) );
  XNOR U22582 ( .A(n22557), .B(n22558), .Z(n22556) );
  XNOR U22583 ( .A(n22559), .B(n22560), .Z(n22555) );
  XNOR U22584 ( .A(key[260]), .B(n22561), .Z(n22560) );
  XOR U22585 ( .A(n22505), .B(n22519), .Z(n22548) );
  XOR U22586 ( .A(n22562), .B(n22563), .Z(n22519) );
  XNOR U22587 ( .A(n22525), .B(n22564), .Z(n22563) );
  XNOR U22588 ( .A(n22565), .B(n22566), .Z(n22564) );
  XOR U22589 ( .A(n22567), .B(n22568), .Z(n22525) );
  XOR U22590 ( .A(n21540), .B(n21520), .Z(n22568) );
  XNOR U22591 ( .A(key[257]), .B(n22569), .Z(n22567) );
  XNOR U22592 ( .A(n21521), .B(n22570), .Z(n22562) );
  XNOR U22593 ( .A(key[259]), .B(n22571), .Z(n22570) );
  IV U22594 ( .A(n22572), .Z(n21521) );
  XOR U22595 ( .A(n22573), .B(n22574), .Z(n22505) );
  XNOR U22596 ( .A(n22575), .B(n22576), .Z(n22574) );
  XNOR U22597 ( .A(key[256]), .B(n22577), .Z(n22573) );
  XOR U22598 ( .A(n20623), .B(n20670), .Z(n15309) );
  XNOR U22599 ( .A(n20629), .B(n22578), .Z(n20670) );
  XNOR U22600 ( .A(n20626), .B(n22579), .Z(n22578) );
  NAND U22601 ( .A(n22580), .B(n20579), .Z(n22579) );
  XOR U22602 ( .A(n20627), .B(n20579), .Z(n20681) );
  XOR U22603 ( .A(n22583), .B(n20572), .Z(n22582) );
  OR U22604 ( .A(n20692), .B(n22584), .Z(n20572) );
  XNOR U22605 ( .A(n20574), .B(n20687), .Z(n20692) );
  NOR U22606 ( .A(n22585), .B(n20687), .Z(n22583) );
  XNOR U22607 ( .A(n22586), .B(n20631), .Z(n20629) );
  OR U22608 ( .A(n20699), .B(n22587), .Z(n20631) );
  XOR U22609 ( .A(n22588), .B(n20633), .Z(n20699) );
  XOR U22610 ( .A(n20687), .B(n20579), .Z(n20633) );
  XOR U22611 ( .A(n22589), .B(n22590), .Z(n20579) );
  NANDN U22612 ( .A(n22591), .B(n22592), .Z(n22590) );
  XNOR U22613 ( .A(n22593), .B(n22594), .Z(n20687) );
  OR U22614 ( .A(n22591), .B(n22595), .Z(n22594) );
  ANDN U22615 ( .B(n22588), .A(n22596), .Z(n22586) );
  IV U22616 ( .A(n20702), .Z(n22588) );
  XOR U22617 ( .A(n20574), .B(n20627), .Z(n20702) );
  XNOR U22618 ( .A(n22597), .B(n22589), .Z(n20627) );
  NANDN U22619 ( .A(n22598), .B(n22599), .Z(n22589) );
  ANDN U22620 ( .B(n22600), .A(n22601), .Z(n22597) );
  NANDN U22621 ( .A(n22598), .B(n22603), .Z(n22593) );
  XOR U22622 ( .A(n22604), .B(n22591), .Z(n22598) );
  XNOR U22623 ( .A(n22605), .B(n22606), .Z(n22591) );
  XOR U22624 ( .A(n22607), .B(n22600), .Z(n22606) );
  XNOR U22625 ( .A(n22608), .B(n22609), .Z(n22605) );
  XNOR U22626 ( .A(n22610), .B(n22611), .Z(n22609) );
  ANDN U22627 ( .B(n22600), .A(n22612), .Z(n22610) );
  IV U22628 ( .A(n22613), .Z(n22600) );
  ANDN U22629 ( .B(n22604), .A(n22612), .Z(n22602) );
  IV U22630 ( .A(n22608), .Z(n22612) );
  IV U22631 ( .A(n22601), .Z(n22604) );
  XNOR U22632 ( .A(n22607), .B(n22614), .Z(n22601) );
  XOR U22633 ( .A(n22615), .B(n22611), .Z(n22614) );
  NAND U22634 ( .A(n22603), .B(n22599), .Z(n22611) );
  XNOR U22635 ( .A(n22592), .B(n22613), .Z(n22599) );
  XOR U22636 ( .A(n22616), .B(n22617), .Z(n22613) );
  XOR U22637 ( .A(n22618), .B(n22619), .Z(n22617) );
  XNOR U22638 ( .A(n20688), .B(n22620), .Z(n22619) );
  XNOR U22639 ( .A(n22621), .B(n22622), .Z(n22616) );
  XNOR U22640 ( .A(n22623), .B(n22624), .Z(n22622) );
  ANDN U22641 ( .B(n22625), .A(n20575), .Z(n22623) );
  XNOR U22642 ( .A(n22608), .B(n22595), .Z(n22603) );
  XOR U22643 ( .A(n22626), .B(n22627), .Z(n22608) );
  XNOR U22644 ( .A(n22628), .B(n22620), .Z(n22627) );
  XOR U22645 ( .A(n22629), .B(n22630), .Z(n22620) );
  XNOR U22646 ( .A(n22631), .B(n22632), .Z(n22630) );
  NAND U22647 ( .A(n20634), .B(n20697), .Z(n22632) );
  XNOR U22648 ( .A(n22633), .B(n22634), .Z(n22626) );
  ANDN U22649 ( .B(n22635), .A(n20628), .Z(n22633) );
  ANDN U22650 ( .B(n22592), .A(n22595), .Z(n22615) );
  XOR U22651 ( .A(n22595), .B(n22592), .Z(n22607) );
  XNOR U22652 ( .A(n22636), .B(n22637), .Z(n22592) );
  XNOR U22653 ( .A(n22629), .B(n22638), .Z(n22637) );
  XOR U22654 ( .A(n22628), .B(n20691), .Z(n22638) );
  XOR U22655 ( .A(n20575), .B(n22639), .Z(n22636) );
  XNOR U22656 ( .A(n22640), .B(n22624), .Z(n22639) );
  OR U22657 ( .A(n20693), .B(n22584), .Z(n22624) );
  XNOR U22658 ( .A(n20575), .B(n22585), .Z(n22584) );
  XOR U22659 ( .A(n20691), .B(n20688), .Z(n20693) );
  ANDN U22660 ( .B(n20688), .A(n22585), .Z(n22640) );
  XOR U22661 ( .A(n22641), .B(n22642), .Z(n22595) );
  XOR U22662 ( .A(n22629), .B(n22618), .Z(n22642) );
  XOR U22663 ( .A(n22580), .B(n20580), .Z(n22618) );
  XOR U22664 ( .A(n22643), .B(n22631), .Z(n22629) );
  NANDN U22665 ( .A(n22587), .B(n20700), .Z(n22631) );
  XOR U22666 ( .A(n20701), .B(n20697), .Z(n20700) );
  XNOR U22667 ( .A(n22635), .B(n22644), .Z(n20688) );
  XNOR U22668 ( .A(n22645), .B(n22646), .Z(n22644) );
  XOR U22669 ( .A(n22596), .B(n20634), .Z(n22587) );
  XNOR U22670 ( .A(n22585), .B(n22580), .Z(n20634) );
  IV U22671 ( .A(n22621), .Z(n22585) );
  XOR U22672 ( .A(n22647), .B(n22648), .Z(n22621) );
  XOR U22673 ( .A(n22649), .B(n22650), .Z(n22648) );
  XNOR U22674 ( .A(n20575), .B(n22651), .Z(n22647) );
  ANDN U22675 ( .B(n20701), .A(n22596), .Z(n22643) );
  XNOR U22676 ( .A(n20575), .B(n20628), .Z(n22596) );
  XOR U22677 ( .A(n22635), .B(n22625), .Z(n20701) );
  IV U22678 ( .A(n20691), .Z(n22625) );
  XOR U22679 ( .A(n22652), .B(n22653), .Z(n20691) );
  XOR U22680 ( .A(n22654), .B(n22650), .Z(n22653) );
  XNOR U22681 ( .A(n22655), .B(n22656), .Z(n22650) );
  XNOR U22682 ( .A(n20287), .B(n19124), .Z(n22656) );
  XOR U22683 ( .A(n20289), .B(n18223), .Z(n19124) );
  XNOR U22684 ( .A(n22657), .B(n18194), .Z(n18223) );
  XNOR U22685 ( .A(n19126), .B(n22659), .Z(n22655) );
  XNOR U22686 ( .A(key[476]), .B(n18225), .Z(n22659) );
  XNOR U22687 ( .A(n18218), .B(n20275), .Z(n18225) );
  XOR U22688 ( .A(n18242), .B(n19143), .Z(n19126) );
  XOR U22689 ( .A(n22660), .B(n22661), .Z(n19143) );
  XNOR U22690 ( .A(n22662), .B(n22663), .Z(n22661) );
  XNOR U22691 ( .A(n22664), .B(n22665), .Z(n22660) );
  XOR U22692 ( .A(n22666), .B(n22667), .Z(n22665) );
  ANDN U22693 ( .B(n22668), .A(n22669), .Z(n22667) );
  IV U22694 ( .A(n20683), .Z(n22635) );
  XOR U22695 ( .A(n22628), .B(n22670), .Z(n22641) );
  XNOR U22696 ( .A(n22671), .B(n22634), .Z(n22670) );
  OR U22697 ( .A(n20682), .B(n22581), .Z(n22634) );
  XNOR U22698 ( .A(n22672), .B(n22580), .Z(n22581) );
  XNOR U22699 ( .A(n20683), .B(n20580), .Z(n20682) );
  ANDN U22700 ( .B(n22580), .A(n20580), .Z(n22671) );
  XOR U22701 ( .A(n22652), .B(n22673), .Z(n20580) );
  XOR U22702 ( .A(n22645), .B(n22674), .Z(n22673) );
  XOR U22703 ( .A(n22654), .B(n22652), .Z(n22580) );
  XNOR U22704 ( .A(n20628), .B(n20683), .Z(n22628) );
  XOR U22705 ( .A(n22652), .B(n22675), .Z(n20683) );
  XNOR U22706 ( .A(n22654), .B(n22649), .Z(n22675) );
  XOR U22707 ( .A(n22676), .B(n22677), .Z(n22649) );
  XOR U22708 ( .A(n19134), .B(n20267), .Z(n22677) );
  XOR U22709 ( .A(n22678), .B(n22679), .Z(n20267) );
  XOR U22710 ( .A(n22680), .B(n22681), .Z(n22679) );
  XOR U22711 ( .A(n22682), .B(n22683), .Z(n22678) );
  XOR U22712 ( .A(n18218), .B(n18242), .Z(n19134) );
  XNOR U22713 ( .A(key[479]), .B(n19119), .Z(n22676) );
  XOR U22714 ( .A(n20282), .B(n20269), .Z(n19119) );
  XNOR U22715 ( .A(n22684), .B(n22685), .Z(n20269) );
  XOR U22716 ( .A(n22686), .B(n22687), .Z(n22685) );
  XNOR U22717 ( .A(n22688), .B(n22689), .Z(n22684) );
  XNOR U22718 ( .A(n22690), .B(n22691), .Z(n22652) );
  XNOR U22719 ( .A(n20276), .B(n19136), .Z(n22691) );
  XOR U22720 ( .A(n22692), .B(n22693), .Z(n19136) );
  XNOR U22721 ( .A(n22694), .B(n22695), .Z(n20276) );
  XNOR U22722 ( .A(n22696), .B(n22681), .Z(n22695) );
  XNOR U22723 ( .A(n22697), .B(n22698), .Z(n22681) );
  XNOR U22724 ( .A(n22699), .B(n22700), .Z(n22698) );
  OR U22725 ( .A(n22701), .B(n22702), .Z(n22700) );
  XNOR U22726 ( .A(n22658), .B(n22703), .Z(n22694) );
  XNOR U22727 ( .A(n22704), .B(n22705), .Z(n22703) );
  ANDN U22728 ( .B(n22706), .A(n22707), .Z(n22704) );
  XNOR U22729 ( .A(n19141), .B(n22708), .Z(n22690) );
  XNOR U22730 ( .A(key[477]), .B(n20272), .Z(n22708) );
  XNOR U22731 ( .A(n20275), .B(n18209), .Z(n19141) );
  XNOR U22732 ( .A(n22709), .B(n22710), .Z(n18209) );
  XNOR U22733 ( .A(n22711), .B(n22687), .Z(n22710) );
  XNOR U22734 ( .A(n22712), .B(n22713), .Z(n22687) );
  XNOR U22735 ( .A(n22714), .B(n22715), .Z(n22713) );
  NANDN U22736 ( .A(n22716), .B(n22717), .Z(n22715) );
  XNOR U22737 ( .A(n22657), .B(n22718), .Z(n22709) );
  XOR U22738 ( .A(n22719), .B(n22720), .Z(n22718) );
  ANDN U22739 ( .B(n22721), .A(n22722), .Z(n22720) );
  XNOR U22740 ( .A(n22723), .B(n22724), .Z(n20275) );
  XNOR U22741 ( .A(n22725), .B(n22726), .Z(n22724) );
  XNOR U22742 ( .A(n22727), .B(n22728), .Z(n22723) );
  XOR U22743 ( .A(n22729), .B(n22730), .Z(n22728) );
  ANDN U22744 ( .B(n22731), .A(n22732), .Z(n22730) );
  IV U22745 ( .A(n22672), .Z(n20628) );
  XNOR U22746 ( .A(n22646), .B(n22733), .Z(n22672) );
  XOR U22747 ( .A(n22651), .B(n22674), .Z(n22733) );
  IV U22748 ( .A(n22654), .Z(n22674) );
  XOR U22749 ( .A(n22734), .B(n22735), .Z(n22654) );
  XNOR U22750 ( .A(n18206), .B(n19138), .Z(n22735) );
  XNOR U22751 ( .A(n18211), .B(n19118), .Z(n19138) );
  XOR U22752 ( .A(n18242), .B(n20283), .Z(n19118) );
  XOR U22753 ( .A(n22736), .B(n22737), .Z(n20283) );
  XNOR U22754 ( .A(n22692), .B(n22663), .Z(n22737) );
  XNOR U22755 ( .A(n22738), .B(n22739), .Z(n22663) );
  XNOR U22756 ( .A(n22740), .B(n22741), .Z(n22739) );
  OR U22757 ( .A(n22742), .B(n22743), .Z(n22741) );
  XOR U22758 ( .A(n20272), .B(n18204), .Z(n18211) );
  XNOR U22759 ( .A(n22744), .B(n22745), .Z(n18204) );
  XOR U22760 ( .A(n22748), .B(n22749), .Z(n20272) );
  XOR U22761 ( .A(n18218), .B(n20282), .Z(n18206) );
  XOR U22762 ( .A(n22750), .B(n22751), .Z(n20282) );
  XOR U22763 ( .A(n22748), .B(n22726), .Z(n22751) );
  XNOR U22764 ( .A(n22752), .B(n22753), .Z(n22726) );
  XNOR U22765 ( .A(n22754), .B(n22755), .Z(n22753) );
  NANDN U22766 ( .A(n22756), .B(n22757), .Z(n22755) );
  XOR U22767 ( .A(n22758), .B(n22759), .Z(n22750) );
  XOR U22768 ( .A(n20270), .B(n22760), .Z(n22734) );
  XOR U22769 ( .A(key[478]), .B(n20575), .Z(n22760) );
  XNOR U22770 ( .A(n22761), .B(n22762), .Z(n20575) );
  XOR U22771 ( .A(n20298), .B(n20296), .Z(n22762) );
  XOR U22772 ( .A(n22764), .B(n22765), .Z(n22763) );
  XNOR U22773 ( .A(n22766), .B(n22767), .Z(n22692) );
  XNOR U22774 ( .A(n18243), .B(n22768), .Z(n22761) );
  XNOR U22775 ( .A(key[472]), .B(n22769), .Z(n22768) );
  XNOR U22776 ( .A(n20286), .B(n20268), .Z(n18243) );
  XOR U22777 ( .A(n22746), .B(n22657), .Z(n20268) );
  XNOR U22778 ( .A(n22712), .B(n22770), .Z(n22657) );
  XNOR U22779 ( .A(n22771), .B(n22772), .Z(n22770) );
  NANDN U22780 ( .A(n22773), .B(n22774), .Z(n22772) );
  XNOR U22781 ( .A(n22775), .B(n22776), .Z(n22712) );
  XNOR U22782 ( .A(n22777), .B(n22778), .Z(n22776) );
  NAND U22783 ( .A(n22779), .B(n22780), .Z(n22778) );
  IV U22784 ( .A(n19120), .Z(n20286) );
  XOR U22785 ( .A(n22781), .B(n22658), .Z(n19120) );
  XNOR U22786 ( .A(n22697), .B(n22782), .Z(n22658) );
  XOR U22787 ( .A(n22783), .B(n22784), .Z(n22782) );
  NOR U22788 ( .A(n22785), .B(n22786), .Z(n22783) );
  XNOR U22789 ( .A(n22787), .B(n22788), .Z(n22697) );
  XNOR U22790 ( .A(n22789), .B(n22790), .Z(n22788) );
  NAND U22791 ( .A(n22791), .B(n22792), .Z(n22790) );
  XOR U22792 ( .A(n22793), .B(n22682), .Z(n20270) );
  XOR U22793 ( .A(n22794), .B(n22795), .Z(n22651) );
  XNOR U22794 ( .A(n20301), .B(n22796), .Z(n22795) );
  XOR U22795 ( .A(n22645), .B(n18196), .Z(n22796) );
  XOR U22796 ( .A(n20300), .B(n18236), .Z(n18196) );
  XNOR U22797 ( .A(n22797), .B(n22798), .Z(n18236) );
  XOR U22798 ( .A(n22799), .B(n22744), .Z(n22798) );
  XNOR U22799 ( .A(n22800), .B(n22801), .Z(n22744) );
  XNOR U22800 ( .A(n22802), .B(n22719), .Z(n22801) );
  NOR U22801 ( .A(n22803), .B(n22804), .Z(n22719) );
  ANDN U22802 ( .B(n22774), .A(n22805), .Z(n22802) );
  XNOR U22803 ( .A(n22747), .B(n22689), .Z(n22797) );
  XOR U22804 ( .A(n22806), .B(n22807), .Z(n22645) );
  XOR U22805 ( .A(n20295), .B(n18241), .Z(n22807) );
  XOR U22806 ( .A(n20298), .B(n18235), .Z(n18241) );
  XOR U22807 ( .A(n22686), .B(n22808), .Z(n18235) );
  XOR U22808 ( .A(n22688), .B(n22689), .Z(n22808) );
  XNOR U22809 ( .A(n22746), .B(n22747), .Z(n22688) );
  XNOR U22810 ( .A(n22711), .B(n22809), .Z(n22747) );
  XNOR U22811 ( .A(n22810), .B(n22811), .Z(n22809) );
  NANDN U22812 ( .A(n22812), .B(n22813), .Z(n22811) );
  IV U22813 ( .A(n22799), .Z(n22686) );
  XOR U22814 ( .A(n22800), .B(n22814), .Z(n22799) );
  XOR U22815 ( .A(n22815), .B(n22810), .Z(n22814) );
  OR U22816 ( .A(n22816), .B(n22817), .Z(n22810) );
  AND U22817 ( .A(n22717), .B(n22818), .Z(n22815) );
  XOR U22818 ( .A(n22711), .B(n22819), .Z(n22800) );
  XNOR U22819 ( .A(n22820), .B(n22821), .Z(n22819) );
  NAND U22820 ( .A(n22822), .B(n22779), .Z(n22821) );
  XOR U22821 ( .A(n22823), .B(n22820), .Z(n22711) );
  NANDN U22822 ( .A(n22824), .B(n22825), .Z(n22820) );
  ANDN U22823 ( .B(n22826), .A(n22827), .Z(n22823) );
  XNOR U22824 ( .A(n22748), .B(n22828), .Z(n20298) );
  XOR U22825 ( .A(n22829), .B(n22759), .Z(n22828) );
  XOR U22826 ( .A(n22830), .B(n22831), .Z(n22748) );
  XNOR U22827 ( .A(n22680), .B(n22832), .Z(n20295) );
  XOR U22828 ( .A(n22682), .B(n22833), .Z(n22832) );
  XNOR U22829 ( .A(n22835), .B(n22836), .Z(n22806) );
  XNOR U22830 ( .A(key[473]), .B(n20260), .Z(n22836) );
  IV U22831 ( .A(n20257), .Z(n20301) );
  XNOR U22832 ( .A(n22837), .B(n22838), .Z(n20257) );
  XNOR U22833 ( .A(n22839), .B(n22840), .Z(n22793) );
  XNOR U22834 ( .A(n22705), .B(n22841), .Z(n22840) );
  OR U22835 ( .A(n22786), .B(n22842), .Z(n22841) );
  NANDN U22836 ( .A(n22843), .B(n22844), .Z(n22705) );
  XOR U22837 ( .A(n22839), .B(n22845), .Z(n22680) );
  XNOR U22838 ( .A(n22846), .B(n22847), .Z(n22845) );
  OR U22839 ( .A(n22701), .B(n22848), .Z(n22847) );
  XNOR U22840 ( .A(n22696), .B(n22849), .Z(n22839) );
  XNOR U22841 ( .A(n22850), .B(n22851), .Z(n22849) );
  NAND U22842 ( .A(n22852), .B(n22791), .Z(n22851) );
  XNOR U22843 ( .A(n22834), .B(n22833), .Z(n22837) );
  IV U22844 ( .A(n22683), .Z(n22833) );
  XNOR U22845 ( .A(n22696), .B(n22853), .Z(n22834) );
  XOR U22846 ( .A(n22854), .B(n22846), .Z(n22853) );
  OR U22847 ( .A(n22855), .B(n22856), .Z(n22846) );
  AND U22848 ( .A(n22857), .B(n22858), .Z(n22854) );
  XOR U22849 ( .A(n22859), .B(n22850), .Z(n22696) );
  NANDN U22850 ( .A(n22860), .B(n22861), .Z(n22850) );
  ANDN U22851 ( .B(n22862), .A(n22863), .Z(n22859) );
  XNOR U22852 ( .A(n19114), .B(n22864), .Z(n22794) );
  XNOR U22853 ( .A(key[475]), .B(n18238), .Z(n22864) );
  XOR U22854 ( .A(n18218), .B(n20289), .Z(n18238) );
  XNOR U22855 ( .A(n22727), .B(n20260), .Z(n20289) );
  IV U22856 ( .A(n22865), .Z(n20260) );
  IV U22857 ( .A(n22769), .Z(n18218) );
  XOR U22858 ( .A(n22727), .B(n22830), .Z(n22769) );
  XNOR U22859 ( .A(n22752), .B(n22866), .Z(n22727) );
  XOR U22860 ( .A(n22867), .B(n22868), .Z(n22866) );
  XNOR U22861 ( .A(n22871), .B(n22872), .Z(n22752) );
  XNOR U22862 ( .A(n22873), .B(n22874), .Z(n22872) );
  NANDN U22863 ( .A(n22875), .B(n22876), .Z(n22874) );
  XOR U22864 ( .A(n18242), .B(n19128), .Z(n19114) );
  XOR U22865 ( .A(n22662), .B(n19098), .Z(n19128) );
  IV U22866 ( .A(n22835), .Z(n19098) );
  XNOR U22867 ( .A(n22764), .B(n22767), .Z(n22835) );
  XOR U22868 ( .A(n22767), .B(n22662), .Z(n18242) );
  XNOR U22869 ( .A(n22738), .B(n22877), .Z(n22662) );
  XOR U22870 ( .A(n22878), .B(n22879), .Z(n22877) );
  ANDN U22871 ( .B(n22880), .A(n22881), .Z(n22878) );
  XOR U22872 ( .A(n22882), .B(n22883), .Z(n22738) );
  XNOR U22873 ( .A(n22884), .B(n22885), .Z(n22883) );
  NANDN U22874 ( .A(n22886), .B(n22887), .Z(n22885) );
  XOR U22875 ( .A(n22889), .B(n22740), .Z(n22888) );
  OR U22876 ( .A(n22890), .B(n22891), .Z(n22740) );
  NOR U22877 ( .A(n22892), .B(n22893), .Z(n22889) );
  XOR U22878 ( .A(n22894), .B(n22895), .Z(n22646) );
  XOR U22879 ( .A(n20258), .B(n19107), .Z(n22895) );
  XNOR U22880 ( .A(n22736), .B(n22896), .Z(n19107) );
  XNOR U22881 ( .A(n22766), .B(n22693), .Z(n22896) );
  XNOR U22882 ( .A(n22897), .B(n22898), .Z(n22693) );
  XNOR U22883 ( .A(n22899), .B(n22666), .Z(n22898) );
  ANDN U22884 ( .B(n22900), .A(n22901), .Z(n22666) );
  ANDN U22885 ( .B(n22880), .A(n22902), .Z(n22899) );
  XNOR U22886 ( .A(n22664), .B(n22903), .Z(n22766) );
  XNOR U22887 ( .A(n22904), .B(n22905), .Z(n22903) );
  NANDN U22888 ( .A(n22893), .B(n22906), .Z(n22905) );
  XNOR U22889 ( .A(n22764), .B(n22765), .Z(n22736) );
  XNOR U22890 ( .A(n22904), .B(n22908), .Z(n22907) );
  OR U22891 ( .A(n22742), .B(n22909), .Z(n22908) );
  OR U22892 ( .A(n22890), .B(n22910), .Z(n22904) );
  XNOR U22893 ( .A(n22742), .B(n22893), .Z(n22890) );
  XNOR U22894 ( .A(n22664), .B(n22911), .Z(n22897) );
  XNOR U22895 ( .A(n22912), .B(n22913), .Z(n22911) );
  NANDN U22896 ( .A(n22886), .B(n22914), .Z(n22913) );
  XOR U22897 ( .A(n22915), .B(n22912), .Z(n22664) );
  NANDN U22898 ( .A(n22916), .B(n22917), .Z(n22912) );
  ANDN U22899 ( .B(n22918), .A(n22919), .Z(n22915) );
  XOR U22900 ( .A(n22882), .B(n22920), .Z(n22764) );
  XNOR U22901 ( .A(n22879), .B(n22921), .Z(n22920) );
  NAND U22902 ( .A(n22922), .B(n22668), .Z(n22921) );
  XOR U22903 ( .A(n22880), .B(n22668), .Z(n22900) );
  XNOR U22904 ( .A(n22924), .B(n22884), .Z(n22882) );
  OR U22905 ( .A(n22916), .B(n22925), .Z(n22884) );
  XOR U22906 ( .A(n22926), .B(n22886), .Z(n22916) );
  XOR U22907 ( .A(n22893), .B(n22668), .Z(n22886) );
  XOR U22908 ( .A(n22927), .B(n22928), .Z(n22668) );
  NANDN U22909 ( .A(n22929), .B(n22930), .Z(n22928) );
  XNOR U22910 ( .A(n22931), .B(n22932), .Z(n22893) );
  OR U22911 ( .A(n22929), .B(n22933), .Z(n22932) );
  ANDN U22912 ( .B(n22926), .A(n22934), .Z(n22924) );
  IV U22913 ( .A(n22919), .Z(n22926) );
  XOR U22914 ( .A(n22742), .B(n22880), .Z(n22919) );
  XNOR U22915 ( .A(n22935), .B(n22927), .Z(n22880) );
  NANDN U22916 ( .A(n22936), .B(n22937), .Z(n22927) );
  ANDN U22917 ( .B(n22938), .A(n22939), .Z(n22935) );
  NANDN U22918 ( .A(n22936), .B(n22941), .Z(n22931) );
  XOR U22919 ( .A(n22942), .B(n22929), .Z(n22936) );
  XNOR U22920 ( .A(n22943), .B(n22944), .Z(n22929) );
  XOR U22921 ( .A(n22945), .B(n22938), .Z(n22944) );
  XNOR U22922 ( .A(n22946), .B(n22947), .Z(n22943) );
  XNOR U22923 ( .A(n22948), .B(n22949), .Z(n22947) );
  ANDN U22924 ( .B(n22938), .A(n22950), .Z(n22948) );
  IV U22925 ( .A(n22951), .Z(n22938) );
  ANDN U22926 ( .B(n22942), .A(n22950), .Z(n22940) );
  IV U22927 ( .A(n22946), .Z(n22950) );
  IV U22928 ( .A(n22939), .Z(n22942) );
  XNOR U22929 ( .A(n22945), .B(n22952), .Z(n22939) );
  XOR U22930 ( .A(n22953), .B(n22949), .Z(n22952) );
  NAND U22931 ( .A(n22941), .B(n22937), .Z(n22949) );
  XNOR U22932 ( .A(n22930), .B(n22951), .Z(n22937) );
  XOR U22933 ( .A(n22954), .B(n22955), .Z(n22951) );
  XOR U22934 ( .A(n22956), .B(n22957), .Z(n22955) );
  XNOR U22935 ( .A(n22906), .B(n22958), .Z(n22957) );
  XNOR U22936 ( .A(n22959), .B(n22960), .Z(n22954) );
  XNOR U22937 ( .A(n22961), .B(n22962), .Z(n22960) );
  ANDN U22938 ( .B(n22963), .A(n22743), .Z(n22961) );
  XNOR U22939 ( .A(n22946), .B(n22933), .Z(n22941) );
  XOR U22940 ( .A(n22964), .B(n22965), .Z(n22946) );
  XNOR U22941 ( .A(n22966), .B(n22958), .Z(n22965) );
  XOR U22942 ( .A(n22967), .B(n22968), .Z(n22958) );
  XNOR U22943 ( .A(n22969), .B(n22970), .Z(n22968) );
  NAND U22944 ( .A(n22887), .B(n22914), .Z(n22970) );
  XNOR U22945 ( .A(n22971), .B(n22972), .Z(n22964) );
  ANDN U22946 ( .B(n22973), .A(n22881), .Z(n22971) );
  ANDN U22947 ( .B(n22930), .A(n22933), .Z(n22953) );
  XOR U22948 ( .A(n22933), .B(n22930), .Z(n22945) );
  XNOR U22949 ( .A(n22974), .B(n22975), .Z(n22930) );
  XNOR U22950 ( .A(n22967), .B(n22976), .Z(n22975) );
  XOR U22951 ( .A(n22966), .B(n22909), .Z(n22976) );
  XOR U22952 ( .A(n22743), .B(n22977), .Z(n22974) );
  XNOR U22953 ( .A(n22978), .B(n22962), .Z(n22977) );
  OR U22954 ( .A(n22910), .B(n22891), .Z(n22962) );
  XNOR U22955 ( .A(n22743), .B(n22892), .Z(n22891) );
  XOR U22956 ( .A(n22909), .B(n22906), .Z(n22910) );
  ANDN U22957 ( .B(n22906), .A(n22892), .Z(n22978) );
  XOR U22958 ( .A(n22979), .B(n22980), .Z(n22933) );
  XOR U22959 ( .A(n22967), .B(n22956), .Z(n22980) );
  XOR U22960 ( .A(n22922), .B(n22669), .Z(n22956) );
  XOR U22961 ( .A(n22981), .B(n22969), .Z(n22967) );
  NANDN U22962 ( .A(n22925), .B(n22917), .Z(n22969) );
  XOR U22963 ( .A(n22918), .B(n22914), .Z(n22917) );
  XNOR U22964 ( .A(n22973), .B(n22982), .Z(n22906) );
  XOR U22965 ( .A(n22983), .B(n22984), .Z(n22982) );
  XOR U22966 ( .A(n22934), .B(n22887), .Z(n22925) );
  XNOR U22967 ( .A(n22892), .B(n22922), .Z(n22887) );
  IV U22968 ( .A(n22959), .Z(n22892) );
  XOR U22969 ( .A(n22985), .B(n22986), .Z(n22959) );
  XOR U22970 ( .A(n22987), .B(n22988), .Z(n22986) );
  XNOR U22971 ( .A(n22743), .B(n22989), .Z(n22985) );
  ANDN U22972 ( .B(n22918), .A(n22934), .Z(n22981) );
  XNOR U22973 ( .A(n22743), .B(n22881), .Z(n22934) );
  XOR U22974 ( .A(n22973), .B(n22963), .Z(n22918) );
  IV U22975 ( .A(n22909), .Z(n22963) );
  XOR U22976 ( .A(n22990), .B(n22991), .Z(n22909) );
  XOR U22977 ( .A(n22992), .B(n22988), .Z(n22991) );
  XNOR U22978 ( .A(n22993), .B(n22994), .Z(n22988) );
  XOR U22979 ( .A(n21222), .B(n22228), .Z(n22994) );
  XNOR U22980 ( .A(n22995), .B(n22996), .Z(n22228) );
  XOR U22981 ( .A(n22231), .B(n22997), .Z(n21222) );
  XNOR U22982 ( .A(n21221), .B(n22998), .Z(n22993) );
  XNOR U22983 ( .A(key[348]), .B(n22999), .Z(n22998) );
  XOR U22984 ( .A(n22246), .B(n21209), .Z(n21221) );
  IV U22985 ( .A(n22902), .Z(n22973) );
  XOR U22986 ( .A(n22966), .B(n23000), .Z(n22979) );
  XNOR U22987 ( .A(n23001), .B(n22972), .Z(n23000) );
  OR U22988 ( .A(n22901), .B(n22923), .Z(n22972) );
  XNOR U22989 ( .A(n23002), .B(n22922), .Z(n22923) );
  XNOR U22990 ( .A(n22902), .B(n22669), .Z(n22901) );
  ANDN U22991 ( .B(n22922), .A(n22669), .Z(n23001) );
  XOR U22992 ( .A(n22990), .B(n23003), .Z(n22669) );
  XNOR U22993 ( .A(n23004), .B(n22992), .Z(n23003) );
  XOR U22994 ( .A(n22992), .B(n22990), .Z(n22922) );
  XNOR U22995 ( .A(n22881), .B(n22902), .Z(n22966) );
  XOR U22996 ( .A(n22990), .B(n23005), .Z(n22902) );
  XNOR U22997 ( .A(n22992), .B(n22987), .Z(n23005) );
  XOR U22998 ( .A(n23006), .B(n23007), .Z(n22987) );
  XNOR U22999 ( .A(n23008), .B(n21217), .Z(n23007) );
  XNOR U23000 ( .A(n23009), .B(n23010), .Z(n21217) );
  XOR U23001 ( .A(key[351]), .B(n21243), .Z(n23006) );
  XNOR U23002 ( .A(n23011), .B(n23012), .Z(n22990) );
  XNOR U23003 ( .A(n23013), .B(n21210), .Z(n23012) );
  XNOR U23004 ( .A(n22217), .B(n22996), .Z(n21210) );
  XNOR U23005 ( .A(n21206), .B(n23014), .Z(n23011) );
  XNOR U23006 ( .A(key[349]), .B(n23015), .Z(n23014) );
  IV U23007 ( .A(n23002), .Z(n22881) );
  XNOR U23008 ( .A(n22984), .B(n23016), .Z(n23002) );
  XOR U23009 ( .A(n23017), .B(n23018), .Z(n22992) );
  XOR U23010 ( .A(n22743), .B(n22209), .Z(n23018) );
  XOR U23011 ( .A(n22224), .B(n23010), .Z(n22209) );
  XNOR U23012 ( .A(n23019), .B(n23020), .Z(n22743) );
  XOR U23013 ( .A(n23021), .B(n22245), .Z(n23020) );
  XNOR U23014 ( .A(n23022), .B(n23023), .Z(n23019) );
  XOR U23015 ( .A(key[344]), .B(n22995), .Z(n23023) );
  IV U23016 ( .A(n22224), .Z(n22995) );
  XOR U23017 ( .A(n21203), .B(n23024), .Z(n23017) );
  XNOR U23018 ( .A(key[350]), .B(n23025), .Z(n23024) );
  XNOR U23019 ( .A(n22216), .B(n21216), .Z(n21203) );
  XOR U23020 ( .A(n22246), .B(n23026), .Z(n21216) );
  XOR U23021 ( .A(n23015), .B(n22210), .Z(n22216) );
  XOR U23022 ( .A(n23027), .B(n23028), .Z(n22989) );
  XOR U23023 ( .A(n22236), .B(n23029), .Z(n23028) );
  XNOR U23024 ( .A(n21228), .B(n23004), .Z(n23029) );
  IV U23025 ( .A(n22983), .Z(n23004) );
  XNOR U23026 ( .A(n23030), .B(n23031), .Z(n22983) );
  XNOR U23027 ( .A(n23032), .B(n21234), .Z(n23031) );
  XNOR U23028 ( .A(n22239), .B(n23033), .Z(n21234) );
  XNOR U23029 ( .A(n23034), .B(n23035), .Z(n23030) );
  XNOR U23030 ( .A(key[345]), .B(n23036), .Z(n23035) );
  XNOR U23031 ( .A(n22246), .B(n21225), .Z(n21228) );
  XOR U23032 ( .A(n22224), .B(n22997), .Z(n22236) );
  XOR U23033 ( .A(n21230), .B(n23037), .Z(n23027) );
  XNOR U23034 ( .A(key[347]), .B(n23038), .Z(n23037) );
  XNOR U23035 ( .A(n23039), .B(n22235), .Z(n21230) );
  XOR U23036 ( .A(n23040), .B(n23041), .Z(n22984) );
  XNOR U23037 ( .A(n23042), .B(n21195), .Z(n23041) );
  XOR U23038 ( .A(n22202), .B(n23032), .Z(n21195) );
  XNOR U23039 ( .A(n23039), .B(n23043), .Z(n23040) );
  XNOR U23040 ( .A(key[346]), .B(n21238), .Z(n23043) );
  XOR U23041 ( .A(n22781), .B(n22683), .Z(n20258) );
  XNOR U23042 ( .A(n22787), .B(n23044), .Z(n22683) );
  XNOR U23043 ( .A(n22784), .B(n23045), .Z(n23044) );
  NAND U23044 ( .A(n23046), .B(n22706), .Z(n23045) );
  NANDN U23045 ( .A(n23047), .B(n22844), .Z(n22784) );
  XNOR U23046 ( .A(n22786), .B(n22706), .Z(n22844) );
  XOR U23047 ( .A(n22787), .B(n23048), .Z(n22781) );
  XOR U23048 ( .A(n23049), .B(n22699), .Z(n23048) );
  OR U23049 ( .A(n23050), .B(n22855), .Z(n22699) );
  XOR U23050 ( .A(n22701), .B(n22858), .Z(n22855) );
  ANDN U23051 ( .B(n22858), .A(n23051), .Z(n23049) );
  XOR U23052 ( .A(n23052), .B(n22789), .Z(n22787) );
  OR U23053 ( .A(n23053), .B(n22860), .Z(n22789) );
  XOR U23054 ( .A(n22863), .B(n22791), .Z(n22860) );
  XOR U23055 ( .A(n22858), .B(n22706), .Z(n22791) );
  XOR U23056 ( .A(n23054), .B(n23055), .Z(n22706) );
  NANDN U23057 ( .A(n23056), .B(n23057), .Z(n23055) );
  XOR U23058 ( .A(n23058), .B(n23059), .Z(n22858) );
  OR U23059 ( .A(n23056), .B(n23060), .Z(n23059) );
  IV U23060 ( .A(n23061), .Z(n22863) );
  ANDN U23061 ( .B(n23061), .A(n23062), .Z(n23052) );
  XOR U23062 ( .A(n22701), .B(n22786), .Z(n23061) );
  XOR U23063 ( .A(n23063), .B(n23054), .Z(n22786) );
  NANDN U23064 ( .A(n23064), .B(n23065), .Z(n23054) );
  ANDN U23065 ( .B(n23066), .A(n23067), .Z(n23063) );
  NANDN U23066 ( .A(n23064), .B(n23069), .Z(n23058) );
  XOR U23067 ( .A(n23070), .B(n23056), .Z(n23064) );
  XNOR U23068 ( .A(n23071), .B(n23072), .Z(n23056) );
  XOR U23069 ( .A(n23073), .B(n23066), .Z(n23072) );
  XNOR U23070 ( .A(n23074), .B(n23075), .Z(n23071) );
  XNOR U23071 ( .A(n23076), .B(n23077), .Z(n23075) );
  ANDN U23072 ( .B(n23066), .A(n23078), .Z(n23076) );
  IV U23073 ( .A(n23079), .Z(n23066) );
  ANDN U23074 ( .B(n23070), .A(n23078), .Z(n23068) );
  IV U23075 ( .A(n23074), .Z(n23078) );
  IV U23076 ( .A(n23067), .Z(n23070) );
  XNOR U23077 ( .A(n23073), .B(n23080), .Z(n23067) );
  XOR U23078 ( .A(n23081), .B(n23077), .Z(n23080) );
  NAND U23079 ( .A(n23069), .B(n23065), .Z(n23077) );
  XNOR U23080 ( .A(n23057), .B(n23079), .Z(n23065) );
  XOR U23081 ( .A(n23082), .B(n23083), .Z(n23079) );
  XOR U23082 ( .A(n23084), .B(n23085), .Z(n23083) );
  XNOR U23083 ( .A(n22857), .B(n23086), .Z(n23085) );
  XNOR U23084 ( .A(n23087), .B(n23088), .Z(n23082) );
  XNOR U23085 ( .A(n23089), .B(n23090), .Z(n23088) );
  ANDN U23086 ( .B(n23091), .A(n22702), .Z(n23089) );
  XNOR U23087 ( .A(n23074), .B(n23060), .Z(n23069) );
  XOR U23088 ( .A(n23092), .B(n23093), .Z(n23074) );
  XNOR U23089 ( .A(n23094), .B(n23086), .Z(n23093) );
  XOR U23090 ( .A(n23095), .B(n23096), .Z(n23086) );
  XNOR U23091 ( .A(n23097), .B(n23098), .Z(n23096) );
  NAND U23092 ( .A(n22792), .B(n22852), .Z(n23098) );
  XNOR U23093 ( .A(n23099), .B(n23100), .Z(n23092) );
  ANDN U23094 ( .B(n23101), .A(n22785), .Z(n23099) );
  ANDN U23095 ( .B(n23057), .A(n23060), .Z(n23081) );
  XOR U23096 ( .A(n23060), .B(n23057), .Z(n23073) );
  XNOR U23097 ( .A(n23102), .B(n23103), .Z(n23057) );
  XNOR U23098 ( .A(n23095), .B(n23104), .Z(n23103) );
  XOR U23099 ( .A(n23094), .B(n22848), .Z(n23104) );
  XOR U23100 ( .A(n22702), .B(n23105), .Z(n23102) );
  XNOR U23101 ( .A(n23106), .B(n23090), .Z(n23105) );
  OR U23102 ( .A(n22856), .B(n23050), .Z(n23090) );
  XNOR U23103 ( .A(n22702), .B(n23051), .Z(n23050) );
  XOR U23104 ( .A(n22848), .B(n22857), .Z(n22856) );
  ANDN U23105 ( .B(n22857), .A(n23051), .Z(n23106) );
  XOR U23106 ( .A(n23107), .B(n23108), .Z(n23060) );
  XOR U23107 ( .A(n23095), .B(n23084), .Z(n23108) );
  XOR U23108 ( .A(n23046), .B(n22707), .Z(n23084) );
  XOR U23109 ( .A(n23109), .B(n23097), .Z(n23095) );
  NANDN U23110 ( .A(n23053), .B(n22861), .Z(n23097) );
  XOR U23111 ( .A(n22862), .B(n22852), .Z(n22861) );
  XNOR U23112 ( .A(n23101), .B(n23110), .Z(n22857) );
  XOR U23113 ( .A(n23111), .B(n23112), .Z(n23110) );
  XOR U23114 ( .A(n23062), .B(n22792), .Z(n23053) );
  XNOR U23115 ( .A(n23051), .B(n23046), .Z(n22792) );
  IV U23116 ( .A(n23087), .Z(n23051) );
  XOR U23117 ( .A(n23113), .B(n23114), .Z(n23087) );
  XOR U23118 ( .A(n23115), .B(n23116), .Z(n23114) );
  XNOR U23119 ( .A(n22702), .B(n23117), .Z(n23113) );
  ANDN U23120 ( .B(n22862), .A(n23062), .Z(n23109) );
  XNOR U23121 ( .A(n22702), .B(n22785), .Z(n23062) );
  XOR U23122 ( .A(n23101), .B(n23091), .Z(n22862) );
  IV U23123 ( .A(n22848), .Z(n23091) );
  XOR U23124 ( .A(n23118), .B(n23119), .Z(n22848) );
  XOR U23125 ( .A(n23120), .B(n23116), .Z(n23119) );
  XNOR U23126 ( .A(n23121), .B(n22388), .Z(n23116) );
  XOR U23127 ( .A(n23122), .B(n23123), .Z(n22388) );
  XNOR U23128 ( .A(n21347), .B(n23124), .Z(n23123) );
  XOR U23129 ( .A(n23125), .B(n23126), .Z(n23122) );
  XNOR U23130 ( .A(n21344), .B(n23127), .Z(n23121) );
  XOR U23131 ( .A(key[356]), .B(n23128), .Z(n23127) );
  XOR U23132 ( .A(n23129), .B(n22404), .Z(n21344) );
  IV U23133 ( .A(n22842), .Z(n23101) );
  XOR U23134 ( .A(n23094), .B(n23130), .Z(n23107) );
  XNOR U23135 ( .A(n23131), .B(n23100), .Z(n23130) );
  OR U23136 ( .A(n22843), .B(n23047), .Z(n23100) );
  XNOR U23137 ( .A(n23132), .B(n23046), .Z(n23047) );
  XNOR U23138 ( .A(n22842), .B(n22707), .Z(n22843) );
  ANDN U23139 ( .B(n23046), .A(n22707), .Z(n23131) );
  XOR U23140 ( .A(n23118), .B(n23133), .Z(n22707) );
  XNOR U23141 ( .A(n23112), .B(n23134), .Z(n23133) );
  XOR U23142 ( .A(n23120), .B(n23118), .Z(n23046) );
  XNOR U23143 ( .A(n22785), .B(n22842), .Z(n23094) );
  XOR U23144 ( .A(n23118), .B(n23135), .Z(n22842) );
  XNOR U23145 ( .A(n23120), .B(n23115), .Z(n23135) );
  XOR U23146 ( .A(n23136), .B(n23137), .Z(n23115) );
  XNOR U23147 ( .A(n23138), .B(n22384), .Z(n23137) );
  XNOR U23148 ( .A(n21356), .B(n23139), .Z(n22384) );
  XNOR U23149 ( .A(key[359]), .B(n23129), .Z(n23136) );
  XNOR U23150 ( .A(n23140), .B(n23141), .Z(n23118) );
  XNOR U23151 ( .A(n23126), .B(n22405), .Z(n23141) );
  XOR U23152 ( .A(n21361), .B(n23142), .Z(n22405) );
  XNOR U23153 ( .A(key[357]), .B(n23143), .Z(n23140) );
  IV U23154 ( .A(n23132), .Z(n22785) );
  XOR U23155 ( .A(n23134), .B(n23144), .Z(n23132) );
  XNOR U23156 ( .A(n23111), .B(n23117), .Z(n23144) );
  XOR U23157 ( .A(n23145), .B(n23146), .Z(n23117) );
  XOR U23158 ( .A(n23112), .B(n23147), .Z(n23146) );
  XOR U23159 ( .A(n21382), .B(n22373), .Z(n23147) );
  XNOR U23160 ( .A(n23148), .B(n23128), .Z(n22373) );
  XNOR U23161 ( .A(n23129), .B(n22389), .Z(n21382) );
  XNOR U23162 ( .A(n23149), .B(n23150), .Z(n23112) );
  XOR U23163 ( .A(n22398), .B(n21398), .Z(n23150) );
  XOR U23164 ( .A(key[353]), .B(n22378), .Z(n23149) );
  XOR U23165 ( .A(n22372), .B(n23151), .Z(n23145) );
  XOR U23166 ( .A(key[355]), .B(n23152), .Z(n23151) );
  XOR U23167 ( .A(n23153), .B(n23154), .Z(n23111) );
  XOR U23168 ( .A(n21392), .B(n22376), .Z(n23154) );
  XOR U23169 ( .A(key[354]), .B(n22363), .Z(n23153) );
  IV U23170 ( .A(n23120), .Z(n23134) );
  XOR U23171 ( .A(n23155), .B(n23156), .Z(n23120) );
  XNOR U23172 ( .A(n22702), .B(n22394), .Z(n23156) );
  XOR U23173 ( .A(n23157), .B(n23138), .Z(n22394) );
  XOR U23174 ( .A(n23125), .B(n23158), .Z(n23138) );
  XNOR U23175 ( .A(n23159), .B(n23160), .Z(n22702) );
  XOR U23176 ( .A(n21387), .B(n21373), .Z(n23160) );
  XNOR U23177 ( .A(n23148), .B(n22397), .Z(n21373) );
  XNOR U23178 ( .A(key[352]), .B(n23161), .Z(n23159) );
  XNOR U23179 ( .A(n21369), .B(n23162), .Z(n23155) );
  XOR U23180 ( .A(key[358]), .B(n23163), .Z(n23162) );
  XNOR U23181 ( .A(n23129), .B(n22385), .Z(n21369) );
  XNOR U23182 ( .A(n18233), .B(n23164), .Z(n22894) );
  XOR U23183 ( .A(key[474]), .B(n20300), .Z(n23164) );
  XNOR U23184 ( .A(n23165), .B(n23166), .Z(n20300) );
  XOR U23185 ( .A(n22831), .B(n22749), .Z(n23166) );
  XNOR U23186 ( .A(n23167), .B(n23168), .Z(n22749) );
  XNOR U23187 ( .A(n23169), .B(n22729), .Z(n23168) );
  ANDN U23188 ( .B(n23170), .A(n23171), .Z(n22729) );
  ANDN U23189 ( .B(n22870), .A(n23172), .Z(n23169) );
  XOR U23190 ( .A(n22725), .B(n23173), .Z(n22831) );
  XNOR U23191 ( .A(n23174), .B(n23175), .Z(n23173) );
  NANDN U23192 ( .A(n23176), .B(n23177), .Z(n23175) );
  XNOR U23193 ( .A(n22829), .B(n22759), .Z(n23165) );
  XNOR U23194 ( .A(n23174), .B(n23179), .Z(n23178) );
  NANDN U23195 ( .A(n23180), .B(n22757), .Z(n23179) );
  OR U23196 ( .A(n23181), .B(n23182), .Z(n23174) );
  XNOR U23197 ( .A(n22725), .B(n23183), .Z(n23167) );
  XNOR U23198 ( .A(n23184), .B(n23185), .Z(n23183) );
  NANDN U23199 ( .A(n22875), .B(n23186), .Z(n23185) );
  XOR U23200 ( .A(n23187), .B(n23184), .Z(n22725) );
  NANDN U23201 ( .A(n23188), .B(n23189), .Z(n23184) );
  ANDN U23202 ( .B(n23190), .A(n23191), .Z(n23187) );
  IV U23203 ( .A(n22758), .Z(n22829) );
  IV U23204 ( .A(n19097), .Z(n18233) );
  XOR U23205 ( .A(n22865), .B(n18194), .Z(n19097) );
  XNOR U23206 ( .A(n22746), .B(n22689), .Z(n18194) );
  XOR U23207 ( .A(n22775), .B(n23192), .Z(n22689) );
  XNOR U23208 ( .A(n22771), .B(n23193), .Z(n23192) );
  NANDN U23209 ( .A(n22722), .B(n23194), .Z(n23193) );
  OR U23210 ( .A(n23195), .B(n22803), .Z(n22771) );
  XNOR U23211 ( .A(n22774), .B(n23196), .Z(n22803) );
  XNOR U23212 ( .A(n22775), .B(n23197), .Z(n22746) );
  XOR U23213 ( .A(n23198), .B(n22714), .Z(n23197) );
  OR U23214 ( .A(n23199), .B(n22816), .Z(n22714) );
  XOR U23215 ( .A(n22717), .B(n22812), .Z(n22816) );
  NOR U23216 ( .A(n23200), .B(n22812), .Z(n23198) );
  XOR U23217 ( .A(n23201), .B(n22777), .Z(n22775) );
  OR U23218 ( .A(n23202), .B(n22824), .Z(n22777) );
  XOR U23219 ( .A(n22827), .B(n22779), .Z(n22824) );
  XOR U23220 ( .A(n22812), .B(n22722), .Z(n22779) );
  IV U23221 ( .A(n23196), .Z(n22722) );
  XOR U23222 ( .A(n23203), .B(n23204), .Z(n23196) );
  NANDN U23223 ( .A(n23205), .B(n23206), .Z(n23204) );
  XNOR U23224 ( .A(n23207), .B(n23208), .Z(n22812) );
  OR U23225 ( .A(n23205), .B(n23209), .Z(n23208) );
  ANDN U23226 ( .B(n23210), .A(n22827), .Z(n23201) );
  XNOR U23227 ( .A(n22717), .B(n22774), .Z(n22827) );
  XOR U23228 ( .A(n23203), .B(n23211), .Z(n22774) );
  NANDN U23229 ( .A(n23212), .B(n23213), .Z(n23211) );
  NANDN U23230 ( .A(n23214), .B(n23215), .Z(n23203) );
  OR U23231 ( .A(n23217), .B(n23214), .Z(n23207) );
  XOR U23232 ( .A(n23218), .B(n23205), .Z(n23214) );
  XNOR U23233 ( .A(n23219), .B(n23220), .Z(n23205) );
  XOR U23234 ( .A(n23221), .B(n23213), .Z(n23220) );
  XNOR U23235 ( .A(n23222), .B(n23223), .Z(n23219) );
  XNOR U23236 ( .A(n23224), .B(n23225), .Z(n23223) );
  ANDN U23237 ( .B(n23213), .A(n23226), .Z(n23224) );
  IV U23238 ( .A(n23227), .Z(n23213) );
  ANDN U23239 ( .B(n23218), .A(n23226), .Z(n23216) );
  IV U23240 ( .A(n23212), .Z(n23218) );
  XNOR U23241 ( .A(n23221), .B(n23228), .Z(n23212) );
  XNOR U23242 ( .A(n23225), .B(n23229), .Z(n23228) );
  NANDN U23243 ( .A(n23209), .B(n23206), .Z(n23229) );
  NANDN U23244 ( .A(n23217), .B(n23215), .Z(n23225) );
  XNOR U23245 ( .A(n23206), .B(n23227), .Z(n23215) );
  XOR U23246 ( .A(n23230), .B(n23231), .Z(n23227) );
  XOR U23247 ( .A(n23232), .B(n23233), .Z(n23231) );
  XNOR U23248 ( .A(n22813), .B(n23234), .Z(n23233) );
  XNOR U23249 ( .A(n23235), .B(n23236), .Z(n23230) );
  XNOR U23250 ( .A(n23237), .B(n23238), .Z(n23236) );
  ANDN U23251 ( .B(n22818), .A(n22716), .Z(n23237) );
  XNOR U23252 ( .A(n23226), .B(n23209), .Z(n23217) );
  IV U23253 ( .A(n23222), .Z(n23226) );
  XOR U23254 ( .A(n23239), .B(n23240), .Z(n23222) );
  XNOR U23255 ( .A(n23241), .B(n23234), .Z(n23240) );
  XOR U23256 ( .A(n23242), .B(n23243), .Z(n23234) );
  XNOR U23257 ( .A(n23244), .B(n23245), .Z(n23243) );
  NAND U23258 ( .A(n22780), .B(n22822), .Z(n23245) );
  XNOR U23259 ( .A(n23246), .B(n23247), .Z(n23239) );
  ANDN U23260 ( .B(n23248), .A(n22773), .Z(n23246) );
  XOR U23261 ( .A(n23209), .B(n23206), .Z(n23221) );
  XNOR U23262 ( .A(n23249), .B(n23250), .Z(n23206) );
  XNOR U23263 ( .A(n23242), .B(n23251), .Z(n23250) );
  XNOR U23264 ( .A(n23241), .B(n22818), .Z(n23251) );
  XNOR U23265 ( .A(n23252), .B(n23253), .Z(n23249) );
  XNOR U23266 ( .A(n23254), .B(n23238), .Z(n23253) );
  OR U23267 ( .A(n22817), .B(n23199), .Z(n23238) );
  XNOR U23268 ( .A(n23252), .B(n23235), .Z(n23199) );
  XNOR U23269 ( .A(n22818), .B(n22813), .Z(n22817) );
  ANDN U23270 ( .B(n22813), .A(n23200), .Z(n23254) );
  XOR U23271 ( .A(n23255), .B(n23256), .Z(n23209) );
  XOR U23272 ( .A(n23242), .B(n23232), .Z(n23256) );
  XNOR U23273 ( .A(n23194), .B(n22721), .Z(n23232) );
  XOR U23274 ( .A(n23257), .B(n23244), .Z(n23242) );
  NANDN U23275 ( .A(n23202), .B(n22825), .Z(n23244) );
  XOR U23276 ( .A(n22826), .B(n22822), .Z(n22825) );
  XOR U23277 ( .A(n22721), .B(n22813), .Z(n22822) );
  XNOR U23278 ( .A(n23248), .B(n23258), .Z(n22813) );
  XOR U23279 ( .A(n23259), .B(n23260), .Z(n23258) );
  XNOR U23280 ( .A(n23210), .B(n22780), .Z(n23202) );
  XNOR U23281 ( .A(n23200), .B(n23194), .Z(n22780) );
  IV U23282 ( .A(n23235), .Z(n23200) );
  XOR U23283 ( .A(n23261), .B(n23262), .Z(n23235) );
  XOR U23284 ( .A(n23263), .B(n23264), .Z(n23262) );
  XOR U23285 ( .A(n23252), .B(n23265), .Z(n23261) );
  AND U23286 ( .A(n22826), .B(n23210), .Z(n23257) );
  XOR U23287 ( .A(n23248), .B(n22818), .Z(n22826) );
  XNOR U23288 ( .A(n23266), .B(n23267), .Z(n22818) );
  XOR U23289 ( .A(n23268), .B(n23264), .Z(n23267) );
  XNOR U23290 ( .A(n23269), .B(n23270), .Z(n23264) );
  XOR U23291 ( .A(n21526), .B(n22558), .Z(n23270) );
  XNOR U23292 ( .A(n22554), .B(n23271), .Z(n22558) );
  XNOR U23293 ( .A(n23272), .B(n23273), .Z(n21526) );
  XNOR U23294 ( .A(n23274), .B(n21547), .Z(n23273) );
  XOR U23295 ( .A(n22577), .B(n22561), .Z(n23272) );
  XOR U23296 ( .A(key[268]), .B(n23275), .Z(n23269) );
  XOR U23297 ( .A(n23241), .B(n23276), .Z(n23255) );
  XNOR U23298 ( .A(n23277), .B(n23247), .Z(n23276) );
  OR U23299 ( .A(n22804), .B(n23195), .Z(n23247) );
  XNOR U23300 ( .A(n23278), .B(n23194), .Z(n23195) );
  XNOR U23301 ( .A(n23248), .B(n22721), .Z(n22804) );
  IV U23302 ( .A(n22805), .Z(n23248) );
  AND U23303 ( .A(n22721), .B(n23194), .Z(n23277) );
  XOR U23304 ( .A(n23268), .B(n23266), .Z(n23194) );
  XNOR U23305 ( .A(n23266), .B(n23279), .Z(n22721) );
  XNOR U23306 ( .A(n23260), .B(n23280), .Z(n23279) );
  XNOR U23307 ( .A(n22773), .B(n22805), .Z(n23241) );
  XOR U23308 ( .A(n23266), .B(n23281), .Z(n22805) );
  XNOR U23309 ( .A(n23268), .B(n23263), .Z(n23281) );
  XOR U23310 ( .A(n23282), .B(n23283), .Z(n23263) );
  XNOR U23311 ( .A(n23284), .B(n21532), .Z(n23283) );
  XNOR U23312 ( .A(n23285), .B(n23286), .Z(n21532) );
  XNOR U23313 ( .A(key[271]), .B(n21541), .Z(n23282) );
  XNOR U23314 ( .A(n23287), .B(n23288), .Z(n23266) );
  XNOR U23315 ( .A(n23289), .B(n21548), .Z(n23288) );
  XNOR U23316 ( .A(n22547), .B(n23271), .Z(n21548) );
  XOR U23317 ( .A(n21544), .B(n23290), .Z(n23287) );
  XNOR U23318 ( .A(key[269]), .B(n23291), .Z(n23290) );
  XOR U23319 ( .A(n22716), .B(n22773), .Z(n23210) );
  IV U23320 ( .A(n23278), .Z(n22773) );
  XOR U23321 ( .A(n23280), .B(n23292), .Z(n23278) );
  XNOR U23322 ( .A(n23259), .B(n23265), .Z(n23292) );
  XOR U23323 ( .A(n23293), .B(n23294), .Z(n23265) );
  XOR U23324 ( .A(n23260), .B(n23295), .Z(n23294) );
  XOR U23325 ( .A(n21506), .B(n22566), .Z(n23295) );
  XOR U23326 ( .A(n22554), .B(n23274), .Z(n22566) );
  XOR U23327 ( .A(n22577), .B(n21527), .Z(n21506) );
  XNOR U23328 ( .A(n23296), .B(n23297), .Z(n23260) );
  XOR U23329 ( .A(n23298), .B(n21512), .Z(n23297) );
  IV U23330 ( .A(n22576), .Z(n21512) );
  XNOR U23331 ( .A(n23299), .B(n23300), .Z(n22576) );
  XNOR U23332 ( .A(n21519), .B(n23301), .Z(n23296) );
  XNOR U23333 ( .A(key[265]), .B(n23302), .Z(n23301) );
  XOR U23334 ( .A(n21508), .B(n23303), .Z(n23293) );
  XNOR U23335 ( .A(key[267]), .B(n23304), .Z(n23303) );
  XNOR U23336 ( .A(n23305), .B(n22565), .Z(n21508) );
  XOR U23337 ( .A(n23306), .B(n23307), .Z(n23259) );
  XOR U23338 ( .A(n21516), .B(n21520), .Z(n23307) );
  XNOR U23339 ( .A(n23308), .B(n23298), .Z(n21520) );
  XNOR U23340 ( .A(n23309), .B(n23310), .Z(n23306) );
  XNOR U23341 ( .A(key[266]), .B(n23305), .Z(n23310) );
  IV U23342 ( .A(n23268), .Z(n23280) );
  XOR U23343 ( .A(n23311), .B(n23312), .Z(n23268) );
  XNOR U23344 ( .A(n23252), .B(n22539), .Z(n23312) );
  XNOR U23345 ( .A(n22554), .B(n23286), .Z(n22539) );
  XOR U23346 ( .A(n21536), .B(n23313), .Z(n23311) );
  XNOR U23347 ( .A(key[270]), .B(n23314), .Z(n23313) );
  XNOR U23348 ( .A(n22546), .B(n21531), .Z(n21536) );
  XOR U23349 ( .A(n22577), .B(n23315), .Z(n21531) );
  XOR U23350 ( .A(n23291), .B(n22540), .Z(n22546) );
  IV U23351 ( .A(n23316), .Z(n22540) );
  IV U23352 ( .A(n23252), .Z(n22716) );
  XOR U23353 ( .A(n23317), .B(n23318), .Z(n23252) );
  XNOR U23354 ( .A(n23319), .B(n23320), .Z(n23317) );
  XOR U23355 ( .A(key[264]), .B(n22554), .Z(n23320) );
  XOR U23356 ( .A(n22830), .B(n22758), .Z(n22865) );
  XOR U23357 ( .A(n22871), .B(n23321), .Z(n22758) );
  XNOR U23358 ( .A(n22868), .B(n23322), .Z(n23321) );
  NANDN U23359 ( .A(n23323), .B(n22731), .Z(n23322) );
  XOR U23360 ( .A(n22870), .B(n22731), .Z(n23170) );
  XOR U23361 ( .A(n22871), .B(n23325), .Z(n22830) );
  XOR U23362 ( .A(n23326), .B(n22754), .Z(n23325) );
  OR U23363 ( .A(n23327), .B(n23181), .Z(n22754) );
  XNOR U23364 ( .A(n22757), .B(n23177), .Z(n23181) );
  ANDN U23365 ( .B(n23177), .A(n23328), .Z(n23326) );
  XOR U23366 ( .A(n23329), .B(n22873), .Z(n22871) );
  OR U23367 ( .A(n23188), .B(n23330), .Z(n22873) );
  XNOR U23368 ( .A(n23191), .B(n22875), .Z(n23188) );
  XNOR U23369 ( .A(n23177), .B(n22731), .Z(n22875) );
  XOR U23370 ( .A(n23331), .B(n23332), .Z(n22731) );
  NANDN U23371 ( .A(n23333), .B(n23334), .Z(n23332) );
  XOR U23372 ( .A(n23335), .B(n23336), .Z(n23177) );
  NANDN U23373 ( .A(n23333), .B(n23337), .Z(n23336) );
  NOR U23374 ( .A(n23191), .B(n23338), .Z(n23329) );
  XNOR U23375 ( .A(n22870), .B(n22757), .Z(n23191) );
  XNOR U23376 ( .A(n23339), .B(n23335), .Z(n22757) );
  NANDN U23377 ( .A(n23340), .B(n23341), .Z(n23335) );
  XOR U23378 ( .A(n23337), .B(n23342), .Z(n23341) );
  ANDN U23379 ( .B(n23342), .A(n23343), .Z(n23339) );
  XNOR U23380 ( .A(n23344), .B(n23331), .Z(n22870) );
  NANDN U23381 ( .A(n23340), .B(n23345), .Z(n23331) );
  XOR U23382 ( .A(n23346), .B(n23334), .Z(n23345) );
  XNOR U23383 ( .A(n23347), .B(n23348), .Z(n23333) );
  XOR U23384 ( .A(n23349), .B(n23350), .Z(n23348) );
  XNOR U23385 ( .A(n23351), .B(n23352), .Z(n23347) );
  XNOR U23386 ( .A(n23353), .B(n23354), .Z(n23352) );
  ANDN U23387 ( .B(n23346), .A(n23350), .Z(n23353) );
  ANDN U23388 ( .B(n23346), .A(n23343), .Z(n23344) );
  XNOR U23389 ( .A(n23349), .B(n23355), .Z(n23343) );
  XOR U23390 ( .A(n23356), .B(n23354), .Z(n23355) );
  NAND U23391 ( .A(n23357), .B(n23358), .Z(n23354) );
  XNOR U23392 ( .A(n23351), .B(n23334), .Z(n23358) );
  IV U23393 ( .A(n23346), .Z(n23351) );
  XNOR U23394 ( .A(n23337), .B(n23350), .Z(n23357) );
  IV U23395 ( .A(n23342), .Z(n23350) );
  XOR U23396 ( .A(n23359), .B(n23360), .Z(n23342) );
  XNOR U23397 ( .A(n23361), .B(n23362), .Z(n23360) );
  XNOR U23398 ( .A(n23363), .B(n23364), .Z(n23359) );
  NOR U23399 ( .A(n23172), .B(n22869), .Z(n23363) );
  AND U23400 ( .A(n23334), .B(n23337), .Z(n23356) );
  XNOR U23401 ( .A(n23334), .B(n23337), .Z(n23349) );
  XNOR U23402 ( .A(n23365), .B(n23366), .Z(n23337) );
  XNOR U23403 ( .A(n23367), .B(n23362), .Z(n23366) );
  XOR U23404 ( .A(n23368), .B(n23369), .Z(n23365) );
  XNOR U23405 ( .A(n23370), .B(n23364), .Z(n23369) );
  OR U23406 ( .A(n23171), .B(n23324), .Z(n23364) );
  XNOR U23407 ( .A(n22869), .B(n23323), .Z(n23324) );
  XNOR U23408 ( .A(n23172), .B(n22732), .Z(n23171) );
  ANDN U23409 ( .B(n23371), .A(n23323), .Z(n23370) );
  XNOR U23410 ( .A(n23372), .B(n23373), .Z(n23334) );
  XNOR U23411 ( .A(n23362), .B(n23374), .Z(n23373) );
  XOR U23412 ( .A(n23180), .B(n23368), .Z(n23374) );
  XNOR U23413 ( .A(n22869), .B(n23375), .Z(n23362) );
  XOR U23414 ( .A(n22756), .B(n23376), .Z(n23372) );
  XNOR U23415 ( .A(n23377), .B(n23378), .Z(n23376) );
  ANDN U23416 ( .B(n23379), .A(n23328), .Z(n23377) );
  XNOR U23417 ( .A(n23380), .B(n23381), .Z(n23346) );
  XNOR U23418 ( .A(n23367), .B(n23382), .Z(n23381) );
  XNOR U23419 ( .A(n23176), .B(n23361), .Z(n23382) );
  XOR U23420 ( .A(n23368), .B(n23383), .Z(n23361) );
  XNOR U23421 ( .A(n23384), .B(n23385), .Z(n23383) );
  NAND U23422 ( .A(n22876), .B(n23186), .Z(n23385) );
  XNOR U23423 ( .A(n23386), .B(n23384), .Z(n23368) );
  NANDN U23424 ( .A(n23330), .B(n23189), .Z(n23384) );
  XOR U23425 ( .A(n23190), .B(n23186), .Z(n23189) );
  XNOR U23426 ( .A(n23379), .B(n22732), .Z(n23186) );
  XOR U23427 ( .A(n23338), .B(n22876), .Z(n23330) );
  XNOR U23428 ( .A(n23328), .B(n23387), .Z(n22876) );
  ANDN U23429 ( .B(n23190), .A(n23338), .Z(n23386) );
  XNOR U23430 ( .A(n22756), .B(n22869), .Z(n23338) );
  XOR U23431 ( .A(n23388), .B(n23389), .Z(n22869) );
  XNOR U23432 ( .A(n23390), .B(n23391), .Z(n23389) );
  XOR U23433 ( .A(n23387), .B(n23371), .Z(n23367) );
  IV U23434 ( .A(n22732), .Z(n23371) );
  XOR U23435 ( .A(n23392), .B(n23393), .Z(n22732) );
  XNOR U23436 ( .A(n23394), .B(n23391), .Z(n23393) );
  IV U23437 ( .A(n23323), .Z(n23387) );
  XOR U23438 ( .A(n23391), .B(n23395), .Z(n23323) );
  XNOR U23439 ( .A(n23396), .B(n23397), .Z(n23380) );
  XNOR U23440 ( .A(n23398), .B(n23378), .Z(n23397) );
  OR U23441 ( .A(n23182), .B(n23327), .Z(n23378) );
  XNOR U23442 ( .A(n22756), .B(n23328), .Z(n23327) );
  IV U23443 ( .A(n23396), .Z(n23328) );
  XOR U23444 ( .A(n23180), .B(n23379), .Z(n23182) );
  IV U23445 ( .A(n23176), .Z(n23379) );
  XOR U23446 ( .A(n23375), .B(n23399), .Z(n23176) );
  XNOR U23447 ( .A(n23394), .B(n23388), .Z(n23399) );
  XOR U23448 ( .A(n23400), .B(n23401), .Z(n23388) );
  XOR U23449 ( .A(n21684), .B(n22104), .Z(n23401) );
  XNOR U23450 ( .A(key[306]), .B(n22070), .Z(n23400) );
  IV U23451 ( .A(n23172), .Z(n23375) );
  XOR U23452 ( .A(n23392), .B(n23402), .Z(n23172) );
  XOR U23453 ( .A(n23391), .B(n23403), .Z(n23402) );
  NOR U23454 ( .A(n23180), .B(n22756), .Z(n23398) );
  XOR U23455 ( .A(n23392), .B(n23404), .Z(n23180) );
  XOR U23456 ( .A(n23391), .B(n23405), .Z(n23404) );
  XOR U23457 ( .A(n23406), .B(n23407), .Z(n23391) );
  XNOR U23458 ( .A(n22756), .B(n22077), .Z(n23407) );
  XNOR U23459 ( .A(n23408), .B(n23409), .Z(n22077) );
  XNOR U23460 ( .A(n21647), .B(n23410), .Z(n23406) );
  XOR U23461 ( .A(key[310]), .B(n22085), .Z(n23410) );
  XOR U23462 ( .A(n23411), .B(n22091), .Z(n21647) );
  IV U23463 ( .A(n23395), .Z(n23392) );
  XOR U23464 ( .A(n23412), .B(n23413), .Z(n23395) );
  XNOR U23465 ( .A(n23414), .B(n22083), .Z(n23413) );
  XOR U23466 ( .A(n21653), .B(n23415), .Z(n22083) );
  XNOR U23467 ( .A(key[309]), .B(n23416), .Z(n23412) );
  XOR U23468 ( .A(n23417), .B(n23418), .Z(n23396) );
  XNOR U23469 ( .A(n23405), .B(n23403), .Z(n23418) );
  XNOR U23470 ( .A(n23419), .B(n23420), .Z(n23403) );
  XOR U23471 ( .A(n23409), .B(n22090), .Z(n23420) );
  XNOR U23472 ( .A(n21662), .B(n23421), .Z(n22090) );
  XOR U23473 ( .A(n23422), .B(n23423), .Z(n23409) );
  XNOR U23474 ( .A(key[311]), .B(n23411), .Z(n23419) );
  XNOR U23475 ( .A(n23424), .B(n22093), .Z(n23405) );
  XOR U23476 ( .A(n23425), .B(n23426), .Z(n22093) );
  XNOR U23477 ( .A(n21671), .B(n23427), .Z(n23426) );
  XNOR U23478 ( .A(n21668), .B(n23428), .Z(n23424) );
  XOR U23479 ( .A(key[308]), .B(n23429), .Z(n23428) );
  XNOR U23480 ( .A(n23411), .B(n22082), .Z(n21668) );
  XNOR U23481 ( .A(n22756), .B(n23390), .Z(n23417) );
  XOR U23482 ( .A(n23430), .B(n23431), .Z(n23390) );
  XNOR U23483 ( .A(n23394), .B(n23432), .Z(n23431) );
  XOR U23484 ( .A(n21674), .B(n22101), .Z(n23432) );
  XNOR U23485 ( .A(n23422), .B(n23429), .Z(n22101) );
  XNOR U23486 ( .A(n23411), .B(n22094), .Z(n21674) );
  XOR U23487 ( .A(n23433), .B(n23434), .Z(n23394) );
  XOR U23488 ( .A(n22112), .B(n23435), .Z(n23434) );
  XOR U23489 ( .A(key[305]), .B(n22106), .Z(n23433) );
  XOR U23490 ( .A(n22100), .B(n23436), .Z(n23430) );
  XOR U23491 ( .A(key[307]), .B(n23437), .Z(n23436) );
  XNOR U23492 ( .A(n23438), .B(n23439), .Z(n22756) );
  XOR U23493 ( .A(n21679), .B(n21690), .Z(n23439) );
  XNOR U23494 ( .A(n23422), .B(n22111), .Z(n21690) );
  XNOR U23495 ( .A(key[304]), .B(n23440), .Z(n23438) );
  XOR U23496 ( .A(n23441), .B(n23442), .Z(n17102) );
  XNOR U23497 ( .A(n20617), .B(n20582), .Z(n23442) );
  XNOR U23498 ( .A(n23443), .B(n23444), .Z(n20582) );
  XNOR U23499 ( .A(n23445), .B(n20534), .Z(n23444) );
  NOR U23500 ( .A(n23446), .B(n23447), .Z(n20534) );
  ANDN U23501 ( .B(n20707), .A(n23448), .Z(n23445) );
  IV U23502 ( .A(n20603), .Z(n20617) );
  XOR U23503 ( .A(n23443), .B(n23449), .Z(n20603) );
  XOR U23504 ( .A(n23450), .B(n23451), .Z(n23449) );
  AND U23505 ( .A(n20609), .B(n23452), .Z(n23450) );
  XNOR U23506 ( .A(n20530), .B(n23453), .Z(n23443) );
  XNOR U23507 ( .A(n23454), .B(n23455), .Z(n23453) );
  NAND U23508 ( .A(n23456), .B(n20712), .Z(n23455) );
  XNOR U23509 ( .A(n20621), .B(n20619), .Z(n23441) );
  IV U23510 ( .A(n20610), .Z(n20619) );
  XNOR U23511 ( .A(n20708), .B(n23457), .Z(n20610) );
  XNOR U23512 ( .A(n20704), .B(n23458), .Z(n23457) );
  NANDN U23513 ( .A(n20537), .B(n23459), .Z(n23458) );
  OR U23514 ( .A(n23460), .B(n23446), .Z(n20704) );
  XNOR U23515 ( .A(n20707), .B(n23461), .Z(n23446) );
  XOR U23516 ( .A(n23462), .B(n20710), .Z(n20708) );
  OR U23517 ( .A(n23463), .B(n23464), .Z(n20710) );
  ANDN U23518 ( .B(n23465), .A(n23466), .Z(n23462) );
  XNOR U23519 ( .A(n20530), .B(n23467), .Z(n20621) );
  XNOR U23520 ( .A(n23451), .B(n23468), .Z(n23467) );
  NANDN U23521 ( .A(n20719), .B(n23469), .Z(n23468) );
  OR U23522 ( .A(n20717), .B(n23470), .Z(n23451) );
  XOR U23523 ( .A(n20609), .B(n20719), .Z(n20717) );
  XOR U23524 ( .A(n23471), .B(n23454), .Z(n20530) );
  NANDN U23525 ( .A(n23464), .B(n23472), .Z(n23454) );
  XOR U23526 ( .A(n23466), .B(n20712), .Z(n23464) );
  XOR U23527 ( .A(n20719), .B(n20537), .Z(n20712) );
  IV U23528 ( .A(n23461), .Z(n20537) );
  XOR U23529 ( .A(n23473), .B(n23474), .Z(n23461) );
  NANDN U23530 ( .A(n23475), .B(n23476), .Z(n23474) );
  XNOR U23531 ( .A(n23477), .B(n23478), .Z(n20719) );
  OR U23532 ( .A(n23475), .B(n23479), .Z(n23478) );
  ANDN U23533 ( .B(n23480), .A(n23466), .Z(n23471) );
  XNOR U23534 ( .A(n20609), .B(n20707), .Z(n23466) );
  XOR U23535 ( .A(n23473), .B(n23481), .Z(n20707) );
  NANDN U23536 ( .A(n23482), .B(n23483), .Z(n23481) );
  NANDN U23537 ( .A(n23484), .B(n23485), .Z(n23473) );
  OR U23538 ( .A(n23487), .B(n23484), .Z(n23477) );
  XOR U23539 ( .A(n23488), .B(n23475), .Z(n23484) );
  XNOR U23540 ( .A(n23489), .B(n23490), .Z(n23475) );
  XOR U23541 ( .A(n23491), .B(n23483), .Z(n23490) );
  XNOR U23542 ( .A(n23492), .B(n23493), .Z(n23489) );
  XNOR U23543 ( .A(n23494), .B(n23495), .Z(n23493) );
  ANDN U23544 ( .B(n23483), .A(n23496), .Z(n23494) );
  IV U23545 ( .A(n23497), .Z(n23483) );
  ANDN U23546 ( .B(n23488), .A(n23496), .Z(n23486) );
  IV U23547 ( .A(n23482), .Z(n23488) );
  XNOR U23548 ( .A(n23491), .B(n23498), .Z(n23482) );
  XNOR U23549 ( .A(n23495), .B(n23499), .Z(n23498) );
  NANDN U23550 ( .A(n23479), .B(n23476), .Z(n23499) );
  NANDN U23551 ( .A(n23487), .B(n23485), .Z(n23495) );
  XNOR U23552 ( .A(n23476), .B(n23497), .Z(n23485) );
  XOR U23553 ( .A(n23500), .B(n23501), .Z(n23497) );
  XOR U23554 ( .A(n23502), .B(n23503), .Z(n23501) );
  XNOR U23555 ( .A(n23469), .B(n23504), .Z(n23503) );
  XNOR U23556 ( .A(n23505), .B(n23506), .Z(n23500) );
  XNOR U23557 ( .A(n23507), .B(n23508), .Z(n23506) );
  ANDN U23558 ( .B(n23452), .A(n20608), .Z(n23507) );
  XNOR U23559 ( .A(n23496), .B(n23479), .Z(n23487) );
  IV U23560 ( .A(n23492), .Z(n23496) );
  XOR U23561 ( .A(n23509), .B(n23510), .Z(n23492) );
  XNOR U23562 ( .A(n23511), .B(n23504), .Z(n23510) );
  XOR U23563 ( .A(n23512), .B(n23513), .Z(n23504) );
  XNOR U23564 ( .A(n23514), .B(n23515), .Z(n23513) );
  NAND U23565 ( .A(n20713), .B(n23456), .Z(n23515) );
  XNOR U23566 ( .A(n23516), .B(n23517), .Z(n23509) );
  ANDN U23567 ( .B(n23518), .A(n20706), .Z(n23516) );
  XOR U23568 ( .A(n23479), .B(n23476), .Z(n23491) );
  XNOR U23569 ( .A(n23519), .B(n23520), .Z(n23476) );
  XNOR U23570 ( .A(n23512), .B(n23521), .Z(n23520) );
  XNOR U23571 ( .A(n23511), .B(n23452), .Z(n23521) );
  XNOR U23572 ( .A(n23522), .B(n23523), .Z(n23519) );
  XNOR U23573 ( .A(n23524), .B(n23508), .Z(n23523) );
  OR U23574 ( .A(n23470), .B(n20716), .Z(n23508) );
  XNOR U23575 ( .A(n23522), .B(n23505), .Z(n20716) );
  XNOR U23576 ( .A(n23452), .B(n23469), .Z(n23470) );
  ANDN U23577 ( .B(n23469), .A(n20718), .Z(n23524) );
  XOR U23578 ( .A(n23525), .B(n23526), .Z(n23479) );
  XOR U23579 ( .A(n23512), .B(n23502), .Z(n23526) );
  XNOR U23580 ( .A(n23459), .B(n20536), .Z(n23502) );
  XOR U23581 ( .A(n23527), .B(n23514), .Z(n23512) );
  NANDN U23582 ( .A(n23463), .B(n23472), .Z(n23514) );
  XOR U23583 ( .A(n23480), .B(n23456), .Z(n23472) );
  XOR U23584 ( .A(n20536), .B(n23469), .Z(n23456) );
  XNOR U23585 ( .A(n23518), .B(n23528), .Z(n23469) );
  XOR U23586 ( .A(n23529), .B(n23530), .Z(n23528) );
  XNOR U23587 ( .A(n23465), .B(n20713), .Z(n23463) );
  XNOR U23588 ( .A(n20718), .B(n23459), .Z(n20713) );
  IV U23589 ( .A(n23505), .Z(n20718) );
  XOR U23590 ( .A(n23531), .B(n23532), .Z(n23505) );
  XOR U23591 ( .A(n23533), .B(n23534), .Z(n23532) );
  XOR U23592 ( .A(n23522), .B(n23535), .Z(n23531) );
  AND U23593 ( .A(n23480), .B(n23465), .Z(n23527) );
  XOR U23594 ( .A(n20608), .B(n20706), .Z(n23465) );
  IV U23595 ( .A(n23522), .Z(n20608) );
  XOR U23596 ( .A(n23511), .B(n23536), .Z(n23525) );
  XNOR U23597 ( .A(n23537), .B(n23517), .Z(n23536) );
  OR U23598 ( .A(n23447), .B(n23460), .Z(n23517) );
  XNOR U23599 ( .A(n23538), .B(n23459), .Z(n23460) );
  XNOR U23600 ( .A(n23518), .B(n20536), .Z(n23447) );
  AND U23601 ( .A(n20536), .B(n23459), .Z(n23537) );
  XOR U23602 ( .A(n23539), .B(n23540), .Z(n23459) );
  XNOR U23603 ( .A(n23540), .B(n23541), .Z(n20536) );
  XNOR U23604 ( .A(n23530), .B(n23542), .Z(n23541) );
  XNOR U23605 ( .A(n20706), .B(n23448), .Z(n23511) );
  IV U23606 ( .A(n23538), .Z(n20706) );
  XOR U23607 ( .A(n23542), .B(n23543), .Z(n23538) );
  XNOR U23608 ( .A(n23529), .B(n23535), .Z(n23543) );
  XOR U23609 ( .A(n23544), .B(n23545), .Z(n23535) );
  XNOR U23610 ( .A(n18511), .B(n23546), .Z(n23545) );
  XNOR U23611 ( .A(n23530), .B(n19996), .Z(n23546) );
  XNOR U23612 ( .A(n23547), .B(n23548), .Z(n19996) );
  XOR U23613 ( .A(n23549), .B(n23550), .Z(n23548) );
  XNOR U23614 ( .A(n23551), .B(n23552), .Z(n23530) );
  XNOR U23615 ( .A(n18517), .B(n20036), .Z(n23552) );
  XOR U23616 ( .A(n23553), .B(n23554), .Z(n20036) );
  XOR U23617 ( .A(n23555), .B(n23556), .Z(n23554) );
  XNOR U23618 ( .A(n20038), .B(n18508), .Z(n18517) );
  XNOR U23619 ( .A(n23557), .B(n23558), .Z(n18508) );
  XOR U23620 ( .A(n23559), .B(n23560), .Z(n23558) );
  XOR U23621 ( .A(n19409), .B(n23561), .Z(n23551) );
  XNOR U23622 ( .A(key[393]), .B(n19999), .Z(n23561) );
  XOR U23623 ( .A(n18493), .B(n20029), .Z(n18511) );
  XNOR U23624 ( .A(n19420), .B(n23562), .Z(n23544) );
  XOR U23625 ( .A(key[395]), .B(n18469), .Z(n23562) );
  XOR U23626 ( .A(n20040), .B(n18513), .Z(n18469) );
  XNOR U23627 ( .A(n23563), .B(n23564), .Z(n18513) );
  XNOR U23628 ( .A(n23565), .B(n23566), .Z(n23564) );
  XNOR U23629 ( .A(n18516), .B(n19391), .Z(n19420) );
  XNOR U23630 ( .A(n23567), .B(n19409), .Z(n19391) );
  XOR U23631 ( .A(n23568), .B(n23569), .Z(n19409) );
  XOR U23632 ( .A(n23570), .B(n23571), .Z(n23529) );
  XOR U23633 ( .A(n20033), .B(n18510), .Z(n23571) );
  IV U23634 ( .A(n19427), .Z(n20033) );
  XNOR U23635 ( .A(n23572), .B(n23573), .Z(n19427) );
  XNOR U23636 ( .A(n23574), .B(n23575), .Z(n23573) );
  XOR U23637 ( .A(n19997), .B(n23576), .Z(n23570) );
  XOR U23638 ( .A(key[394]), .B(n20040), .Z(n23576) );
  XNOR U23639 ( .A(n23577), .B(n23578), .Z(n20040) );
  XOR U23640 ( .A(n23579), .B(n23580), .Z(n23578) );
  XOR U23641 ( .A(n23581), .B(n23582), .Z(n23577) );
  IV U23642 ( .A(n23539), .Z(n23542) );
  XOR U23643 ( .A(n23518), .B(n23452), .Z(n23480) );
  XNOR U23644 ( .A(n23540), .B(n23583), .Z(n23452) );
  XOR U23645 ( .A(n23539), .B(n23534), .Z(n23583) );
  XNOR U23646 ( .A(n23584), .B(n23585), .Z(n23534) );
  XOR U23647 ( .A(n20027), .B(n18498), .Z(n23585) );
  XNOR U23648 ( .A(n18493), .B(n20014), .Z(n18498) );
  XOR U23649 ( .A(n23586), .B(n19997), .Z(n20027) );
  XOR U23650 ( .A(n23587), .B(n23555), .Z(n19997) );
  XNOR U23651 ( .A(key[396]), .B(n19389), .Z(n23584) );
  XOR U23652 ( .A(n23588), .B(n23589), .Z(n19389) );
  XOR U23653 ( .A(n20015), .B(n18500), .Z(n23589) );
  XNOR U23654 ( .A(n23590), .B(n18471), .Z(n18500) );
  XOR U23655 ( .A(n23591), .B(n23559), .Z(n18471) );
  IV U23656 ( .A(n19400), .Z(n20015) );
  XNOR U23657 ( .A(n23592), .B(n23593), .Z(n19400) );
  XNOR U23658 ( .A(n23567), .B(n23594), .Z(n23593) );
  XNOR U23659 ( .A(n23595), .B(n23596), .Z(n23592) );
  XOR U23660 ( .A(n23597), .B(n23598), .Z(n23596) );
  ANDN U23661 ( .B(n23599), .A(n23600), .Z(n23598) );
  XNOR U23662 ( .A(n23601), .B(n20029), .Z(n23588) );
  XOR U23663 ( .A(n23602), .B(n19999), .Z(n20029) );
  XNOR U23664 ( .A(n23603), .B(n23582), .Z(n19999) );
  IV U23665 ( .A(n23448), .Z(n23518) );
  XOR U23666 ( .A(n23540), .B(n23604), .Z(n23448) );
  XNOR U23667 ( .A(n23539), .B(n23533), .Z(n23604) );
  XOR U23668 ( .A(n23605), .B(n23606), .Z(n23533) );
  XNOR U23669 ( .A(n23547), .B(n23607), .Z(n20006) );
  XNOR U23670 ( .A(n23553), .B(n23608), .Z(n23607) );
  XNOR U23671 ( .A(n23555), .B(n23556), .Z(n23547) );
  XOR U23672 ( .A(n23609), .B(n23610), .Z(n23556) );
  XNOR U23673 ( .A(n23611), .B(n23612), .Z(n23610) );
  NANDN U23674 ( .A(n23613), .B(n23614), .Z(n23612) );
  XNOR U23675 ( .A(n23615), .B(n23616), .Z(n23555) );
  XOR U23676 ( .A(n23617), .B(n23618), .Z(n23616) );
  NANDN U23677 ( .A(n23619), .B(n23620), .Z(n23618) );
  XOR U23678 ( .A(n18493), .B(n23601), .Z(n19430) );
  XNOR U23679 ( .A(key[399]), .B(n19404), .Z(n23605) );
  XOR U23680 ( .A(n20022), .B(n20008), .Z(n19404) );
  XNOR U23681 ( .A(n23563), .B(n23621), .Z(n20008) );
  XNOR U23682 ( .A(n23557), .B(n23622), .Z(n23621) );
  XNOR U23683 ( .A(n23559), .B(n23560), .Z(n23563) );
  XNOR U23684 ( .A(n23623), .B(n23624), .Z(n23560) );
  XNOR U23685 ( .A(n23625), .B(n23626), .Z(n23624) );
  NANDN U23686 ( .A(n23627), .B(n23628), .Z(n23626) );
  XNOR U23687 ( .A(n23629), .B(n23630), .Z(n23559) );
  XOR U23688 ( .A(n23631), .B(n23632), .Z(n23630) );
  NANDN U23689 ( .A(n23633), .B(n23634), .Z(n23632) );
  XOR U23690 ( .A(n23635), .B(n23636), .Z(n23539) );
  XNOR U23691 ( .A(n18481), .B(n19416), .Z(n23636) );
  XNOR U23692 ( .A(n19403), .B(n18486), .Z(n19416) );
  XOR U23693 ( .A(n20011), .B(n18479), .Z(n18486) );
  XOR U23694 ( .A(n23566), .B(n23557), .Z(n18479) );
  XOR U23695 ( .A(n23637), .B(n23565), .Z(n23557) );
  XNOR U23696 ( .A(n23625), .B(n23639), .Z(n23638) );
  NANDN U23697 ( .A(n23640), .B(n23641), .Z(n23639) );
  OR U23698 ( .A(n23642), .B(n23643), .Z(n23625) );
  XOR U23699 ( .A(n23623), .B(n23645), .Z(n23566) );
  XNOR U23700 ( .A(n23646), .B(n23647), .Z(n23645) );
  NOR U23701 ( .A(n23648), .B(n23649), .Z(n23646) );
  XNOR U23702 ( .A(n23644), .B(n23650), .Z(n23623) );
  XNOR U23703 ( .A(n23651), .B(n23652), .Z(n23650) );
  NAND U23704 ( .A(n23653), .B(n23654), .Z(n23652) );
  XOR U23705 ( .A(n18516), .B(n20023), .Z(n19403) );
  XOR U23706 ( .A(n23572), .B(n23655), .Z(n20023) );
  XNOR U23707 ( .A(n23656), .B(n23594), .Z(n23655) );
  XNOR U23708 ( .A(n23657), .B(n23658), .Z(n23594) );
  XNOR U23709 ( .A(n23659), .B(n23660), .Z(n23658) );
  NANDN U23710 ( .A(n23661), .B(n23662), .Z(n23660) );
  XNOR U23711 ( .A(n23663), .B(n23664), .Z(n23572) );
  IV U23712 ( .A(n23601), .Z(n18516) );
  XOR U23713 ( .A(n23569), .B(n23567), .Z(n23601) );
  XNOR U23714 ( .A(n23657), .B(n23665), .Z(n23567) );
  XOR U23715 ( .A(n23666), .B(n23667), .Z(n23665) );
  ANDN U23716 ( .B(n23668), .A(n23669), .Z(n23666) );
  XNOR U23717 ( .A(n23670), .B(n23671), .Z(n23657) );
  XNOR U23718 ( .A(n23672), .B(n23673), .Z(n23671) );
  NANDN U23719 ( .A(n23674), .B(n23675), .Z(n23673) );
  XNOR U23720 ( .A(n18493), .B(n20022), .Z(n18481) );
  XOR U23721 ( .A(n23676), .B(n23677), .Z(n20022) );
  XOR U23722 ( .A(n23579), .B(n23678), .Z(n23677) );
  XNOR U23723 ( .A(n23679), .B(n23582), .Z(n23676) );
  IV U23724 ( .A(n23680), .Z(n23582) );
  XOR U23725 ( .A(n20009), .B(n23681), .Z(n23635) );
  XNOR U23726 ( .A(key[398]), .B(n23522), .Z(n23681) );
  XOR U23727 ( .A(n23682), .B(n23683), .Z(n23522) );
  XNOR U23728 ( .A(n20038), .B(n19425), .Z(n23683) );
  XOR U23729 ( .A(n23656), .B(n23684), .Z(n19425) );
  XOR U23730 ( .A(n23663), .B(n23664), .Z(n23684) );
  XOR U23731 ( .A(n23685), .B(n23686), .Z(n23664) );
  XNOR U23732 ( .A(n23687), .B(n23688), .Z(n23686) );
  NANDN U23733 ( .A(n23689), .B(n23662), .Z(n23688) );
  IV U23734 ( .A(n23568), .Z(n23663) );
  XOR U23735 ( .A(n23670), .B(n23690), .Z(n23568) );
  XNOR U23736 ( .A(n23667), .B(n23691), .Z(n23690) );
  NANDN U23737 ( .A(n23692), .B(n23599), .Z(n23691) );
  XNOR U23738 ( .A(n23579), .B(n23695), .Z(n20038) );
  XNOR U23739 ( .A(n23679), .B(n23680), .Z(n23695) );
  XOR U23740 ( .A(n23696), .B(n23697), .Z(n23680) );
  XOR U23741 ( .A(n23698), .B(n23699), .Z(n23697) );
  NANDN U23742 ( .A(n23700), .B(n23701), .Z(n23699) );
  XNOR U23743 ( .A(n23703), .B(n23704), .Z(n23702) );
  NANDN U23744 ( .A(n23705), .B(n23706), .Z(n23704) );
  XNOR U23745 ( .A(n18493), .B(n23708), .Z(n23682) );
  XNOR U23746 ( .A(key[392]), .B(n18518), .Z(n23708) );
  XNOR U23747 ( .A(n20026), .B(n20007), .Z(n18518) );
  IV U23748 ( .A(n19431), .Z(n20007) );
  XOR U23749 ( .A(n23637), .B(n23590), .Z(n19431) );
  IV U23750 ( .A(n23591), .Z(n23637) );
  XNOR U23751 ( .A(n23629), .B(n23709), .Z(n23591) );
  XOR U23752 ( .A(n23710), .B(n23711), .Z(n23709) );
  ANDN U23753 ( .B(n23641), .A(n23712), .Z(n23710) );
  IV U23754 ( .A(n19405), .Z(n20026) );
  XOR U23755 ( .A(n23713), .B(n23586), .Z(n19405) );
  XNOR U23756 ( .A(n23553), .B(n23550), .Z(n20009) );
  XOR U23757 ( .A(n23609), .B(n23714), .Z(n23550) );
  XNOR U23758 ( .A(n23715), .B(n23716), .Z(n23714) );
  ANDN U23759 ( .B(n23717), .A(n23718), .Z(n23715) );
  XNOR U23760 ( .A(n23719), .B(n23720), .Z(n23609) );
  XNOR U23761 ( .A(n23721), .B(n23722), .Z(n23720) );
  NANDN U23762 ( .A(n23723), .B(n23724), .Z(n23722) );
  XOR U23763 ( .A(n23713), .B(n23549), .Z(n23553) );
  XNOR U23764 ( .A(n23719), .B(n23725), .Z(n23549) );
  XNOR U23765 ( .A(n23611), .B(n23726), .Z(n23725) );
  NANDN U23766 ( .A(n23727), .B(n23728), .Z(n23726) );
  OR U23767 ( .A(n23729), .B(n23730), .Z(n23611) );
  IV U23768 ( .A(n23587), .Z(n23713) );
  XNOR U23769 ( .A(n23615), .B(n23731), .Z(n23587) );
  XOR U23770 ( .A(n23732), .B(n23733), .Z(n23731) );
  ANDN U23771 ( .B(n23728), .A(n23734), .Z(n23732) );
  XNOR U23772 ( .A(n23735), .B(n23736), .Z(n23540) );
  XNOR U23773 ( .A(n19398), .B(n20016), .Z(n23736) );
  XOR U23774 ( .A(n23737), .B(n23738), .Z(n20016) );
  XNOR U23775 ( .A(n23719), .B(n23608), .Z(n23738) );
  XNOR U23776 ( .A(n23739), .B(n23740), .Z(n23608) );
  XNOR U23777 ( .A(n23733), .B(n23741), .Z(n23740) );
  NANDN U23778 ( .A(n23742), .B(n23614), .Z(n23741) );
  OR U23779 ( .A(n23743), .B(n23729), .Z(n23733) );
  XNOR U23780 ( .A(n23614), .B(n23728), .Z(n23729) );
  XOR U23781 ( .A(n23744), .B(n23721), .Z(n23719) );
  NANDN U23782 ( .A(n23745), .B(n23746), .Z(n23721) );
  ANDN U23783 ( .B(n23747), .A(n23748), .Z(n23744) );
  XNOR U23784 ( .A(n23586), .B(n23749), .Z(n23737) );
  XOR U23785 ( .A(n23716), .B(n23750), .Z(n23749) );
  ANDN U23786 ( .B(n23620), .A(n23751), .Z(n23750) );
  NOR U23787 ( .A(n23752), .B(n23753), .Z(n23716) );
  XNOR U23788 ( .A(n23739), .B(n23754), .Z(n23586) );
  XNOR U23789 ( .A(n23755), .B(n23617), .Z(n23754) );
  XNOR U23790 ( .A(n23717), .B(n23620), .Z(n23752) );
  ANDN U23791 ( .B(n23717), .A(n23757), .Z(n23755) );
  XNOR U23792 ( .A(n23615), .B(n23758), .Z(n23739) );
  XNOR U23793 ( .A(n23759), .B(n23760), .Z(n23758) );
  NANDN U23794 ( .A(n23723), .B(n23761), .Z(n23760) );
  XOR U23795 ( .A(n23762), .B(n23759), .Z(n23615) );
  OR U23796 ( .A(n23745), .B(n23763), .Z(n23759) );
  XOR U23797 ( .A(n23764), .B(n23723), .Z(n23745) );
  XNOR U23798 ( .A(n23728), .B(n23620), .Z(n23723) );
  XOR U23799 ( .A(n23765), .B(n23766), .Z(n23620) );
  NANDN U23800 ( .A(n23767), .B(n23768), .Z(n23766) );
  XOR U23801 ( .A(n23769), .B(n23770), .Z(n23728) );
  NANDN U23802 ( .A(n23767), .B(n23771), .Z(n23770) );
  ANDN U23803 ( .B(n23764), .A(n23772), .Z(n23762) );
  IV U23804 ( .A(n23748), .Z(n23764) );
  XNOR U23805 ( .A(n23717), .B(n23614), .Z(n23748) );
  XNOR U23806 ( .A(n23773), .B(n23769), .Z(n23614) );
  NANDN U23807 ( .A(n23774), .B(n23775), .Z(n23769) );
  XOR U23808 ( .A(n23771), .B(n23776), .Z(n23775) );
  ANDN U23809 ( .B(n23776), .A(n23777), .Z(n23773) );
  XNOR U23810 ( .A(n23778), .B(n23765), .Z(n23717) );
  NANDN U23811 ( .A(n23774), .B(n23779), .Z(n23765) );
  XOR U23812 ( .A(n23780), .B(n23768), .Z(n23779) );
  XNOR U23813 ( .A(n23781), .B(n23782), .Z(n23767) );
  XOR U23814 ( .A(n23783), .B(n23784), .Z(n23782) );
  XNOR U23815 ( .A(n23785), .B(n23786), .Z(n23781) );
  XNOR U23816 ( .A(n23787), .B(n23788), .Z(n23786) );
  ANDN U23817 ( .B(n23780), .A(n23784), .Z(n23787) );
  ANDN U23818 ( .B(n23780), .A(n23777), .Z(n23778) );
  XNOR U23819 ( .A(n23783), .B(n23789), .Z(n23777) );
  XOR U23820 ( .A(n23790), .B(n23788), .Z(n23789) );
  NAND U23821 ( .A(n23791), .B(n23792), .Z(n23788) );
  XNOR U23822 ( .A(n23785), .B(n23768), .Z(n23792) );
  IV U23823 ( .A(n23780), .Z(n23785) );
  XNOR U23824 ( .A(n23771), .B(n23784), .Z(n23791) );
  IV U23825 ( .A(n23776), .Z(n23784) );
  XOR U23826 ( .A(n23793), .B(n23794), .Z(n23776) );
  XNOR U23827 ( .A(n23795), .B(n23796), .Z(n23794) );
  XNOR U23828 ( .A(n23797), .B(n23798), .Z(n23793) );
  NOR U23829 ( .A(n23718), .B(n23757), .Z(n23797) );
  AND U23830 ( .A(n23768), .B(n23771), .Z(n23790) );
  XNOR U23831 ( .A(n23768), .B(n23771), .Z(n23783) );
  XNOR U23832 ( .A(n23799), .B(n23800), .Z(n23771) );
  XNOR U23833 ( .A(n23801), .B(n23796), .Z(n23800) );
  XOR U23834 ( .A(n23802), .B(n23803), .Z(n23799) );
  XNOR U23835 ( .A(n23804), .B(n23798), .Z(n23803) );
  OR U23836 ( .A(n23753), .B(n23756), .Z(n23798) );
  XNOR U23837 ( .A(n23757), .B(n23619), .Z(n23756) );
  XNOR U23838 ( .A(n23718), .B(n23751), .Z(n23753) );
  ANDN U23839 ( .B(n23805), .A(n23619), .Z(n23804) );
  XNOR U23840 ( .A(n23806), .B(n23807), .Z(n23768) );
  XNOR U23841 ( .A(n23796), .B(n23808), .Z(n23807) );
  XOR U23842 ( .A(n23613), .B(n23802), .Z(n23808) );
  XNOR U23843 ( .A(n23757), .B(n23809), .Z(n23796) );
  XOR U23844 ( .A(n23742), .B(n23810), .Z(n23806) );
  XNOR U23845 ( .A(n23811), .B(n23812), .Z(n23810) );
  ANDN U23846 ( .B(n23813), .A(n23734), .Z(n23811) );
  XNOR U23847 ( .A(n23814), .B(n23815), .Z(n23780) );
  XNOR U23848 ( .A(n23801), .B(n23816), .Z(n23815) );
  XNOR U23849 ( .A(n23727), .B(n23795), .Z(n23816) );
  XOR U23850 ( .A(n23802), .B(n23817), .Z(n23795) );
  XNOR U23851 ( .A(n23818), .B(n23819), .Z(n23817) );
  NAND U23852 ( .A(n23761), .B(n23724), .Z(n23819) );
  XNOR U23853 ( .A(n23820), .B(n23818), .Z(n23802) );
  NANDN U23854 ( .A(n23763), .B(n23746), .Z(n23818) );
  XOR U23855 ( .A(n23747), .B(n23724), .Z(n23746) );
  XNOR U23856 ( .A(n23813), .B(n23751), .Z(n23724) );
  XOR U23857 ( .A(n23772), .B(n23761), .Z(n23763) );
  XNOR U23858 ( .A(n23734), .B(n23821), .Z(n23761) );
  ANDN U23859 ( .B(n23747), .A(n23772), .Z(n23820) );
  XNOR U23860 ( .A(n23742), .B(n23757), .Z(n23772) );
  XOR U23861 ( .A(n23822), .B(n23823), .Z(n23757) );
  XNOR U23862 ( .A(n23824), .B(n23825), .Z(n23823) );
  XOR U23863 ( .A(n23821), .B(n23805), .Z(n23801) );
  IV U23864 ( .A(n23751), .Z(n23805) );
  XOR U23865 ( .A(n23826), .B(n23827), .Z(n23751) );
  XNOR U23866 ( .A(n23828), .B(n23825), .Z(n23827) );
  IV U23867 ( .A(n23619), .Z(n23821) );
  XOR U23868 ( .A(n23825), .B(n23829), .Z(n23619) );
  XNOR U23869 ( .A(n23830), .B(n23831), .Z(n23814) );
  XNOR U23870 ( .A(n23832), .B(n23812), .Z(n23831) );
  OR U23871 ( .A(n23730), .B(n23743), .Z(n23812) );
  XNOR U23872 ( .A(n23742), .B(n23734), .Z(n23743) );
  IV U23873 ( .A(n23830), .Z(n23734) );
  XOR U23874 ( .A(n23613), .B(n23813), .Z(n23730) );
  IV U23875 ( .A(n23727), .Z(n23813) );
  XOR U23876 ( .A(n23809), .B(n23833), .Z(n23727) );
  XNOR U23877 ( .A(n23828), .B(n23822), .Z(n23833) );
  XOR U23878 ( .A(n23834), .B(n23835), .Z(n23822) );
  XOR U23879 ( .A(n22372), .B(n21398), .Z(n23835) );
  XOR U23880 ( .A(n21388), .B(n22376), .Z(n21398) );
  XOR U23881 ( .A(n21401), .B(n21384), .Z(n22372) );
  XOR U23882 ( .A(n23836), .B(n23837), .Z(n21384) );
  XOR U23883 ( .A(n23838), .B(n23839), .Z(n23837) );
  XOR U23884 ( .A(n23840), .B(n23841), .Z(n23836) );
  XNOR U23885 ( .A(key[370]), .B(n21389), .Z(n23834) );
  IV U23886 ( .A(n23718), .Z(n23809) );
  XOR U23887 ( .A(n23826), .B(n23842), .Z(n23718) );
  XOR U23888 ( .A(n23825), .B(n23843), .Z(n23842) );
  NOR U23889 ( .A(n23613), .B(n23742), .Z(n23832) );
  XOR U23890 ( .A(n23826), .B(n23844), .Z(n23613) );
  XOR U23891 ( .A(n23825), .B(n23845), .Z(n23844) );
  XOR U23892 ( .A(n23846), .B(n23847), .Z(n23825) );
  XNOR U23893 ( .A(n22401), .B(n21379), .Z(n23847) );
  XNOR U23894 ( .A(n23143), .B(n23848), .Z(n21379) );
  XNOR U23895 ( .A(n21363), .B(n23163), .Z(n23143) );
  IV U23896 ( .A(n22407), .Z(n23163) );
  XNOR U23897 ( .A(n23849), .B(n23850), .Z(n22407) );
  XNOR U23898 ( .A(n23851), .B(n23852), .Z(n21363) );
  XOR U23899 ( .A(n22397), .B(n21356), .Z(n22401) );
  XNOR U23900 ( .A(n23853), .B(n23854), .Z(n21356) );
  XNOR U23901 ( .A(n23855), .B(n23856), .Z(n23854) );
  XNOR U23902 ( .A(n23840), .B(n23857), .Z(n23853) );
  XOR U23903 ( .A(n21365), .B(n23858), .Z(n23846) );
  XOR U23904 ( .A(key[374]), .B(n23742), .Z(n23858) );
  IV U23905 ( .A(n23829), .Z(n23826) );
  XOR U23906 ( .A(n23859), .B(n23860), .Z(n23829) );
  XNOR U23907 ( .A(n23157), .B(n21362), .Z(n23860) );
  XOR U23908 ( .A(n23126), .B(n22404), .Z(n21362) );
  XNOR U23909 ( .A(n23861), .B(n23862), .Z(n22404) );
  XNOR U23910 ( .A(n23863), .B(n23864), .Z(n23862) );
  XOR U23911 ( .A(n23865), .B(n23866), .Z(n23861) );
  XOR U23912 ( .A(n23867), .B(n23868), .Z(n23866) );
  ANDN U23913 ( .B(n23869), .A(n23870), .Z(n23868) );
  XOR U23914 ( .A(n23871), .B(n23872), .Z(n23126) );
  XNOR U23915 ( .A(n23873), .B(n23874), .Z(n23872) );
  XNOR U23916 ( .A(n23875), .B(n23876), .Z(n23871) );
  XNOR U23917 ( .A(n23877), .B(n23878), .Z(n23876) );
  ANDN U23918 ( .B(n23879), .A(n23880), .Z(n23878) );
  XNOR U23919 ( .A(n21365), .B(n21377), .Z(n23157) );
  XOR U23920 ( .A(n23855), .B(n23839), .Z(n21377) );
  XNOR U23921 ( .A(n23881), .B(n23882), .Z(n23839) );
  XNOR U23922 ( .A(n23883), .B(n23884), .Z(n23882) );
  NOR U23923 ( .A(n23885), .B(n23886), .Z(n23883) );
  XNOR U23924 ( .A(n23887), .B(n23888), .Z(n21365) );
  XOR U23925 ( .A(key[373]), .B(n23142), .Z(n23859) );
  XOR U23926 ( .A(n23889), .B(n23890), .Z(n23830) );
  XNOR U23927 ( .A(n23845), .B(n23843), .Z(n23890) );
  XNOR U23928 ( .A(n23891), .B(n23892), .Z(n23843) );
  XNOR U23929 ( .A(n23848), .B(n21357), .Z(n23892) );
  XOR U23930 ( .A(n23893), .B(n23894), .Z(n22385) );
  XNOR U23931 ( .A(n23895), .B(n23864), .Z(n23894) );
  XNOR U23932 ( .A(n23896), .B(n23897), .Z(n23864) );
  XNOR U23933 ( .A(n23898), .B(n23899), .Z(n23897) );
  NANDN U23934 ( .A(n23900), .B(n23901), .Z(n23899) );
  XOR U23935 ( .A(n23902), .B(n23851), .Z(n23893) );
  XOR U23936 ( .A(n23903), .B(n23904), .Z(n23158) );
  XNOR U23937 ( .A(n23849), .B(n23874), .Z(n23904) );
  XNOR U23938 ( .A(n23905), .B(n23906), .Z(n23874) );
  XNOR U23939 ( .A(n23907), .B(n23908), .Z(n23906) );
  OR U23940 ( .A(n23909), .B(n23910), .Z(n23908) );
  XOR U23941 ( .A(n23161), .B(n23139), .Z(n23848) );
  XNOR U23942 ( .A(n23911), .B(n23912), .Z(n23139) );
  XNOR U23943 ( .A(n23913), .B(n23914), .Z(n23912) );
  XOR U23944 ( .A(n23915), .B(n23887), .Z(n23911) );
  XNOR U23945 ( .A(key[375]), .B(n22397), .Z(n23891) );
  XNOR U23946 ( .A(n23916), .B(n23917), .Z(n23845) );
  XNOR U23947 ( .A(n21345), .B(n21343), .Z(n23917) );
  XOR U23948 ( .A(n23128), .B(n22389), .Z(n21343) );
  XNOR U23949 ( .A(n23918), .B(n21388), .Z(n22389) );
  XOR U23950 ( .A(n23921), .B(n23922), .Z(n22376) );
  XOR U23951 ( .A(n23161), .B(n23142), .Z(n21345) );
  XNOR U23952 ( .A(n23923), .B(n23924), .Z(n23142) );
  XNOR U23953 ( .A(n23925), .B(n23914), .Z(n23924) );
  XNOR U23954 ( .A(n23926), .B(n23927), .Z(n23914) );
  XNOR U23955 ( .A(n23928), .B(n23929), .Z(n23927) );
  NANDN U23956 ( .A(n23930), .B(n23931), .Z(n23929) );
  XNOR U23957 ( .A(n23932), .B(n23933), .Z(n23923) );
  XOR U23958 ( .A(n23934), .B(n23935), .Z(n23933) );
  ANDN U23959 ( .B(n23936), .A(n23937), .Z(n23935) );
  XNOR U23960 ( .A(n22391), .B(n23938), .Z(n23916) );
  XOR U23961 ( .A(key[372]), .B(n23124), .Z(n23938) );
  XNOR U23962 ( .A(n22397), .B(n21361), .Z(n22391) );
  XOR U23963 ( .A(n23939), .B(n23940), .Z(n21361) );
  XNOR U23964 ( .A(n23941), .B(n23856), .Z(n23940) );
  XNOR U23965 ( .A(n23942), .B(n23943), .Z(n23856) );
  XNOR U23966 ( .A(n23944), .B(n23945), .Z(n23943) );
  NANDN U23967 ( .A(n23946), .B(n23947), .Z(n23945) );
  XNOR U23968 ( .A(n23948), .B(n23949), .Z(n23939) );
  XOR U23969 ( .A(n23884), .B(n23950), .Z(n23949) );
  ANDN U23970 ( .B(n23951), .A(n23952), .Z(n23950) );
  ANDN U23971 ( .B(n23953), .A(n23954), .Z(n23884) );
  XNOR U23972 ( .A(n23742), .B(n23824), .Z(n23889) );
  XOR U23973 ( .A(n23955), .B(n23956), .Z(n23824) );
  XNOR U23974 ( .A(n21392), .B(n23957), .Z(n23956) );
  XNOR U23975 ( .A(n23828), .B(n21394), .Z(n23957) );
  XOR U23976 ( .A(n23161), .B(n23124), .Z(n21394) );
  XOR U23977 ( .A(n23932), .B(n21389), .Z(n23124) );
  IV U23978 ( .A(n23958), .Z(n21389) );
  XOR U23979 ( .A(n23959), .B(n23960), .Z(n23828) );
  XNOR U23980 ( .A(n22363), .B(n21387), .Z(n23960) );
  XOR U23981 ( .A(n22398), .B(n21372), .Z(n21387) );
  XNOR U23982 ( .A(n23919), .B(n23961), .Z(n21372) );
  XNOR U23983 ( .A(n23902), .B(n23851), .Z(n23961) );
  XOR U23984 ( .A(n23920), .B(n23962), .Z(n23851) );
  XOR U23985 ( .A(n23849), .B(n23963), .Z(n22398) );
  XNOR U23986 ( .A(n23922), .B(n23964), .Z(n23963) );
  XNOR U23987 ( .A(n23921), .B(n23965), .Z(n23849) );
  IV U23988 ( .A(n23966), .Z(n23921) );
  XOR U23989 ( .A(n21399), .B(n23958), .Z(n22363) );
  XOR U23990 ( .A(n23967), .B(n23913), .Z(n23958) );
  XNOR U23991 ( .A(key[369]), .B(n21374), .Z(n23959) );
  XOR U23992 ( .A(n22361), .B(n21397), .Z(n21392) );
  XNOR U23993 ( .A(n23968), .B(n23969), .Z(n21397) );
  XNOR U23994 ( .A(n23895), .B(n23852), .Z(n23969) );
  XNOR U23995 ( .A(n23970), .B(n23971), .Z(n23852) );
  XNOR U23996 ( .A(n23972), .B(n23867), .Z(n23971) );
  ANDN U23997 ( .B(n23973), .A(n23974), .Z(n23867) );
  NOR U23998 ( .A(n23975), .B(n23976), .Z(n23972) );
  IV U23999 ( .A(n23919), .Z(n23895) );
  XOR U24000 ( .A(n23977), .B(n23978), .Z(n23919) );
  XOR U24001 ( .A(n23979), .B(n23980), .Z(n23978) );
  NANDN U24002 ( .A(n23981), .B(n23869), .Z(n23980) );
  XOR U24003 ( .A(n23902), .B(n23962), .Z(n23968) );
  XOR U24004 ( .A(n23863), .B(n23982), .Z(n23962) );
  XNOR U24005 ( .A(n23983), .B(n23984), .Z(n23982) );
  NANDN U24006 ( .A(n23985), .B(n23986), .Z(n23984) );
  XNOR U24007 ( .A(n23983), .B(n23988), .Z(n23987) );
  NANDN U24008 ( .A(n23989), .B(n23901), .Z(n23988) );
  OR U24009 ( .A(n23990), .B(n23991), .Z(n23983) );
  XNOR U24010 ( .A(n23863), .B(n23992), .Z(n23970) );
  XNOR U24011 ( .A(n23993), .B(n23994), .Z(n23992) );
  NAND U24012 ( .A(n23995), .B(n23996), .Z(n23994) );
  XOR U24013 ( .A(n23997), .B(n23993), .Z(n23863) );
  NANDN U24014 ( .A(n23998), .B(n23999), .Z(n23993) );
  ANDN U24015 ( .B(n24000), .A(n24001), .Z(n23997) );
  IV U24016 ( .A(n23152), .Z(n22361) );
  XNOR U24017 ( .A(n23903), .B(n24002), .Z(n23152) );
  XOR U24018 ( .A(n23965), .B(n23850), .Z(n24002) );
  XNOR U24019 ( .A(n24003), .B(n24004), .Z(n23850) );
  XOR U24020 ( .A(n24005), .B(n23877), .Z(n24004) );
  NANDN U24021 ( .A(n24006), .B(n24007), .Z(n23877) );
  NOR U24022 ( .A(n24008), .B(n24009), .Z(n24005) );
  XOR U24023 ( .A(n23873), .B(n24010), .Z(n23965) );
  XNOR U24024 ( .A(n24011), .B(n24012), .Z(n24010) );
  NANDN U24025 ( .A(n24013), .B(n24014), .Z(n24012) );
  XOR U24026 ( .A(n23922), .B(n23964), .Z(n23903) );
  XOR U24027 ( .A(n24003), .B(n24015), .Z(n23964) );
  XNOR U24028 ( .A(n24011), .B(n24016), .Z(n24015) );
  OR U24029 ( .A(n23909), .B(n24017), .Z(n24016) );
  OR U24030 ( .A(n24018), .B(n24019), .Z(n24011) );
  XNOR U24031 ( .A(n23873), .B(n24020), .Z(n24003) );
  XNOR U24032 ( .A(n24021), .B(n24022), .Z(n24020) );
  NAND U24033 ( .A(n24023), .B(n24024), .Z(n24022) );
  XOR U24034 ( .A(n24025), .B(n24021), .Z(n23873) );
  NANDN U24035 ( .A(n24026), .B(n24027), .Z(n24021) );
  AND U24036 ( .A(n24028), .B(n24029), .Z(n24025) );
  XOR U24037 ( .A(n24030), .B(n24031), .Z(n23922) );
  XNOR U24038 ( .A(n24032), .B(n24033), .Z(n24031) );
  NAND U24039 ( .A(n24034), .B(n23879), .Z(n24033) );
  XNOR U24040 ( .A(n22380), .B(n24035), .Z(n23955) );
  XNOR U24041 ( .A(key[371]), .B(n21401), .Z(n24035) );
  XOR U24042 ( .A(n24036), .B(n24037), .Z(n21401) );
  XNOR U24043 ( .A(n23913), .B(n23888), .Z(n24037) );
  XNOR U24044 ( .A(n24038), .B(n24039), .Z(n23888) );
  XNOR U24045 ( .A(n24040), .B(n23934), .Z(n24039) );
  ANDN U24046 ( .B(n24041), .A(n24042), .Z(n23934) );
  NOR U24047 ( .A(n24043), .B(n24044), .Z(n24040) );
  IV U24048 ( .A(n24045), .Z(n23913) );
  XNOR U24049 ( .A(n23915), .B(n24046), .Z(n24036) );
  XNOR U24050 ( .A(n22397), .B(n21347), .Z(n22380) );
  XOR U24051 ( .A(n23941), .B(n21399), .Z(n21347) );
  XNOR U24052 ( .A(n23840), .B(n24047), .Z(n21399) );
  XOR U24053 ( .A(n24047), .B(n23941), .Z(n22397) );
  XNOR U24054 ( .A(n23942), .B(n24048), .Z(n23941) );
  XOR U24055 ( .A(n24049), .B(n24050), .Z(n24048) );
  ANDN U24056 ( .B(n24051), .A(n23886), .Z(n24049) );
  XOR U24057 ( .A(n24052), .B(n24053), .Z(n23942) );
  XNOR U24058 ( .A(n24054), .B(n24055), .Z(n24053) );
  NAND U24059 ( .A(n24056), .B(n24057), .Z(n24055) );
  XNOR U24060 ( .A(n24058), .B(n24059), .Z(n23742) );
  XOR U24061 ( .A(n23148), .B(n22378), .Z(n24059) );
  XNOR U24062 ( .A(n21391), .B(n21374), .Z(n22378) );
  XOR U24063 ( .A(n24045), .B(n24060), .Z(n21374) );
  XNOR U24064 ( .A(n23915), .B(n23887), .Z(n24060) );
  XOR U24065 ( .A(n23967), .B(n24046), .Z(n23887) );
  XNOR U24066 ( .A(n23925), .B(n24061), .Z(n24046) );
  XNOR U24067 ( .A(n24062), .B(n24063), .Z(n24061) );
  NANDN U24068 ( .A(n24064), .B(n24065), .Z(n24063) );
  XNOR U24069 ( .A(n24062), .B(n24067), .Z(n24066) );
  NANDN U24070 ( .A(n24068), .B(n23931), .Z(n24067) );
  OR U24071 ( .A(n24069), .B(n24070), .Z(n24062) );
  XNOR U24072 ( .A(n23925), .B(n24071), .Z(n24038) );
  XNOR U24073 ( .A(n24072), .B(n24073), .Z(n24071) );
  NAND U24074 ( .A(n24074), .B(n24075), .Z(n24073) );
  XOR U24075 ( .A(n24076), .B(n24072), .Z(n23925) );
  NANDN U24076 ( .A(n24077), .B(n24078), .Z(n24072) );
  ANDN U24077 ( .B(n24079), .A(n24080), .Z(n24076) );
  XOR U24078 ( .A(n24081), .B(n24082), .Z(n24045) );
  XOR U24079 ( .A(n24083), .B(n24084), .Z(n24082) );
  NANDN U24080 ( .A(n24085), .B(n23936), .Z(n24084) );
  XNOR U24081 ( .A(n23840), .B(n23841), .Z(n24086) );
  IV U24082 ( .A(n23857), .Z(n23841) );
  XOR U24083 ( .A(n23881), .B(n24087), .Z(n23857) );
  XNOR U24084 ( .A(n24088), .B(n24089), .Z(n24087) );
  NANDN U24085 ( .A(n24090), .B(n23947), .Z(n24089) );
  XNOR U24086 ( .A(n23948), .B(n24091), .Z(n23881) );
  XNOR U24087 ( .A(n24092), .B(n24093), .Z(n24091) );
  NAND U24088 ( .A(n24094), .B(n24056), .Z(n24093) );
  XNOR U24089 ( .A(n24050), .B(n24096), .Z(n24095) );
  NANDN U24090 ( .A(n24097), .B(n23951), .Z(n24096) );
  XNOR U24091 ( .A(n23886), .B(n23951), .Z(n23953) );
  XNOR U24092 ( .A(n24047), .B(n23838), .Z(n23855) );
  XOR U24093 ( .A(n23948), .B(n24099), .Z(n23838) );
  XNOR U24094 ( .A(n24088), .B(n24100), .Z(n24099) );
  NANDN U24095 ( .A(n24101), .B(n24102), .Z(n24100) );
  OR U24096 ( .A(n24103), .B(n24104), .Z(n24088) );
  XOR U24097 ( .A(n24105), .B(n24092), .Z(n23948) );
  NANDN U24098 ( .A(n24106), .B(n24107), .Z(n24092) );
  ANDN U24099 ( .B(n24108), .A(n24109), .Z(n24105) );
  XNOR U24100 ( .A(n24052), .B(n24110), .Z(n24047) );
  XOR U24101 ( .A(n24111), .B(n23944), .Z(n24110) );
  OR U24102 ( .A(n24112), .B(n24103), .Z(n23944) );
  XNOR U24103 ( .A(n23947), .B(n24102), .Z(n24103) );
  ANDN U24104 ( .B(n24102), .A(n24113), .Z(n24111) );
  XNOR U24105 ( .A(n24114), .B(n24054), .Z(n24052) );
  OR U24106 ( .A(n24106), .B(n24115), .Z(n24054) );
  XNOR U24107 ( .A(n24116), .B(n24056), .Z(n24106) );
  XOR U24108 ( .A(n24102), .B(n23951), .Z(n24056) );
  XOR U24109 ( .A(n24117), .B(n24118), .Z(n23951) );
  NANDN U24110 ( .A(n24119), .B(n24120), .Z(n24118) );
  XOR U24111 ( .A(n24121), .B(n24122), .Z(n24102) );
  NANDN U24112 ( .A(n24119), .B(n24123), .Z(n24122) );
  ANDN U24113 ( .B(n24116), .A(n24124), .Z(n24114) );
  IV U24114 ( .A(n24109), .Z(n24116) );
  XOR U24115 ( .A(n23886), .B(n23947), .Z(n24109) );
  XNOR U24116 ( .A(n24125), .B(n24121), .Z(n23947) );
  NANDN U24117 ( .A(n24126), .B(n24127), .Z(n24121) );
  XOR U24118 ( .A(n24123), .B(n24128), .Z(n24127) );
  ANDN U24119 ( .B(n24128), .A(n24129), .Z(n24125) );
  XOR U24120 ( .A(n24130), .B(n24117), .Z(n23886) );
  NANDN U24121 ( .A(n24126), .B(n24131), .Z(n24117) );
  XOR U24122 ( .A(n24132), .B(n24120), .Z(n24131) );
  XNOR U24123 ( .A(n24133), .B(n24134), .Z(n24119) );
  XOR U24124 ( .A(n24135), .B(n24136), .Z(n24134) );
  XNOR U24125 ( .A(n24137), .B(n24138), .Z(n24133) );
  XNOR U24126 ( .A(n24139), .B(n24140), .Z(n24138) );
  ANDN U24127 ( .B(n24132), .A(n24136), .Z(n24139) );
  ANDN U24128 ( .B(n24132), .A(n24129), .Z(n24130) );
  XNOR U24129 ( .A(n24135), .B(n24141), .Z(n24129) );
  XOR U24130 ( .A(n24142), .B(n24140), .Z(n24141) );
  NAND U24131 ( .A(n24143), .B(n24144), .Z(n24140) );
  XNOR U24132 ( .A(n24137), .B(n24120), .Z(n24144) );
  IV U24133 ( .A(n24132), .Z(n24137) );
  XNOR U24134 ( .A(n24123), .B(n24136), .Z(n24143) );
  IV U24135 ( .A(n24128), .Z(n24136) );
  XOR U24136 ( .A(n24145), .B(n24146), .Z(n24128) );
  XNOR U24137 ( .A(n24147), .B(n24148), .Z(n24146) );
  XNOR U24138 ( .A(n24149), .B(n24150), .Z(n24145) );
  ANDN U24139 ( .B(n24051), .A(n23885), .Z(n24149) );
  AND U24140 ( .A(n24120), .B(n24123), .Z(n24142) );
  XNOR U24141 ( .A(n24120), .B(n24123), .Z(n24135) );
  XNOR U24142 ( .A(n24151), .B(n24152), .Z(n24123) );
  XNOR U24143 ( .A(n24153), .B(n24148), .Z(n24152) );
  XOR U24144 ( .A(n24154), .B(n24155), .Z(n24151) );
  XNOR U24145 ( .A(n24156), .B(n24150), .Z(n24155) );
  OR U24146 ( .A(n23954), .B(n24098), .Z(n24150) );
  XNOR U24147 ( .A(n24051), .B(n24157), .Z(n24098) );
  XNOR U24148 ( .A(n23885), .B(n23952), .Z(n23954) );
  ANDN U24149 ( .B(n24158), .A(n24097), .Z(n24156) );
  XNOR U24150 ( .A(n24159), .B(n24160), .Z(n24120) );
  XNOR U24151 ( .A(n24148), .B(n24161), .Z(n24160) );
  XOR U24152 ( .A(n24090), .B(n24154), .Z(n24161) );
  XNOR U24153 ( .A(n24051), .B(n23885), .Z(n24148) );
  XOR U24154 ( .A(n23946), .B(n24162), .Z(n24159) );
  XNOR U24155 ( .A(n24163), .B(n24164), .Z(n24162) );
  ANDN U24156 ( .B(n24165), .A(n24113), .Z(n24163) );
  XNOR U24157 ( .A(n24166), .B(n24167), .Z(n24132) );
  XNOR U24158 ( .A(n24153), .B(n24168), .Z(n24167) );
  XNOR U24159 ( .A(n24101), .B(n24147), .Z(n24168) );
  XOR U24160 ( .A(n24154), .B(n24169), .Z(n24147) );
  XNOR U24161 ( .A(n24170), .B(n24171), .Z(n24169) );
  NAND U24162 ( .A(n24057), .B(n24094), .Z(n24171) );
  XNOR U24163 ( .A(n24172), .B(n24170), .Z(n24154) );
  NANDN U24164 ( .A(n24115), .B(n24107), .Z(n24170) );
  XOR U24165 ( .A(n24108), .B(n24094), .Z(n24107) );
  XNOR U24166 ( .A(n24165), .B(n23952), .Z(n24094) );
  XOR U24167 ( .A(n24124), .B(n24057), .Z(n24115) );
  XNOR U24168 ( .A(n24113), .B(n24157), .Z(n24057) );
  ANDN U24169 ( .B(n24108), .A(n24124), .Z(n24172) );
  XOR U24170 ( .A(n23946), .B(n24051), .Z(n24124) );
  XNOR U24171 ( .A(n24173), .B(n24174), .Z(n24051) );
  XNOR U24172 ( .A(n24175), .B(n24176), .Z(n24174) );
  XOR U24173 ( .A(n24157), .B(n24158), .Z(n24153) );
  IV U24174 ( .A(n23952), .Z(n24158) );
  XOR U24175 ( .A(n24177), .B(n24178), .Z(n23952) );
  XNOR U24176 ( .A(n24179), .B(n24176), .Z(n24178) );
  IV U24177 ( .A(n24097), .Z(n24157) );
  XOR U24178 ( .A(n24176), .B(n24180), .Z(n24097) );
  XNOR U24179 ( .A(n24181), .B(n24182), .Z(n24166) );
  XNOR U24180 ( .A(n24183), .B(n24164), .Z(n24182) );
  OR U24181 ( .A(n24104), .B(n24112), .Z(n24164) );
  XNOR U24182 ( .A(n23946), .B(n24113), .Z(n24112) );
  IV U24183 ( .A(n24181), .Z(n24113) );
  XOR U24184 ( .A(n24090), .B(n24165), .Z(n24104) );
  IV U24185 ( .A(n24101), .Z(n24165) );
  XNOR U24186 ( .A(n24179), .B(n24173), .Z(n24184) );
  XOR U24187 ( .A(n24185), .B(n24186), .Z(n24173) );
  XNOR U24188 ( .A(n24187), .B(n24188), .Z(n24186) );
  XOR U24189 ( .A(key[210]), .B(n24189), .Z(n24185) );
  XOR U24190 ( .A(n24177), .B(n24190), .Z(n23885) );
  XOR U24191 ( .A(n24176), .B(n24191), .Z(n24190) );
  NOR U24192 ( .A(n24090), .B(n23946), .Z(n24183) );
  XOR U24193 ( .A(n24177), .B(n24192), .Z(n24090) );
  XOR U24194 ( .A(n24176), .B(n24193), .Z(n24192) );
  XOR U24195 ( .A(n24194), .B(n24195), .Z(n24176) );
  XNOR U24196 ( .A(n24196), .B(n24197), .Z(n24195) );
  XNOR U24197 ( .A(n24198), .B(n24199), .Z(n24194) );
  XOR U24198 ( .A(key[214]), .B(n23946), .Z(n24199) );
  IV U24199 ( .A(n24180), .Z(n24177) );
  XOR U24200 ( .A(n24200), .B(n24201), .Z(n24180) );
  XNOR U24201 ( .A(n24202), .B(n24203), .Z(n24201) );
  XNOR U24202 ( .A(key[213]), .B(n24204), .Z(n24200) );
  XOR U24203 ( .A(n24205), .B(n24206), .Z(n24181) );
  XNOR U24204 ( .A(n24193), .B(n24191), .Z(n24206) );
  XNOR U24205 ( .A(n24207), .B(n24208), .Z(n24191) );
  XNOR U24206 ( .A(n24209), .B(n24210), .Z(n24208) );
  XNOR U24207 ( .A(key[215]), .B(n24211), .Z(n24207) );
  XNOR U24208 ( .A(n24212), .B(n24213), .Z(n24193) );
  XOR U24209 ( .A(n24214), .B(n24215), .Z(n24213) );
  XNOR U24210 ( .A(n24216), .B(n24217), .Z(n24212) );
  XNOR U24211 ( .A(key[212]), .B(n24218), .Z(n24217) );
  XNOR U24212 ( .A(n23946), .B(n24175), .Z(n24205) );
  XOR U24213 ( .A(n24219), .B(n24220), .Z(n24175) );
  XNOR U24214 ( .A(n24221), .B(n24222), .Z(n24220) );
  XNOR U24215 ( .A(n24179), .B(n24223), .Z(n24222) );
  XOR U24216 ( .A(n24224), .B(n24225), .Z(n24179) );
  XNOR U24217 ( .A(n24226), .B(n24227), .Z(n24225) );
  XOR U24218 ( .A(key[209]), .B(n24228), .Z(n24224) );
  XOR U24219 ( .A(n24229), .B(n24230), .Z(n24219) );
  XNOR U24220 ( .A(key[211]), .B(n24231), .Z(n24230) );
  XNOR U24221 ( .A(n24232), .B(n24233), .Z(n23946) );
  XNOR U24222 ( .A(key[208]), .B(n24236), .Z(n24232) );
  IV U24223 ( .A(n23125), .Z(n23148) );
  XOR U24224 ( .A(n23966), .B(n23875), .Z(n23125) );
  XNOR U24225 ( .A(n23905), .B(n24237), .Z(n23875) );
  XOR U24226 ( .A(n24238), .B(n24032), .Z(n24237) );
  NANDN U24227 ( .A(n24239), .B(n24007), .Z(n24032) );
  XNOR U24228 ( .A(n24009), .B(n23879), .Z(n24007) );
  NOR U24229 ( .A(n24240), .B(n24009), .Z(n24238) );
  XNOR U24230 ( .A(n24030), .B(n24241), .Z(n23905) );
  XNOR U24231 ( .A(n24242), .B(n24243), .Z(n24241) );
  NAND U24232 ( .A(n24024), .B(n24244), .Z(n24243) );
  XNOR U24233 ( .A(n24030), .B(n24245), .Z(n23966) );
  XOR U24234 ( .A(n24246), .B(n23907), .Z(n24245) );
  OR U24235 ( .A(n24247), .B(n24018), .Z(n23907) );
  XNOR U24236 ( .A(n23909), .B(n24013), .Z(n24018) );
  NOR U24237 ( .A(n24248), .B(n24013), .Z(n24246) );
  XOR U24238 ( .A(n24249), .B(n24242), .Z(n24030) );
  OR U24239 ( .A(n24026), .B(n24250), .Z(n24242) );
  XNOR U24240 ( .A(n24028), .B(n24024), .Z(n24026) );
  XNOR U24241 ( .A(n24013), .B(n23879), .Z(n24024) );
  XOR U24242 ( .A(n24251), .B(n24252), .Z(n23879) );
  NANDN U24243 ( .A(n24253), .B(n24254), .Z(n24252) );
  XNOR U24244 ( .A(n24255), .B(n24256), .Z(n24013) );
  OR U24245 ( .A(n24253), .B(n24257), .Z(n24256) );
  ANDN U24246 ( .B(n24028), .A(n24258), .Z(n24249) );
  XOR U24247 ( .A(n23909), .B(n24009), .Z(n24028) );
  XOR U24248 ( .A(n24259), .B(n24251), .Z(n24009) );
  NANDN U24249 ( .A(n24260), .B(n24261), .Z(n24251) );
  ANDN U24250 ( .B(n24262), .A(n24263), .Z(n24259) );
  NANDN U24251 ( .A(n24260), .B(n24265), .Z(n24255) );
  XOR U24252 ( .A(n24266), .B(n24253), .Z(n24260) );
  XNOR U24253 ( .A(n24267), .B(n24268), .Z(n24253) );
  XOR U24254 ( .A(n24269), .B(n24262), .Z(n24268) );
  XNOR U24255 ( .A(n24270), .B(n24271), .Z(n24267) );
  XNOR U24256 ( .A(n24272), .B(n24273), .Z(n24271) );
  ANDN U24257 ( .B(n24262), .A(n24274), .Z(n24272) );
  IV U24258 ( .A(n24275), .Z(n24262) );
  ANDN U24259 ( .B(n24266), .A(n24274), .Z(n24264) );
  IV U24260 ( .A(n24270), .Z(n24274) );
  IV U24261 ( .A(n24263), .Z(n24266) );
  XNOR U24262 ( .A(n24269), .B(n24276), .Z(n24263) );
  XOR U24263 ( .A(n24277), .B(n24273), .Z(n24276) );
  NAND U24264 ( .A(n24265), .B(n24261), .Z(n24273) );
  XNOR U24265 ( .A(n24254), .B(n24275), .Z(n24261) );
  XOR U24266 ( .A(n24278), .B(n24279), .Z(n24275) );
  XOR U24267 ( .A(n24280), .B(n24281), .Z(n24279) );
  XNOR U24268 ( .A(n24014), .B(n24282), .Z(n24281) );
  XNOR U24269 ( .A(n24283), .B(n24284), .Z(n24278) );
  XNOR U24270 ( .A(n24285), .B(n24286), .Z(n24284) );
  ANDN U24271 ( .B(n24287), .A(n23910), .Z(n24285) );
  XNOR U24272 ( .A(n24270), .B(n24257), .Z(n24265) );
  XOR U24273 ( .A(n24288), .B(n24289), .Z(n24270) );
  XNOR U24274 ( .A(n24290), .B(n24282), .Z(n24289) );
  XOR U24275 ( .A(n24291), .B(n24292), .Z(n24282) );
  XNOR U24276 ( .A(n24293), .B(n24294), .Z(n24292) );
  NAND U24277 ( .A(n24244), .B(n24023), .Z(n24294) );
  XNOR U24278 ( .A(n24295), .B(n24296), .Z(n24288) );
  ANDN U24279 ( .B(n24297), .A(n24240), .Z(n24295) );
  ANDN U24280 ( .B(n24254), .A(n24257), .Z(n24277) );
  XOR U24281 ( .A(n24257), .B(n24254), .Z(n24269) );
  XNOR U24282 ( .A(n24298), .B(n24299), .Z(n24254) );
  XNOR U24283 ( .A(n24291), .B(n24300), .Z(n24299) );
  XOR U24284 ( .A(n24290), .B(n24017), .Z(n24300) );
  XOR U24285 ( .A(n23910), .B(n24301), .Z(n24298) );
  XNOR U24286 ( .A(n24302), .B(n24286), .Z(n24301) );
  OR U24287 ( .A(n24019), .B(n24247), .Z(n24286) );
  XNOR U24288 ( .A(n23910), .B(n24248), .Z(n24247) );
  XOR U24289 ( .A(n24017), .B(n24014), .Z(n24019) );
  ANDN U24290 ( .B(n24014), .A(n24248), .Z(n24302) );
  XOR U24291 ( .A(n24303), .B(n24304), .Z(n24257) );
  XOR U24292 ( .A(n24291), .B(n24280), .Z(n24304) );
  XOR U24293 ( .A(n24034), .B(n23880), .Z(n24280) );
  XOR U24294 ( .A(n24305), .B(n24293), .Z(n24291) );
  NANDN U24295 ( .A(n24250), .B(n24027), .Z(n24293) );
  XOR U24296 ( .A(n24029), .B(n24023), .Z(n24027) );
  XNOR U24297 ( .A(n24297), .B(n24306), .Z(n24014) );
  XNOR U24298 ( .A(n24307), .B(n24308), .Z(n24306) );
  XOR U24299 ( .A(n24258), .B(n24244), .Z(n24250) );
  XNOR U24300 ( .A(n24248), .B(n24034), .Z(n24244) );
  IV U24301 ( .A(n24283), .Z(n24248) );
  XOR U24302 ( .A(n24309), .B(n24310), .Z(n24283) );
  XOR U24303 ( .A(n24311), .B(n24312), .Z(n24310) );
  XNOR U24304 ( .A(n23910), .B(n24313), .Z(n24309) );
  ANDN U24305 ( .B(n24029), .A(n24258), .Z(n24305) );
  XNOR U24306 ( .A(n23910), .B(n24240), .Z(n24258) );
  XOR U24307 ( .A(n24297), .B(n24287), .Z(n24029) );
  IV U24308 ( .A(n24017), .Z(n24287) );
  XOR U24309 ( .A(n24314), .B(n24315), .Z(n24017) );
  XOR U24310 ( .A(n24316), .B(n24312), .Z(n24315) );
  XNOR U24311 ( .A(n24317), .B(n24318), .Z(n24312) );
  XNOR U24312 ( .A(n24319), .B(n24320), .Z(n24318) );
  XNOR U24313 ( .A(n24321), .B(n24322), .Z(n24317) );
  XNOR U24314 ( .A(key[252]), .B(n24323), .Z(n24322) );
  IV U24315 ( .A(n24008), .Z(n24297) );
  XOR U24316 ( .A(n24290), .B(n24324), .Z(n24303) );
  XNOR U24317 ( .A(n24325), .B(n24296), .Z(n24324) );
  OR U24318 ( .A(n24006), .B(n24239), .Z(n24296) );
  XNOR U24319 ( .A(n24326), .B(n24034), .Z(n24239) );
  XNOR U24320 ( .A(n24008), .B(n23880), .Z(n24006) );
  ANDN U24321 ( .B(n24034), .A(n23880), .Z(n24325) );
  XOR U24322 ( .A(n24314), .B(n24327), .Z(n23880) );
  XOR U24323 ( .A(n24307), .B(n24328), .Z(n24327) );
  XOR U24324 ( .A(n24316), .B(n24314), .Z(n24034) );
  XNOR U24325 ( .A(n24240), .B(n24008), .Z(n24290) );
  XOR U24326 ( .A(n24314), .B(n24329), .Z(n24008) );
  XNOR U24327 ( .A(n24316), .B(n24311), .Z(n24329) );
  XOR U24328 ( .A(n24330), .B(n24331), .Z(n24311) );
  XOR U24329 ( .A(n24332), .B(n24333), .Z(n24331) );
  XNOR U24330 ( .A(key[255]), .B(n24334), .Z(n24330) );
  XNOR U24331 ( .A(n24335), .B(n24336), .Z(n24314) );
  XOR U24332 ( .A(n24337), .B(n24338), .Z(n24336) );
  XOR U24333 ( .A(n24339), .B(n24340), .Z(n24335) );
  XNOR U24334 ( .A(key[253]), .B(n24341), .Z(n24340) );
  IV U24335 ( .A(n24326), .Z(n24240) );
  XNOR U24336 ( .A(n24308), .B(n24342), .Z(n24326) );
  XOR U24337 ( .A(n24313), .B(n24328), .Z(n24342) );
  IV U24338 ( .A(n24316), .Z(n24328) );
  XOR U24339 ( .A(n24343), .B(n24344), .Z(n24316) );
  XOR U24340 ( .A(n24345), .B(n24346), .Z(n24344) );
  XOR U24341 ( .A(n24347), .B(n24348), .Z(n24343) );
  XOR U24342 ( .A(key[254]), .B(n23910), .Z(n24348) );
  XNOR U24343 ( .A(n24349), .B(n24350), .Z(n23910) );
  XOR U24344 ( .A(n24351), .B(n24352), .Z(n24350) );
  XNOR U24345 ( .A(n24353), .B(n24354), .Z(n24349) );
  XOR U24346 ( .A(key[248]), .B(n24355), .Z(n24354) );
  XOR U24347 ( .A(n24356), .B(n24357), .Z(n24313) );
  XOR U24348 ( .A(n24358), .B(n24359), .Z(n24357) );
  XOR U24349 ( .A(n24307), .B(n24360), .Z(n24359) );
  XOR U24350 ( .A(n24361), .B(n24362), .Z(n24307) );
  XOR U24351 ( .A(n24363), .B(n24364), .Z(n24362) );
  XNOR U24352 ( .A(n24365), .B(n24366), .Z(n24361) );
  XNOR U24353 ( .A(key[249]), .B(n24367), .Z(n24366) );
  XNOR U24354 ( .A(n24368), .B(n24369), .Z(n24356) );
  XNOR U24355 ( .A(key[251]), .B(n24370), .Z(n24369) );
  XOR U24356 ( .A(n24371), .B(n24372), .Z(n24308) );
  XOR U24357 ( .A(n24373), .B(n24374), .Z(n24372) );
  XOR U24358 ( .A(n24375), .B(n24376), .Z(n24371) );
  XNOR U24359 ( .A(key[250]), .B(n24377), .Z(n24376) );
  XOR U24360 ( .A(n23161), .B(n21376), .Z(n21358) );
  IV U24361 ( .A(n23129), .Z(n21376) );
  XNOR U24362 ( .A(n23865), .B(n23920), .Z(n23129) );
  XOR U24363 ( .A(n23977), .B(n24378), .Z(n23920) );
  XOR U24364 ( .A(n24379), .B(n23898), .Z(n24378) );
  OR U24365 ( .A(n24380), .B(n23990), .Z(n23898) );
  XNOR U24366 ( .A(n23901), .B(n23986), .Z(n23990) );
  ANDN U24367 ( .B(n23986), .A(n24381), .Z(n24379) );
  IV U24368 ( .A(n24382), .Z(n23977) );
  IV U24369 ( .A(n23918), .Z(n23865) );
  XNOR U24370 ( .A(n24384), .B(n23979), .Z(n24383) );
  XNOR U24371 ( .A(n23976), .B(n23869), .Z(n23973) );
  ANDN U24372 ( .B(n24386), .A(n23976), .Z(n24384) );
  XOR U24373 ( .A(n24382), .B(n24387), .Z(n23896) );
  XNOR U24374 ( .A(n24388), .B(n24389), .Z(n24387) );
  NAND U24375 ( .A(n23996), .B(n24390), .Z(n24389) );
  XNOR U24376 ( .A(n24391), .B(n24388), .Z(n24382) );
  OR U24377 ( .A(n24392), .B(n23998), .Z(n24388) );
  XOR U24378 ( .A(n24001), .B(n23996), .Z(n23998) );
  XOR U24379 ( .A(n23986), .B(n23869), .Z(n23996) );
  XOR U24380 ( .A(n24393), .B(n24394), .Z(n23869) );
  NANDN U24381 ( .A(n24395), .B(n24396), .Z(n24394) );
  XOR U24382 ( .A(n24397), .B(n24398), .Z(n23986) );
  NANDN U24383 ( .A(n24395), .B(n24399), .Z(n24398) );
  NOR U24384 ( .A(n24001), .B(n24400), .Z(n24391) );
  XOR U24385 ( .A(n23976), .B(n23901), .Z(n24001) );
  XNOR U24386 ( .A(n24401), .B(n24397), .Z(n23901) );
  NANDN U24387 ( .A(n24402), .B(n24403), .Z(n24397) );
  XOR U24388 ( .A(n24399), .B(n24404), .Z(n24403) );
  ANDN U24389 ( .B(n24404), .A(n24405), .Z(n24401) );
  XOR U24390 ( .A(n24406), .B(n24393), .Z(n23976) );
  NANDN U24391 ( .A(n24402), .B(n24407), .Z(n24393) );
  XOR U24392 ( .A(n24408), .B(n24396), .Z(n24407) );
  XNOR U24393 ( .A(n24409), .B(n24410), .Z(n24395) );
  XOR U24394 ( .A(n24411), .B(n24412), .Z(n24410) );
  XNOR U24395 ( .A(n24413), .B(n24414), .Z(n24409) );
  XNOR U24396 ( .A(n24415), .B(n24416), .Z(n24414) );
  ANDN U24397 ( .B(n24408), .A(n24412), .Z(n24415) );
  ANDN U24398 ( .B(n24408), .A(n24405), .Z(n24406) );
  XNOR U24399 ( .A(n24411), .B(n24417), .Z(n24405) );
  XOR U24400 ( .A(n24418), .B(n24416), .Z(n24417) );
  NAND U24401 ( .A(n24419), .B(n24420), .Z(n24416) );
  XNOR U24402 ( .A(n24413), .B(n24396), .Z(n24420) );
  IV U24403 ( .A(n24408), .Z(n24413) );
  XNOR U24404 ( .A(n24399), .B(n24412), .Z(n24419) );
  IV U24405 ( .A(n24404), .Z(n24412) );
  XOR U24406 ( .A(n24421), .B(n24422), .Z(n24404) );
  XNOR U24407 ( .A(n24423), .B(n24424), .Z(n24422) );
  XNOR U24408 ( .A(n24425), .B(n24426), .Z(n24421) );
  ANDN U24409 ( .B(n24386), .A(n23975), .Z(n24425) );
  AND U24410 ( .A(n24396), .B(n24399), .Z(n24418) );
  XNOR U24411 ( .A(n24396), .B(n24399), .Z(n24411) );
  XNOR U24412 ( .A(n24427), .B(n24428), .Z(n24399) );
  XNOR U24413 ( .A(n24429), .B(n24424), .Z(n24428) );
  XOR U24414 ( .A(n24430), .B(n24431), .Z(n24427) );
  XNOR U24415 ( .A(n24432), .B(n24426), .Z(n24431) );
  OR U24416 ( .A(n23974), .B(n24385), .Z(n24426) );
  XNOR U24417 ( .A(n24386), .B(n24433), .Z(n24385) );
  XNOR U24418 ( .A(n23975), .B(n23870), .Z(n23974) );
  ANDN U24419 ( .B(n24434), .A(n23981), .Z(n24432) );
  XNOR U24420 ( .A(n24435), .B(n24436), .Z(n24396) );
  XNOR U24421 ( .A(n24424), .B(n24437), .Z(n24436) );
  XOR U24422 ( .A(n23989), .B(n24430), .Z(n24437) );
  XNOR U24423 ( .A(n24386), .B(n23975), .Z(n24424) );
  XOR U24424 ( .A(n23900), .B(n24438), .Z(n24435) );
  XNOR U24425 ( .A(n24439), .B(n24440), .Z(n24438) );
  ANDN U24426 ( .B(n24441), .A(n24381), .Z(n24439) );
  XNOR U24427 ( .A(n24442), .B(n24443), .Z(n24408) );
  XNOR U24428 ( .A(n24429), .B(n24444), .Z(n24443) );
  XNOR U24429 ( .A(n23985), .B(n24423), .Z(n24444) );
  XOR U24430 ( .A(n24430), .B(n24445), .Z(n24423) );
  XNOR U24431 ( .A(n24446), .B(n24447), .Z(n24445) );
  NAND U24432 ( .A(n24390), .B(n23995), .Z(n24447) );
  XNOR U24433 ( .A(n24448), .B(n24446), .Z(n24430) );
  NANDN U24434 ( .A(n24392), .B(n23999), .Z(n24446) );
  XOR U24435 ( .A(n24000), .B(n23995), .Z(n23999) );
  XNOR U24436 ( .A(n24441), .B(n23870), .Z(n23995) );
  XOR U24437 ( .A(n24400), .B(n24390), .Z(n24392) );
  XNOR U24438 ( .A(n24381), .B(n24433), .Z(n24390) );
  ANDN U24439 ( .B(n24000), .A(n24400), .Z(n24448) );
  XOR U24440 ( .A(n23900), .B(n24386), .Z(n24400) );
  XNOR U24441 ( .A(n24449), .B(n24450), .Z(n24386) );
  XNOR U24442 ( .A(n24451), .B(n24452), .Z(n24450) );
  XOR U24443 ( .A(n24433), .B(n24434), .Z(n24429) );
  IV U24444 ( .A(n23870), .Z(n24434) );
  XOR U24445 ( .A(n24454), .B(n24455), .Z(n23870) );
  XNOR U24446 ( .A(n24456), .B(n24452), .Z(n24455) );
  IV U24447 ( .A(n23981), .Z(n24433) );
  XOR U24448 ( .A(n24452), .B(n24457), .Z(n23981) );
  XNOR U24449 ( .A(n24458), .B(n24459), .Z(n24442) );
  XNOR U24450 ( .A(n24460), .B(n24440), .Z(n24459) );
  OR U24451 ( .A(n23991), .B(n24380), .Z(n24440) );
  XNOR U24452 ( .A(n23900), .B(n24381), .Z(n24380) );
  IV U24453 ( .A(n24458), .Z(n24381) );
  XOR U24454 ( .A(n23989), .B(n24441), .Z(n23991) );
  IV U24455 ( .A(n23985), .Z(n24441) );
  XOR U24456 ( .A(n24453), .B(n24461), .Z(n23985) );
  XNOR U24457 ( .A(n24456), .B(n24449), .Z(n24461) );
  XOR U24458 ( .A(n24462), .B(n24463), .Z(n24449) );
  XNOR U24459 ( .A(n24464), .B(n24465), .Z(n24463) );
  XOR U24460 ( .A(key[130]), .B(n24466), .Z(n24462) );
  IV U24461 ( .A(n23975), .Z(n24453) );
  XOR U24462 ( .A(n24454), .B(n24467), .Z(n23975) );
  XOR U24463 ( .A(n24452), .B(n24468), .Z(n24467) );
  NOR U24464 ( .A(n23989), .B(n23900), .Z(n24460) );
  XOR U24465 ( .A(n24454), .B(n24469), .Z(n23989) );
  XOR U24466 ( .A(n24452), .B(n24470), .Z(n24469) );
  XOR U24467 ( .A(n24471), .B(n24472), .Z(n24452) );
  XNOR U24468 ( .A(n24473), .B(n24474), .Z(n24472) );
  XNOR U24469 ( .A(n24475), .B(n24476), .Z(n24471) );
  XOR U24470 ( .A(key[134]), .B(n23900), .Z(n24476) );
  IV U24471 ( .A(n24457), .Z(n24454) );
  XOR U24472 ( .A(n24477), .B(n24478), .Z(n24457) );
  XNOR U24473 ( .A(n24479), .B(n24480), .Z(n24478) );
  XNOR U24474 ( .A(key[133]), .B(n24481), .Z(n24477) );
  XOR U24475 ( .A(n24482), .B(n24483), .Z(n24458) );
  XNOR U24476 ( .A(n24470), .B(n24468), .Z(n24483) );
  XNOR U24477 ( .A(n24484), .B(n24485), .Z(n24468) );
  XOR U24478 ( .A(n24486), .B(n24487), .Z(n24485) );
  XNOR U24479 ( .A(key[135]), .B(n24488), .Z(n24484) );
  XNOR U24480 ( .A(n24489), .B(n24490), .Z(n24470) );
  XNOR U24481 ( .A(n24491), .B(n24492), .Z(n24490) );
  XNOR U24482 ( .A(n24493), .B(n24494), .Z(n24489) );
  XNOR U24483 ( .A(key[132]), .B(n24495), .Z(n24494) );
  XNOR U24484 ( .A(n23900), .B(n24451), .Z(n24482) );
  XOR U24485 ( .A(n24496), .B(n24497), .Z(n24451) );
  XOR U24486 ( .A(n24498), .B(n24499), .Z(n24497) );
  XNOR U24487 ( .A(n24456), .B(n24500), .Z(n24499) );
  XOR U24488 ( .A(n24501), .B(n24502), .Z(n24456) );
  XOR U24489 ( .A(key[129]), .B(n24505), .Z(n24501) );
  XOR U24490 ( .A(n24506), .B(n24507), .Z(n24496) );
  XNOR U24491 ( .A(key[131]), .B(n24508), .Z(n24507) );
  XNOR U24492 ( .A(n24509), .B(n24510), .Z(n23900) );
  XOR U24493 ( .A(n24511), .B(n24512), .Z(n24510) );
  XNOR U24494 ( .A(key[128]), .B(n24513), .Z(n24509) );
  XNOR U24495 ( .A(n23932), .B(n23967), .Z(n23161) );
  XNOR U24496 ( .A(n24081), .B(n24514), .Z(n23967) );
  XOR U24497 ( .A(n24515), .B(n23928), .Z(n24514) );
  OR U24498 ( .A(n24516), .B(n24069), .Z(n23928) );
  XNOR U24499 ( .A(n23931), .B(n24065), .Z(n24069) );
  ANDN U24500 ( .B(n24065), .A(n24517), .Z(n24515) );
  IV U24501 ( .A(n24518), .Z(n24081) );
  XNOR U24502 ( .A(n23926), .B(n24519), .Z(n23932) );
  XNOR U24503 ( .A(n24520), .B(n24083), .Z(n24519) );
  XNOR U24504 ( .A(n24044), .B(n23936), .Z(n24041) );
  ANDN U24505 ( .B(n24522), .A(n24044), .Z(n24520) );
  XOR U24506 ( .A(n24518), .B(n24523), .Z(n23926) );
  XNOR U24507 ( .A(n24524), .B(n24525), .Z(n24523) );
  NAND U24508 ( .A(n24075), .B(n24526), .Z(n24525) );
  XNOR U24509 ( .A(n24527), .B(n24524), .Z(n24518) );
  OR U24510 ( .A(n24528), .B(n24077), .Z(n24524) );
  XOR U24511 ( .A(n24080), .B(n24075), .Z(n24077) );
  XOR U24512 ( .A(n24065), .B(n23936), .Z(n24075) );
  XOR U24513 ( .A(n24529), .B(n24530), .Z(n23936) );
  NANDN U24514 ( .A(n24531), .B(n24532), .Z(n24530) );
  XOR U24515 ( .A(n24533), .B(n24534), .Z(n24065) );
  NANDN U24516 ( .A(n24531), .B(n24535), .Z(n24534) );
  NOR U24517 ( .A(n24080), .B(n24536), .Z(n24527) );
  XOR U24518 ( .A(n24044), .B(n23931), .Z(n24080) );
  XNOR U24519 ( .A(n24537), .B(n24533), .Z(n23931) );
  NANDN U24520 ( .A(n24538), .B(n24539), .Z(n24533) );
  XOR U24521 ( .A(n24535), .B(n24540), .Z(n24539) );
  ANDN U24522 ( .B(n24540), .A(n24541), .Z(n24537) );
  XOR U24523 ( .A(n24542), .B(n24529), .Z(n24044) );
  NANDN U24524 ( .A(n24538), .B(n24543), .Z(n24529) );
  XOR U24525 ( .A(n24544), .B(n24532), .Z(n24543) );
  XNOR U24526 ( .A(n24545), .B(n24546), .Z(n24531) );
  XOR U24527 ( .A(n24547), .B(n24548), .Z(n24546) );
  XNOR U24528 ( .A(n24549), .B(n24550), .Z(n24545) );
  XNOR U24529 ( .A(n24551), .B(n24552), .Z(n24550) );
  ANDN U24530 ( .B(n24544), .A(n24548), .Z(n24551) );
  ANDN U24531 ( .B(n24544), .A(n24541), .Z(n24542) );
  XNOR U24532 ( .A(n24547), .B(n24553), .Z(n24541) );
  XOR U24533 ( .A(n24554), .B(n24552), .Z(n24553) );
  NAND U24534 ( .A(n24555), .B(n24556), .Z(n24552) );
  XNOR U24535 ( .A(n24549), .B(n24532), .Z(n24556) );
  IV U24536 ( .A(n24544), .Z(n24549) );
  XNOR U24537 ( .A(n24535), .B(n24548), .Z(n24555) );
  IV U24538 ( .A(n24540), .Z(n24548) );
  XOR U24539 ( .A(n24557), .B(n24558), .Z(n24540) );
  XNOR U24540 ( .A(n24559), .B(n24560), .Z(n24558) );
  XNOR U24541 ( .A(n24561), .B(n24562), .Z(n24557) );
  ANDN U24542 ( .B(n24522), .A(n24043), .Z(n24561) );
  AND U24543 ( .A(n24532), .B(n24535), .Z(n24554) );
  XNOR U24544 ( .A(n24532), .B(n24535), .Z(n24547) );
  XNOR U24545 ( .A(n24563), .B(n24564), .Z(n24535) );
  XNOR U24546 ( .A(n24565), .B(n24560), .Z(n24564) );
  XOR U24547 ( .A(n24566), .B(n24567), .Z(n24563) );
  XNOR U24548 ( .A(n24568), .B(n24562), .Z(n24567) );
  OR U24549 ( .A(n24042), .B(n24521), .Z(n24562) );
  XNOR U24550 ( .A(n24522), .B(n24569), .Z(n24521) );
  XNOR U24551 ( .A(n24043), .B(n23937), .Z(n24042) );
  ANDN U24552 ( .B(n24570), .A(n24085), .Z(n24568) );
  XNOR U24553 ( .A(n24571), .B(n24572), .Z(n24532) );
  XNOR U24554 ( .A(n24560), .B(n24573), .Z(n24572) );
  XOR U24555 ( .A(n24068), .B(n24566), .Z(n24573) );
  XNOR U24556 ( .A(n24522), .B(n24043), .Z(n24560) );
  XOR U24557 ( .A(n23930), .B(n24574), .Z(n24571) );
  XNOR U24558 ( .A(n24575), .B(n24576), .Z(n24574) );
  ANDN U24559 ( .B(n24577), .A(n24517), .Z(n24575) );
  XNOR U24560 ( .A(n24578), .B(n24579), .Z(n24544) );
  XNOR U24561 ( .A(n24565), .B(n24580), .Z(n24579) );
  XNOR U24562 ( .A(n24064), .B(n24559), .Z(n24580) );
  XOR U24563 ( .A(n24566), .B(n24581), .Z(n24559) );
  XNOR U24564 ( .A(n24582), .B(n24583), .Z(n24581) );
  NAND U24565 ( .A(n24526), .B(n24074), .Z(n24583) );
  XNOR U24566 ( .A(n24584), .B(n24582), .Z(n24566) );
  NANDN U24567 ( .A(n24528), .B(n24078), .Z(n24582) );
  XOR U24568 ( .A(n24079), .B(n24074), .Z(n24078) );
  XNOR U24569 ( .A(n24577), .B(n23937), .Z(n24074) );
  XOR U24570 ( .A(n24536), .B(n24526), .Z(n24528) );
  XNOR U24571 ( .A(n24517), .B(n24569), .Z(n24526) );
  ANDN U24572 ( .B(n24079), .A(n24536), .Z(n24584) );
  XOR U24573 ( .A(n23930), .B(n24522), .Z(n24536) );
  XNOR U24574 ( .A(n24585), .B(n24586), .Z(n24522) );
  XNOR U24575 ( .A(n24587), .B(n24588), .Z(n24586) );
  XOR U24576 ( .A(n24569), .B(n24570), .Z(n24565) );
  IV U24577 ( .A(n23937), .Z(n24570) );
  XOR U24578 ( .A(n24590), .B(n24591), .Z(n23937) );
  XNOR U24579 ( .A(n24592), .B(n24588), .Z(n24591) );
  IV U24580 ( .A(n24085), .Z(n24569) );
  XOR U24581 ( .A(n24588), .B(n24593), .Z(n24085) );
  XNOR U24582 ( .A(n24594), .B(n24595), .Z(n24578) );
  XNOR U24583 ( .A(n24596), .B(n24576), .Z(n24595) );
  OR U24584 ( .A(n24070), .B(n24516), .Z(n24576) );
  XNOR U24585 ( .A(n23930), .B(n24517), .Z(n24516) );
  IV U24586 ( .A(n24594), .Z(n24517) );
  XOR U24587 ( .A(n24068), .B(n24577), .Z(n24070) );
  IV U24588 ( .A(n24064), .Z(n24577) );
  XOR U24589 ( .A(n24589), .B(n24597), .Z(n24064) );
  XNOR U24590 ( .A(n24592), .B(n24585), .Z(n24597) );
  XOR U24591 ( .A(n24598), .B(n24599), .Z(n24585) );
  XOR U24592 ( .A(n24602), .B(n24603), .Z(n24598) );
  XNOR U24593 ( .A(key[170]), .B(n24604), .Z(n24603) );
  IV U24594 ( .A(n24043), .Z(n24589) );
  XOR U24595 ( .A(n24590), .B(n24605), .Z(n24043) );
  XOR U24596 ( .A(n24588), .B(n24606), .Z(n24605) );
  NOR U24597 ( .A(n24068), .B(n23930), .Z(n24596) );
  XOR U24598 ( .A(n24590), .B(n24607), .Z(n24068) );
  XOR U24599 ( .A(n24588), .B(n24608), .Z(n24607) );
  XOR U24600 ( .A(n24609), .B(n24610), .Z(n24588) );
  XNOR U24601 ( .A(n24613), .B(n24614), .Z(n24609) );
  XOR U24602 ( .A(key[174]), .B(n23930), .Z(n24614) );
  IV U24603 ( .A(n24593), .Z(n24590) );
  XOR U24604 ( .A(n24615), .B(n24616), .Z(n24593) );
  XOR U24605 ( .A(n24617), .B(n24618), .Z(n24616) );
  XNOR U24606 ( .A(n24619), .B(n24620), .Z(n24615) );
  XOR U24607 ( .A(key[173]), .B(n24621), .Z(n24620) );
  XOR U24608 ( .A(n24622), .B(n24623), .Z(n24594) );
  XNOR U24609 ( .A(n24608), .B(n24606), .Z(n24623) );
  XNOR U24610 ( .A(n24624), .B(n24625), .Z(n24606) );
  XOR U24611 ( .A(n24626), .B(n24627), .Z(n24625) );
  XNOR U24612 ( .A(key[175]), .B(n24628), .Z(n24624) );
  XNOR U24613 ( .A(n24629), .B(n24630), .Z(n24608) );
  XNOR U24614 ( .A(n24631), .B(n24632), .Z(n24630) );
  XNOR U24615 ( .A(n24633), .B(n24634), .Z(n24629) );
  XNOR U24616 ( .A(key[172]), .B(n24635), .Z(n24634) );
  XNOR U24617 ( .A(n23930), .B(n24587), .Z(n24622) );
  XOR U24618 ( .A(n24636), .B(n24637), .Z(n24587) );
  XNOR U24619 ( .A(n24638), .B(n24639), .Z(n24637) );
  XOR U24620 ( .A(n24592), .B(n24640), .Z(n24639) );
  XOR U24621 ( .A(n24641), .B(n24642), .Z(n24592) );
  XNOR U24622 ( .A(n24643), .B(n24644), .Z(n24642) );
  XNOR U24623 ( .A(n24645), .B(n24646), .Z(n24641) );
  XNOR U24624 ( .A(key[169]), .B(n24647), .Z(n24646) );
  XNOR U24625 ( .A(n24648), .B(n24649), .Z(n24636) );
  XNOR U24626 ( .A(key[171]), .B(n24650), .Z(n24649) );
  XNOR U24627 ( .A(n24651), .B(n24652), .Z(n23930) );
  XOR U24628 ( .A(n24653), .B(n24654), .Z(n24652) );
  XNOR U24629 ( .A(n24655), .B(n24656), .Z(n24651) );
  XOR U24630 ( .A(key[168]), .B(n24657), .Z(n24656) );
  XNOR U24631 ( .A(n20014), .B(n18484), .Z(n19398) );
  XNOR U24632 ( .A(n24658), .B(n24659), .Z(n18484) );
  XOR U24633 ( .A(n23644), .B(n23622), .Z(n24659) );
  XNOR U24634 ( .A(n24660), .B(n24661), .Z(n23622) );
  XNOR U24635 ( .A(n23711), .B(n24662), .Z(n24661) );
  NANDN U24636 ( .A(n24663), .B(n23628), .Z(n24662) );
  OR U24637 ( .A(n24664), .B(n23642), .Z(n23711) );
  XNOR U24638 ( .A(n23628), .B(n23641), .Z(n23642) );
  XNOR U24639 ( .A(n24665), .B(n23651), .Z(n23644) );
  NANDN U24640 ( .A(n24666), .B(n24667), .Z(n23651) );
  ANDN U24641 ( .B(n24668), .A(n24669), .Z(n24665) );
  XNOR U24642 ( .A(n23590), .B(n24670), .Z(n24658) );
  XOR U24643 ( .A(n23647), .B(n24671), .Z(n24670) );
  ANDN U24644 ( .B(n23634), .A(n24672), .Z(n24671) );
  ANDN U24645 ( .B(n24673), .A(n24674), .Z(n23647) );
  XNOR U24646 ( .A(n24660), .B(n24675), .Z(n23590) );
  XNOR U24647 ( .A(n24676), .B(n23631), .Z(n24675) );
  XNOR U24648 ( .A(n23649), .B(n23634), .Z(n24673) );
  ANDN U24649 ( .B(n24678), .A(n23649), .Z(n24676) );
  XNOR U24650 ( .A(n23629), .B(n24679), .Z(n24660) );
  XNOR U24651 ( .A(n24680), .B(n24681), .Z(n24679) );
  NAND U24652 ( .A(n23654), .B(n24682), .Z(n24681) );
  XOR U24653 ( .A(n24683), .B(n24680), .Z(n23629) );
  OR U24654 ( .A(n24666), .B(n24684), .Z(n24680) );
  XNOR U24655 ( .A(n24685), .B(n23654), .Z(n24666) );
  XOR U24656 ( .A(n23641), .B(n23634), .Z(n23654) );
  XOR U24657 ( .A(n24686), .B(n24687), .Z(n23634) );
  NANDN U24658 ( .A(n24688), .B(n24689), .Z(n24687) );
  XOR U24659 ( .A(n24690), .B(n24691), .Z(n23641) );
  NANDN U24660 ( .A(n24688), .B(n24692), .Z(n24691) );
  ANDN U24661 ( .B(n24685), .A(n24693), .Z(n24683) );
  IV U24662 ( .A(n24669), .Z(n24685) );
  XOR U24663 ( .A(n23649), .B(n23628), .Z(n24669) );
  XNOR U24664 ( .A(n24694), .B(n24690), .Z(n23628) );
  NANDN U24665 ( .A(n24695), .B(n24696), .Z(n24690) );
  XOR U24666 ( .A(n24692), .B(n24697), .Z(n24696) );
  ANDN U24667 ( .B(n24697), .A(n24698), .Z(n24694) );
  XOR U24668 ( .A(n24699), .B(n24686), .Z(n23649) );
  NANDN U24669 ( .A(n24695), .B(n24700), .Z(n24686) );
  XOR U24670 ( .A(n24701), .B(n24689), .Z(n24700) );
  XNOR U24671 ( .A(n24702), .B(n24703), .Z(n24688) );
  XOR U24672 ( .A(n24704), .B(n24705), .Z(n24703) );
  XNOR U24673 ( .A(n24706), .B(n24707), .Z(n24702) );
  XNOR U24674 ( .A(n24708), .B(n24709), .Z(n24707) );
  ANDN U24675 ( .B(n24701), .A(n24705), .Z(n24708) );
  ANDN U24676 ( .B(n24701), .A(n24698), .Z(n24699) );
  XNOR U24677 ( .A(n24704), .B(n24710), .Z(n24698) );
  XOR U24678 ( .A(n24711), .B(n24709), .Z(n24710) );
  NAND U24679 ( .A(n24712), .B(n24713), .Z(n24709) );
  XNOR U24680 ( .A(n24706), .B(n24689), .Z(n24713) );
  IV U24681 ( .A(n24701), .Z(n24706) );
  XNOR U24682 ( .A(n24692), .B(n24705), .Z(n24712) );
  IV U24683 ( .A(n24697), .Z(n24705) );
  XOR U24684 ( .A(n24714), .B(n24715), .Z(n24697) );
  XNOR U24685 ( .A(n24716), .B(n24717), .Z(n24715) );
  XNOR U24686 ( .A(n24718), .B(n24719), .Z(n24714) );
  ANDN U24687 ( .B(n24678), .A(n23648), .Z(n24718) );
  AND U24688 ( .A(n24689), .B(n24692), .Z(n24711) );
  XNOR U24689 ( .A(n24689), .B(n24692), .Z(n24704) );
  XNOR U24690 ( .A(n24720), .B(n24721), .Z(n24692) );
  XNOR U24691 ( .A(n24722), .B(n24717), .Z(n24721) );
  XOR U24692 ( .A(n24723), .B(n24724), .Z(n24720) );
  XNOR U24693 ( .A(n24725), .B(n24719), .Z(n24724) );
  OR U24694 ( .A(n24674), .B(n24677), .Z(n24719) );
  XNOR U24695 ( .A(n24678), .B(n24726), .Z(n24677) );
  XNOR U24696 ( .A(n23648), .B(n24672), .Z(n24674) );
  ANDN U24697 ( .B(n24727), .A(n23633), .Z(n24725) );
  XNOR U24698 ( .A(n24728), .B(n24729), .Z(n24689) );
  XNOR U24699 ( .A(n24717), .B(n24730), .Z(n24729) );
  XOR U24700 ( .A(n23627), .B(n24723), .Z(n24730) );
  XNOR U24701 ( .A(n24678), .B(n23648), .Z(n24717) );
  XOR U24702 ( .A(n24663), .B(n24731), .Z(n24728) );
  XNOR U24703 ( .A(n24732), .B(n24733), .Z(n24731) );
  ANDN U24704 ( .B(n24734), .A(n23712), .Z(n24732) );
  XNOR U24705 ( .A(n24735), .B(n24736), .Z(n24701) );
  XNOR U24706 ( .A(n24722), .B(n24737), .Z(n24736) );
  XNOR U24707 ( .A(n23640), .B(n24716), .Z(n24737) );
  XOR U24708 ( .A(n24723), .B(n24738), .Z(n24716) );
  XNOR U24709 ( .A(n24739), .B(n24740), .Z(n24738) );
  NAND U24710 ( .A(n24682), .B(n23653), .Z(n24740) );
  XNOR U24711 ( .A(n24741), .B(n24739), .Z(n24723) );
  NANDN U24712 ( .A(n24684), .B(n24667), .Z(n24739) );
  XOR U24713 ( .A(n24668), .B(n23653), .Z(n24667) );
  XNOR U24714 ( .A(n24734), .B(n24672), .Z(n23653) );
  XOR U24715 ( .A(n24693), .B(n24682), .Z(n24684) );
  XNOR U24716 ( .A(n23712), .B(n24726), .Z(n24682) );
  ANDN U24717 ( .B(n24668), .A(n24693), .Z(n24741) );
  XOR U24718 ( .A(n24663), .B(n24678), .Z(n24693) );
  XNOR U24719 ( .A(n24742), .B(n24743), .Z(n24678) );
  XNOR U24720 ( .A(n24744), .B(n24745), .Z(n24743) );
  XOR U24721 ( .A(n24726), .B(n24727), .Z(n24722) );
  IV U24722 ( .A(n24672), .Z(n24727) );
  XOR U24723 ( .A(n24747), .B(n24748), .Z(n24672) );
  XNOR U24724 ( .A(n24749), .B(n24745), .Z(n24748) );
  IV U24725 ( .A(n23633), .Z(n24726) );
  XOR U24726 ( .A(n24745), .B(n24750), .Z(n23633) );
  XNOR U24727 ( .A(n24751), .B(n24752), .Z(n24735) );
  XNOR U24728 ( .A(n24753), .B(n24733), .Z(n24752) );
  OR U24729 ( .A(n23643), .B(n24664), .Z(n24733) );
  XNOR U24730 ( .A(n24663), .B(n23712), .Z(n24664) );
  IV U24731 ( .A(n24751), .Z(n23712) );
  XOR U24732 ( .A(n23627), .B(n24734), .Z(n23643) );
  IV U24733 ( .A(n23640), .Z(n24734) );
  XOR U24734 ( .A(n24746), .B(n24754), .Z(n23640) );
  XNOR U24735 ( .A(n24749), .B(n24742), .Z(n24754) );
  XOR U24736 ( .A(n24755), .B(n24756), .Z(n24742) );
  XNOR U24737 ( .A(n22565), .B(n24757), .Z(n24756) );
  XNOR U24738 ( .A(n24758), .B(n24759), .Z(n22565) );
  XOR U24739 ( .A(n24760), .B(n24761), .Z(n24759) );
  XOR U24740 ( .A(n24762), .B(n24763), .Z(n24758) );
  XNOR U24741 ( .A(key[282]), .B(n23304), .Z(n24764) );
  IV U24742 ( .A(n23648), .Z(n24746) );
  XOR U24743 ( .A(n24747), .B(n24765), .Z(n23648) );
  XOR U24744 ( .A(n24745), .B(n24766), .Z(n24765) );
  NOR U24745 ( .A(n23627), .B(n24663), .Z(n24753) );
  XOR U24746 ( .A(n24747), .B(n24767), .Z(n23627) );
  XOR U24747 ( .A(n24745), .B(n24768), .Z(n24767) );
  XOR U24748 ( .A(n24769), .B(n24770), .Z(n24745) );
  XNOR U24749 ( .A(n22542), .B(n21542), .Z(n24770) );
  XOR U24750 ( .A(n21533), .B(n23284), .Z(n21542) );
  XNOR U24751 ( .A(n21549), .B(n22552), .Z(n22542) );
  XNOR U24752 ( .A(n21539), .B(n23285), .Z(n22552) );
  XOR U24753 ( .A(n24771), .B(n24772), .Z(n23285) );
  XNOR U24754 ( .A(n24773), .B(n24774), .Z(n24772) );
  XNOR U24755 ( .A(n24762), .B(n24775), .Z(n24771) );
  XNOR U24756 ( .A(n24776), .B(n21544), .Z(n21549) );
  XNOR U24757 ( .A(n24777), .B(n24778), .Z(n21544) );
  XNOR U24758 ( .A(n23291), .B(n24779), .Z(n24769) );
  XOR U24759 ( .A(key[286]), .B(n24663), .Z(n24779) );
  XOR U24760 ( .A(n24780), .B(n24781), .Z(n23291) );
  IV U24761 ( .A(n24750), .Z(n24747) );
  XOR U24762 ( .A(n24782), .B(n24783), .Z(n24750) );
  XOR U24763 ( .A(n23271), .B(n22545), .Z(n24783) );
  XNOR U24764 ( .A(n23289), .B(n21547), .Z(n22545) );
  XNOR U24765 ( .A(n24784), .B(n24785), .Z(n21547) );
  XNOR U24766 ( .A(n24786), .B(n24787), .Z(n24785) );
  XNOR U24767 ( .A(n24788), .B(n24789), .Z(n24784) );
  XOR U24768 ( .A(n24790), .B(n24791), .Z(n24789) );
  ANDN U24769 ( .B(n24792), .A(n24793), .Z(n24791) );
  XNOR U24770 ( .A(n24794), .B(n24795), .Z(n23271) );
  XNOR U24771 ( .A(n24796), .B(n24797), .Z(n24795) );
  XNOR U24772 ( .A(n24798), .B(n24799), .Z(n24794) );
  XNOR U24773 ( .A(n24800), .B(n24801), .Z(n24799) );
  ANDN U24774 ( .B(n24802), .A(n24803), .Z(n24801) );
  XOR U24775 ( .A(n23316), .B(n24804), .Z(n24782) );
  XOR U24776 ( .A(key[285]), .B(n24776), .Z(n24804) );
  IV U24777 ( .A(n23314), .Z(n24776) );
  XOR U24778 ( .A(n24805), .B(n24806), .Z(n23314) );
  XOR U24779 ( .A(n24773), .B(n24761), .Z(n23316) );
  XNOR U24780 ( .A(n24807), .B(n24808), .Z(n24761) );
  XNOR U24781 ( .A(n24809), .B(n24810), .Z(n24808) );
  NOR U24782 ( .A(n24811), .B(n24812), .Z(n24809) );
  XOR U24783 ( .A(n24813), .B(n24814), .Z(n24751) );
  XNOR U24784 ( .A(n24768), .B(n24766), .Z(n24814) );
  XNOR U24785 ( .A(n24815), .B(n24816), .Z(n24766) );
  XOR U24786 ( .A(n23286), .B(n22553), .Z(n24816) );
  XNOR U24787 ( .A(n23284), .B(n23315), .Z(n22553) );
  XNOR U24788 ( .A(n24817), .B(n24818), .Z(n23315) );
  XNOR U24789 ( .A(n24819), .B(n24787), .Z(n24818) );
  XNOR U24790 ( .A(n24820), .B(n24821), .Z(n24787) );
  XNOR U24791 ( .A(n24822), .B(n24823), .Z(n24821) );
  NANDN U24792 ( .A(n24824), .B(n24825), .Z(n24823) );
  XOR U24793 ( .A(n24826), .B(n24777), .Z(n24817) );
  XNOR U24794 ( .A(n24827), .B(n24828), .Z(n23284) );
  XNOR U24795 ( .A(n24829), .B(n24830), .Z(n24828) );
  XOR U24796 ( .A(n24831), .B(n24805), .Z(n24827) );
  XNOR U24797 ( .A(n24832), .B(n24833), .Z(n23286) );
  XOR U24798 ( .A(n24781), .B(n24797), .Z(n24833) );
  XNOR U24799 ( .A(n24834), .B(n24835), .Z(n24797) );
  XNOR U24800 ( .A(n24836), .B(n24837), .Z(n24835) );
  OR U24801 ( .A(n24838), .B(n24839), .Z(n24837) );
  XNOR U24802 ( .A(n24840), .B(n24841), .Z(n24832) );
  XNOR U24803 ( .A(key[287]), .B(n22575), .Z(n24815) );
  XOR U24804 ( .A(n24842), .B(n21539), .Z(n22575) );
  XNOR U24805 ( .A(n24843), .B(n24844), .Z(n24768) );
  XNOR U24806 ( .A(n22557), .B(n21525), .Z(n24844) );
  XOR U24807 ( .A(n21533), .B(n23289), .Z(n21525) );
  XNOR U24808 ( .A(n24845), .B(n24846), .Z(n23289) );
  XNOR U24809 ( .A(n24847), .B(n24830), .Z(n24846) );
  XNOR U24810 ( .A(n24848), .B(n24849), .Z(n24830) );
  XNOR U24811 ( .A(n24850), .B(n24851), .Z(n24849) );
  NANDN U24812 ( .A(n24852), .B(n24853), .Z(n24851) );
  XNOR U24813 ( .A(n24854), .B(n24855), .Z(n24845) );
  XOR U24814 ( .A(n24856), .B(n24857), .Z(n24855) );
  ANDN U24815 ( .B(n24858), .A(n24859), .Z(n24857) );
  XNOR U24816 ( .A(n23275), .B(n21527), .Z(n22557) );
  XOR U24817 ( .A(n24788), .B(n21519), .Z(n21527) );
  XOR U24818 ( .A(n23274), .B(n24861), .Z(n24843) );
  XNOR U24819 ( .A(key[284]), .B(n22559), .Z(n24861) );
  XNOR U24820 ( .A(n21539), .B(n22547), .Z(n22559) );
  XOR U24821 ( .A(n24862), .B(n24863), .Z(n22547) );
  XNOR U24822 ( .A(n24864), .B(n24774), .Z(n24863) );
  XNOR U24823 ( .A(n24865), .B(n24866), .Z(n24774) );
  XNOR U24824 ( .A(n24867), .B(n24868), .Z(n24866) );
  OR U24825 ( .A(n24869), .B(n24870), .Z(n24868) );
  XNOR U24826 ( .A(n24871), .B(n24872), .Z(n24862) );
  XOR U24827 ( .A(n24810), .B(n24873), .Z(n24872) );
  ANDN U24828 ( .B(n24874), .A(n24875), .Z(n24873) );
  ANDN U24829 ( .B(n24876), .A(n24877), .Z(n24810) );
  XOR U24830 ( .A(n24798), .B(n23298), .Z(n23274) );
  IV U24831 ( .A(n24757), .Z(n23298) );
  XOR U24832 ( .A(n24878), .B(n24841), .Z(n24757) );
  XNOR U24833 ( .A(n24663), .B(n24744), .Z(n24813) );
  XOR U24834 ( .A(n24879), .B(n24880), .Z(n24744) );
  XNOR U24835 ( .A(n21514), .B(n24881), .Z(n24880) );
  XOR U24836 ( .A(n24749), .B(n22572), .Z(n24881) );
  XOR U24837 ( .A(n21516), .B(n23304), .Z(n22572) );
  XOR U24838 ( .A(n24882), .B(n24883), .Z(n23304) );
  XNOR U24839 ( .A(n24829), .B(n24806), .Z(n24883) );
  XNOR U24840 ( .A(n24884), .B(n24885), .Z(n24806) );
  XNOR U24841 ( .A(n24886), .B(n24856), .Z(n24885) );
  ANDN U24842 ( .B(n24887), .A(n24888), .Z(n24856) );
  NOR U24843 ( .A(n24889), .B(n24890), .Z(n24886) );
  IV U24844 ( .A(n24891), .Z(n24829) );
  XOR U24845 ( .A(n24831), .B(n24892), .Z(n24882) );
  XOR U24846 ( .A(n24893), .B(n24894), .Z(n21516) );
  XNOR U24847 ( .A(n24819), .B(n24778), .Z(n24894) );
  XNOR U24848 ( .A(n24895), .B(n24896), .Z(n24778) );
  XNOR U24849 ( .A(n24897), .B(n24790), .Z(n24896) );
  ANDN U24850 ( .B(n24898), .A(n24899), .Z(n24790) );
  NOR U24851 ( .A(n24900), .B(n24901), .Z(n24897) );
  IV U24852 ( .A(n24902), .Z(n24819) );
  XOR U24853 ( .A(n24826), .B(n24903), .Z(n24893) );
  XOR U24854 ( .A(n24904), .B(n24905), .Z(n24749) );
  XOR U24855 ( .A(n23300), .B(n21540), .Z(n24905) );
  XNOR U24856 ( .A(n24906), .B(n21513), .Z(n21540) );
  XNOR U24857 ( .A(n24902), .B(n24907), .Z(n21513) );
  XNOR U24858 ( .A(n24826), .B(n24777), .Z(n24907) );
  XOR U24859 ( .A(n24860), .B(n24903), .Z(n24777) );
  XOR U24860 ( .A(n24786), .B(n24908), .Z(n24903) );
  XNOR U24861 ( .A(n24909), .B(n24910), .Z(n24908) );
  NANDN U24862 ( .A(n24911), .B(n24912), .Z(n24910) );
  XNOR U24863 ( .A(n24909), .B(n24914), .Z(n24913) );
  NANDN U24864 ( .A(n24915), .B(n24825), .Z(n24914) );
  OR U24865 ( .A(n24916), .B(n24917), .Z(n24909) );
  XNOR U24866 ( .A(n24786), .B(n24918), .Z(n24895) );
  XNOR U24867 ( .A(n24919), .B(n24920), .Z(n24918) );
  NAND U24868 ( .A(n24921), .B(n24922), .Z(n24920) );
  XOR U24869 ( .A(n24923), .B(n24919), .Z(n24786) );
  NANDN U24870 ( .A(n24924), .B(n24925), .Z(n24919) );
  ANDN U24871 ( .B(n24926), .A(n24927), .Z(n24923) );
  XOR U24872 ( .A(n24928), .B(n24929), .Z(n24902) );
  XOR U24873 ( .A(n24930), .B(n24931), .Z(n24929) );
  NANDN U24874 ( .A(n24932), .B(n24792), .Z(n24931) );
  IV U24875 ( .A(n23319), .Z(n23300) );
  XOR U24876 ( .A(n24781), .B(n24933), .Z(n23319) );
  XOR U24877 ( .A(n24840), .B(n24841), .Z(n24933) );
  XOR U24878 ( .A(n24878), .B(n24934), .Z(n24781) );
  IV U24879 ( .A(n24935), .Z(n24878) );
  XNOR U24880 ( .A(n23309), .B(n24936), .Z(n24904) );
  XOR U24881 ( .A(key[281]), .B(n23308), .Z(n24936) );
  XNOR U24882 ( .A(n24842), .B(n23275), .Z(n21514) );
  XOR U24883 ( .A(n24854), .B(n23309), .Z(n23275) );
  XNOR U24884 ( .A(n23305), .B(n24938), .Z(n24879) );
  XNOR U24885 ( .A(key[283]), .B(n22571), .Z(n24938) );
  XNOR U24886 ( .A(n21539), .B(n22561), .Z(n22571) );
  XOR U24887 ( .A(n24864), .B(n23308), .Z(n22561) );
  IV U24888 ( .A(n22532), .Z(n23308) );
  XOR U24889 ( .A(n24762), .B(n24939), .Z(n22532) );
  XOR U24890 ( .A(n24939), .B(n24864), .Z(n21539) );
  XNOR U24891 ( .A(n24865), .B(n24940), .Z(n24864) );
  XNOR U24892 ( .A(n24941), .B(n24942), .Z(n24940) );
  NOR U24893 ( .A(n24943), .B(n24812), .Z(n24941) );
  XOR U24894 ( .A(n24944), .B(n24945), .Z(n24865) );
  XNOR U24895 ( .A(n24946), .B(n24947), .Z(n24945) );
  NAND U24896 ( .A(n24948), .B(n24949), .Z(n24947) );
  XOR U24897 ( .A(n24950), .B(n24951), .Z(n23305) );
  XOR U24898 ( .A(n24841), .B(n24780), .Z(n24951) );
  XNOR U24899 ( .A(n24952), .B(n24953), .Z(n24780) );
  XOR U24900 ( .A(n24954), .B(n24800), .Z(n24953) );
  NANDN U24901 ( .A(n24955), .B(n24956), .Z(n24800) );
  NOR U24902 ( .A(n24957), .B(n24958), .Z(n24954) );
  XOR U24903 ( .A(n24959), .B(n24960), .Z(n24841) );
  XNOR U24904 ( .A(n24961), .B(n24962), .Z(n24960) );
  NAND U24905 ( .A(n24963), .B(n24802), .Z(n24962) );
  XNOR U24906 ( .A(n24840), .B(n24934), .Z(n24950) );
  XOR U24907 ( .A(n24796), .B(n24964), .Z(n24934) );
  XNOR U24908 ( .A(n24965), .B(n24966), .Z(n24964) );
  NANDN U24909 ( .A(n24967), .B(n24968), .Z(n24966) );
  XNOR U24910 ( .A(n24952), .B(n24969), .Z(n24840) );
  XNOR U24911 ( .A(n24965), .B(n24970), .Z(n24969) );
  OR U24912 ( .A(n24838), .B(n24971), .Z(n24970) );
  OR U24913 ( .A(n24972), .B(n24973), .Z(n24965) );
  XNOR U24914 ( .A(n24796), .B(n24974), .Z(n24952) );
  XNOR U24915 ( .A(n24975), .B(n24976), .Z(n24974) );
  NAND U24916 ( .A(n24977), .B(n24978), .Z(n24976) );
  XOR U24917 ( .A(n24979), .B(n24975), .Z(n24796) );
  NANDN U24918 ( .A(n24980), .B(n24981), .Z(n24975) );
  AND U24919 ( .A(n24982), .B(n24983), .Z(n24979) );
  XNOR U24920 ( .A(n24984), .B(n24985), .Z(n24663) );
  XOR U24921 ( .A(n24906), .B(n21541), .Z(n24985) );
  XOR U24922 ( .A(n22577), .B(n22554), .Z(n21541) );
  XOR U24923 ( .A(n24935), .B(n24798), .Z(n22554) );
  XNOR U24924 ( .A(n24834), .B(n24986), .Z(n24798) );
  XOR U24925 ( .A(n24987), .B(n24961), .Z(n24986) );
  NANDN U24926 ( .A(n24988), .B(n24956), .Z(n24961) );
  XNOR U24927 ( .A(n24958), .B(n24802), .Z(n24956) );
  NOR U24928 ( .A(n24989), .B(n24958), .Z(n24987) );
  XNOR U24929 ( .A(n24959), .B(n24990), .Z(n24834) );
  XNOR U24930 ( .A(n24991), .B(n24992), .Z(n24990) );
  NAND U24931 ( .A(n24978), .B(n24993), .Z(n24992) );
  XNOR U24932 ( .A(n24959), .B(n24994), .Z(n24935) );
  XOR U24933 ( .A(n24995), .B(n24836), .Z(n24994) );
  OR U24934 ( .A(n24996), .B(n24972), .Z(n24836) );
  XNOR U24935 ( .A(n24838), .B(n24967), .Z(n24972) );
  NOR U24936 ( .A(n24997), .B(n24967), .Z(n24995) );
  XOR U24937 ( .A(n24998), .B(n24991), .Z(n24959) );
  OR U24938 ( .A(n24980), .B(n24999), .Z(n24991) );
  XNOR U24939 ( .A(n24982), .B(n24978), .Z(n24980) );
  XNOR U24940 ( .A(n24967), .B(n24802), .Z(n24978) );
  XOR U24941 ( .A(n25000), .B(n25001), .Z(n24802) );
  NANDN U24942 ( .A(n25002), .B(n25003), .Z(n25001) );
  XNOR U24943 ( .A(n25004), .B(n25005), .Z(n24967) );
  OR U24944 ( .A(n25002), .B(n25006), .Z(n25005) );
  ANDN U24945 ( .B(n24982), .A(n25007), .Z(n24998) );
  XOR U24946 ( .A(n24838), .B(n24958), .Z(n24982) );
  XOR U24947 ( .A(n25008), .B(n25000), .Z(n24958) );
  NANDN U24948 ( .A(n25009), .B(n25010), .Z(n25000) );
  ANDN U24949 ( .B(n25011), .A(n25012), .Z(n25008) );
  NANDN U24950 ( .A(n25009), .B(n25014), .Z(n25004) );
  XOR U24951 ( .A(n25015), .B(n25002), .Z(n25009) );
  XNOR U24952 ( .A(n25016), .B(n25017), .Z(n25002) );
  XOR U24953 ( .A(n25018), .B(n25011), .Z(n25017) );
  XNOR U24954 ( .A(n25019), .B(n25020), .Z(n25016) );
  XNOR U24955 ( .A(n25021), .B(n25022), .Z(n25020) );
  ANDN U24956 ( .B(n25011), .A(n25023), .Z(n25021) );
  IV U24957 ( .A(n25024), .Z(n25011) );
  ANDN U24958 ( .B(n25015), .A(n25023), .Z(n25013) );
  IV U24959 ( .A(n25019), .Z(n25023) );
  IV U24960 ( .A(n25012), .Z(n25015) );
  XNOR U24961 ( .A(n25018), .B(n25025), .Z(n25012) );
  XOR U24962 ( .A(n25026), .B(n25022), .Z(n25025) );
  NAND U24963 ( .A(n25014), .B(n25010), .Z(n25022) );
  XNOR U24964 ( .A(n25003), .B(n25024), .Z(n25010) );
  XOR U24965 ( .A(n25027), .B(n25028), .Z(n25024) );
  XOR U24966 ( .A(n25029), .B(n25030), .Z(n25028) );
  XNOR U24967 ( .A(n24968), .B(n25031), .Z(n25030) );
  XNOR U24968 ( .A(n25032), .B(n25033), .Z(n25027) );
  XNOR U24969 ( .A(n25034), .B(n25035), .Z(n25033) );
  ANDN U24970 ( .B(n25036), .A(n24839), .Z(n25034) );
  XNOR U24971 ( .A(n25019), .B(n25006), .Z(n25014) );
  XOR U24972 ( .A(n25037), .B(n25038), .Z(n25019) );
  XNOR U24973 ( .A(n25039), .B(n25031), .Z(n25038) );
  XOR U24974 ( .A(n25040), .B(n25041), .Z(n25031) );
  XNOR U24975 ( .A(n25042), .B(n25043), .Z(n25041) );
  NAND U24976 ( .A(n24993), .B(n24977), .Z(n25043) );
  XNOR U24977 ( .A(n25044), .B(n25045), .Z(n25037) );
  ANDN U24978 ( .B(n25046), .A(n24989), .Z(n25044) );
  ANDN U24979 ( .B(n25003), .A(n25006), .Z(n25026) );
  XOR U24980 ( .A(n25006), .B(n25003), .Z(n25018) );
  XNOR U24981 ( .A(n25047), .B(n25048), .Z(n25003) );
  XNOR U24982 ( .A(n25040), .B(n25049), .Z(n25048) );
  XOR U24983 ( .A(n25039), .B(n24971), .Z(n25049) );
  XOR U24984 ( .A(n24839), .B(n25050), .Z(n25047) );
  XNOR U24985 ( .A(n25051), .B(n25035), .Z(n25050) );
  OR U24986 ( .A(n24973), .B(n24996), .Z(n25035) );
  XNOR U24987 ( .A(n24839), .B(n24997), .Z(n24996) );
  XOR U24988 ( .A(n24971), .B(n24968), .Z(n24973) );
  ANDN U24989 ( .B(n24968), .A(n24997), .Z(n25051) );
  XOR U24990 ( .A(n25052), .B(n25053), .Z(n25006) );
  XOR U24991 ( .A(n25040), .B(n25029), .Z(n25053) );
  XOR U24992 ( .A(n24963), .B(n24803), .Z(n25029) );
  XOR U24993 ( .A(n25054), .B(n25042), .Z(n25040) );
  NANDN U24994 ( .A(n24999), .B(n24981), .Z(n25042) );
  XOR U24995 ( .A(n24983), .B(n24977), .Z(n24981) );
  XNOR U24996 ( .A(n25046), .B(n25055), .Z(n24968) );
  XNOR U24997 ( .A(n25056), .B(n25057), .Z(n25055) );
  XOR U24998 ( .A(n25007), .B(n24993), .Z(n24999) );
  XNOR U24999 ( .A(n24997), .B(n24963), .Z(n24993) );
  IV U25000 ( .A(n25032), .Z(n24997) );
  XOR U25001 ( .A(n25058), .B(n25059), .Z(n25032) );
  XOR U25002 ( .A(n25060), .B(n25061), .Z(n25059) );
  XNOR U25003 ( .A(n24839), .B(n25062), .Z(n25058) );
  ANDN U25004 ( .B(n24983), .A(n25007), .Z(n25054) );
  XNOR U25005 ( .A(n24839), .B(n24989), .Z(n25007) );
  XOR U25006 ( .A(n25046), .B(n25036), .Z(n24983) );
  IV U25007 ( .A(n24971), .Z(n25036) );
  XOR U25008 ( .A(n25063), .B(n25064), .Z(n24971) );
  XOR U25009 ( .A(n25065), .B(n25061), .Z(n25064) );
  XNOR U25010 ( .A(n25066), .B(n25067), .Z(n25061) );
  XOR U25011 ( .A(n25068), .B(n25069), .Z(n25067) );
  XOR U25012 ( .A(n25070), .B(n25071), .Z(n25066) );
  XNOR U25013 ( .A(key[164]), .B(n24633), .Z(n25071) );
  XOR U25014 ( .A(n25072), .B(n25073), .Z(n24633) );
  IV U25015 ( .A(n24957), .Z(n25046) );
  XOR U25016 ( .A(n25039), .B(n25074), .Z(n25052) );
  XNOR U25017 ( .A(n25075), .B(n25045), .Z(n25074) );
  OR U25018 ( .A(n24955), .B(n24988), .Z(n25045) );
  XNOR U25019 ( .A(n25076), .B(n24963), .Z(n24988) );
  XNOR U25020 ( .A(n24957), .B(n24803), .Z(n24955) );
  ANDN U25021 ( .B(n24963), .A(n24803), .Z(n25075) );
  XOR U25022 ( .A(n25063), .B(n25077), .Z(n24803) );
  XOR U25023 ( .A(n25056), .B(n25078), .Z(n25077) );
  XOR U25024 ( .A(n25065), .B(n25063), .Z(n24963) );
  XNOR U25025 ( .A(n24989), .B(n24957), .Z(n25039) );
  XOR U25026 ( .A(n25063), .B(n25079), .Z(n24957) );
  XNOR U25027 ( .A(n25065), .B(n25060), .Z(n25079) );
  XOR U25028 ( .A(n25080), .B(n25081), .Z(n25060) );
  XOR U25029 ( .A(n25082), .B(n25083), .Z(n25081) );
  XNOR U25030 ( .A(key[167]), .B(n24655), .Z(n25080) );
  XNOR U25031 ( .A(n25084), .B(n25085), .Z(n25063) );
  XOR U25032 ( .A(n25086), .B(n25087), .Z(n25085) );
  XNOR U25033 ( .A(key[165]), .B(n25088), .Z(n25084) );
  IV U25034 ( .A(n25076), .Z(n24989) );
  XNOR U25035 ( .A(n25057), .B(n25089), .Z(n25076) );
  XOR U25036 ( .A(n25062), .B(n25078), .Z(n25089) );
  IV U25037 ( .A(n25065), .Z(n25078) );
  XOR U25038 ( .A(n25090), .B(n25091), .Z(n25065) );
  XOR U25039 ( .A(n24839), .B(n25092), .Z(n25091) );
  XNOR U25040 ( .A(n25093), .B(n25094), .Z(n24839) );
  XNOR U25041 ( .A(n25095), .B(n24643), .Z(n25094) );
  XOR U25042 ( .A(key[160]), .B(n24657), .Z(n25093) );
  XOR U25043 ( .A(n25096), .B(n25097), .Z(n25090) );
  XNOR U25044 ( .A(key[166]), .B(n24613), .Z(n25097) );
  XOR U25045 ( .A(n25072), .B(n25098), .Z(n24613) );
  XOR U25046 ( .A(n25099), .B(n25100), .Z(n25062) );
  XNOR U25047 ( .A(n25101), .B(n25102), .Z(n25100) );
  XOR U25048 ( .A(n25056), .B(n25103), .Z(n25102) );
  XOR U25049 ( .A(n25104), .B(n25105), .Z(n25056) );
  XOR U25050 ( .A(n24602), .B(n25106), .Z(n25105) );
  XOR U25051 ( .A(key[161]), .B(n25107), .Z(n25104) );
  XNOR U25052 ( .A(n25108), .B(n25109), .Z(n25099) );
  XNOR U25053 ( .A(key[163]), .B(n24648), .Z(n25109) );
  XOR U25054 ( .A(n25072), .B(n25110), .Z(n24648) );
  IV U25055 ( .A(n24655), .Z(n25072) );
  XOR U25056 ( .A(n25111), .B(n25112), .Z(n25057) );
  XNOR U25057 ( .A(n25113), .B(n25114), .Z(n25112) );
  XOR U25058 ( .A(key[162]), .B(n24640), .Z(n25111) );
  XOR U25059 ( .A(n24788), .B(n24860), .Z(n22577) );
  XOR U25060 ( .A(n24928), .B(n25115), .Z(n24860) );
  XOR U25061 ( .A(n25116), .B(n24822), .Z(n25115) );
  OR U25062 ( .A(n25117), .B(n24916), .Z(n24822) );
  XNOR U25063 ( .A(n24825), .B(n24912), .Z(n24916) );
  ANDN U25064 ( .B(n24912), .A(n25118), .Z(n25116) );
  IV U25065 ( .A(n25119), .Z(n24928) );
  XNOR U25066 ( .A(n24820), .B(n25120), .Z(n24788) );
  XNOR U25067 ( .A(n25121), .B(n24930), .Z(n25120) );
  XNOR U25068 ( .A(n24901), .B(n24792), .Z(n24898) );
  ANDN U25069 ( .B(n25123), .A(n24901), .Z(n25121) );
  XOR U25070 ( .A(n25119), .B(n25124), .Z(n24820) );
  XNOR U25071 ( .A(n25125), .B(n25126), .Z(n25124) );
  NAND U25072 ( .A(n24922), .B(n25127), .Z(n25126) );
  XNOR U25073 ( .A(n25128), .B(n25125), .Z(n25119) );
  OR U25074 ( .A(n25129), .B(n24924), .Z(n25125) );
  XOR U25075 ( .A(n24927), .B(n24922), .Z(n24924) );
  XOR U25076 ( .A(n24912), .B(n24792), .Z(n24922) );
  XOR U25077 ( .A(n25130), .B(n25131), .Z(n24792) );
  NANDN U25078 ( .A(n25132), .B(n25133), .Z(n25131) );
  XOR U25079 ( .A(n25134), .B(n25135), .Z(n24912) );
  NANDN U25080 ( .A(n25132), .B(n25136), .Z(n25135) );
  NOR U25081 ( .A(n24927), .B(n25137), .Z(n25128) );
  XOR U25082 ( .A(n24901), .B(n24825), .Z(n24927) );
  XNOR U25083 ( .A(n25138), .B(n25134), .Z(n24825) );
  NANDN U25084 ( .A(n25139), .B(n25140), .Z(n25134) );
  XOR U25085 ( .A(n25136), .B(n25141), .Z(n25140) );
  ANDN U25086 ( .B(n25141), .A(n25142), .Z(n25138) );
  XOR U25087 ( .A(n25143), .B(n25130), .Z(n24901) );
  NANDN U25088 ( .A(n25139), .B(n25144), .Z(n25130) );
  XOR U25089 ( .A(n25145), .B(n25133), .Z(n25144) );
  XNOR U25090 ( .A(n25146), .B(n25147), .Z(n25132) );
  XOR U25091 ( .A(n25148), .B(n25149), .Z(n25147) );
  XNOR U25092 ( .A(n25150), .B(n25151), .Z(n25146) );
  XNOR U25093 ( .A(n25152), .B(n25153), .Z(n25151) );
  ANDN U25094 ( .B(n25145), .A(n25149), .Z(n25152) );
  ANDN U25095 ( .B(n25145), .A(n25142), .Z(n25143) );
  XNOR U25096 ( .A(n25148), .B(n25154), .Z(n25142) );
  XOR U25097 ( .A(n25155), .B(n25153), .Z(n25154) );
  NAND U25098 ( .A(n25156), .B(n25157), .Z(n25153) );
  XNOR U25099 ( .A(n25150), .B(n25133), .Z(n25157) );
  IV U25100 ( .A(n25145), .Z(n25150) );
  XNOR U25101 ( .A(n25136), .B(n25149), .Z(n25156) );
  IV U25102 ( .A(n25141), .Z(n25149) );
  XOR U25103 ( .A(n25158), .B(n25159), .Z(n25141) );
  XNOR U25104 ( .A(n25160), .B(n25161), .Z(n25159) );
  XNOR U25105 ( .A(n25162), .B(n25163), .Z(n25158) );
  ANDN U25106 ( .B(n25123), .A(n24900), .Z(n25162) );
  AND U25107 ( .A(n25133), .B(n25136), .Z(n25155) );
  XNOR U25108 ( .A(n25133), .B(n25136), .Z(n25148) );
  XNOR U25109 ( .A(n25164), .B(n25165), .Z(n25136) );
  XNOR U25110 ( .A(n25166), .B(n25161), .Z(n25165) );
  XOR U25111 ( .A(n25167), .B(n25168), .Z(n25164) );
  XNOR U25112 ( .A(n25169), .B(n25163), .Z(n25168) );
  OR U25113 ( .A(n24899), .B(n25122), .Z(n25163) );
  XNOR U25114 ( .A(n25123), .B(n25170), .Z(n25122) );
  XNOR U25115 ( .A(n24900), .B(n24793), .Z(n24899) );
  ANDN U25116 ( .B(n25171), .A(n24932), .Z(n25169) );
  XNOR U25117 ( .A(n25172), .B(n25173), .Z(n25133) );
  XNOR U25118 ( .A(n25161), .B(n25174), .Z(n25173) );
  XOR U25119 ( .A(n24915), .B(n25167), .Z(n25174) );
  XNOR U25120 ( .A(n25123), .B(n24900), .Z(n25161) );
  XOR U25121 ( .A(n24824), .B(n25175), .Z(n25172) );
  XNOR U25122 ( .A(n25176), .B(n25177), .Z(n25175) );
  ANDN U25123 ( .B(n25178), .A(n25118), .Z(n25176) );
  XNOR U25124 ( .A(n25179), .B(n25180), .Z(n25145) );
  XNOR U25125 ( .A(n25166), .B(n25181), .Z(n25180) );
  XNOR U25126 ( .A(n24911), .B(n25160), .Z(n25181) );
  XOR U25127 ( .A(n25167), .B(n25182), .Z(n25160) );
  XNOR U25128 ( .A(n25183), .B(n25184), .Z(n25182) );
  NAND U25129 ( .A(n25127), .B(n24921), .Z(n25184) );
  XNOR U25130 ( .A(n25185), .B(n25183), .Z(n25167) );
  NANDN U25131 ( .A(n25129), .B(n24925), .Z(n25183) );
  XOR U25132 ( .A(n24926), .B(n24921), .Z(n24925) );
  XNOR U25133 ( .A(n25178), .B(n24793), .Z(n24921) );
  XOR U25134 ( .A(n25137), .B(n25127), .Z(n25129) );
  XNOR U25135 ( .A(n25118), .B(n25170), .Z(n25127) );
  ANDN U25136 ( .B(n24926), .A(n25137), .Z(n25185) );
  XOR U25137 ( .A(n24824), .B(n25123), .Z(n25137) );
  XNOR U25138 ( .A(n25186), .B(n25187), .Z(n25123) );
  XNOR U25139 ( .A(n25188), .B(n25189), .Z(n25187) );
  XOR U25140 ( .A(n25170), .B(n25171), .Z(n25166) );
  IV U25141 ( .A(n24793), .Z(n25171) );
  XOR U25142 ( .A(n25191), .B(n25192), .Z(n24793) );
  XOR U25143 ( .A(n25193), .B(n25189), .Z(n25192) );
  IV U25144 ( .A(n24932), .Z(n25170) );
  XOR U25145 ( .A(n25189), .B(n25194), .Z(n24932) );
  XNOR U25146 ( .A(n25195), .B(n25196), .Z(n25179) );
  XNOR U25147 ( .A(n25197), .B(n25177), .Z(n25196) );
  OR U25148 ( .A(n24917), .B(n25117), .Z(n25177) );
  XNOR U25149 ( .A(n24824), .B(n25118), .Z(n25117) );
  IV U25150 ( .A(n25195), .Z(n25118) );
  XOR U25151 ( .A(n24915), .B(n25178), .Z(n24917) );
  IV U25152 ( .A(n24911), .Z(n25178) );
  XOR U25153 ( .A(n25190), .B(n25198), .Z(n24911) );
  XNOR U25154 ( .A(n25199), .B(n25186), .Z(n25198) );
  XOR U25155 ( .A(n25200), .B(n25201), .Z(n25186) );
  XNOR U25156 ( .A(n25202), .B(n24187), .Z(n25201) );
  XOR U25157 ( .A(n24229), .B(n25203), .Z(n25200) );
  XNOR U25158 ( .A(key[202]), .B(n25204), .Z(n25203) );
  IV U25159 ( .A(n24900), .Z(n25190) );
  XOR U25160 ( .A(n25191), .B(n25205), .Z(n24900) );
  XOR U25161 ( .A(n25189), .B(n25206), .Z(n25205) );
  NOR U25162 ( .A(n24915), .B(n24824), .Z(n25197) );
  XOR U25163 ( .A(n25191), .B(n25207), .Z(n24915) );
  XOR U25164 ( .A(n25189), .B(n25208), .Z(n25207) );
  XOR U25165 ( .A(n25209), .B(n25210), .Z(n25189) );
  XNOR U25166 ( .A(n24824), .B(n25211), .Z(n25210) );
  XOR U25167 ( .A(n25212), .B(n25213), .Z(n25209) );
  XNOR U25168 ( .A(key[206]), .B(n24198), .Z(n25213) );
  XNOR U25169 ( .A(n25214), .B(n24209), .Z(n24198) );
  XOR U25170 ( .A(n25215), .B(n25216), .Z(n24209) );
  IV U25171 ( .A(n25194), .Z(n25191) );
  XOR U25172 ( .A(n25217), .B(n25218), .Z(n25194) );
  XOR U25173 ( .A(n25219), .B(n24202), .Z(n25218) );
  XNOR U25174 ( .A(n25222), .B(n25223), .Z(n25217) );
  XOR U25175 ( .A(key[205]), .B(n25224), .Z(n25223) );
  XOR U25176 ( .A(n25225), .B(n25226), .Z(n25195) );
  XNOR U25177 ( .A(n25208), .B(n25206), .Z(n25226) );
  XNOR U25178 ( .A(n25227), .B(n25228), .Z(n25206) );
  XOR U25179 ( .A(n25229), .B(n24210), .Z(n25228) );
  XNOR U25180 ( .A(n25230), .B(n25231), .Z(n24210) );
  XOR U25181 ( .A(key[207]), .B(n24234), .Z(n25227) );
  XNOR U25182 ( .A(n25232), .B(n25233), .Z(n25208) );
  XNOR U25183 ( .A(n24214), .B(n25234), .Z(n25233) );
  XOR U25184 ( .A(n25235), .B(n25236), .Z(n24214) );
  XNOR U25185 ( .A(n24216), .B(n25237), .Z(n25232) );
  XOR U25186 ( .A(key[204]), .B(n25238), .Z(n25237) );
  XOR U25187 ( .A(n25215), .B(n24204), .Z(n24216) );
  XNOR U25188 ( .A(n24824), .B(n25188), .Z(n25225) );
  XOR U25189 ( .A(n25239), .B(n25240), .Z(n25188) );
  XNOR U25190 ( .A(n25241), .B(n25242), .Z(n25240) );
  XOR U25191 ( .A(n25243), .B(n25199), .Z(n25242) );
  IV U25192 ( .A(n25193), .Z(n25199) );
  XNOR U25193 ( .A(n25244), .B(n25245), .Z(n25193) );
  XOR U25194 ( .A(n24189), .B(n25246), .Z(n25245) );
  XOR U25195 ( .A(n24226), .B(n25247), .Z(n25244) );
  XNOR U25196 ( .A(key[201]), .B(n25248), .Z(n25247) );
  XNOR U25197 ( .A(n24223), .B(n25249), .Z(n25239) );
  XNOR U25198 ( .A(key[203]), .B(n24231), .Z(n25249) );
  IV U25199 ( .A(n25250), .Z(n24231) );
  XOR U25200 ( .A(n25215), .B(n24218), .Z(n24223) );
  XNOR U25201 ( .A(n25251), .B(n25252), .Z(n24824) );
  XNOR U25202 ( .A(n25253), .B(n25254), .Z(n25252) );
  XNOR U25203 ( .A(n25255), .B(n25256), .Z(n25251) );
  XOR U25204 ( .A(key[200]), .B(n24228), .Z(n25256) );
  IV U25205 ( .A(n23302), .Z(n24906) );
  XOR U25206 ( .A(n24891), .B(n25257), .Z(n23302) );
  XNOR U25207 ( .A(n24831), .B(n24805), .Z(n25257) );
  XOR U25208 ( .A(n24937), .B(n24892), .Z(n24805) );
  XOR U25209 ( .A(n24847), .B(n25258), .Z(n24892) );
  XNOR U25210 ( .A(n25259), .B(n25260), .Z(n25258) );
  NANDN U25211 ( .A(n25261), .B(n25262), .Z(n25260) );
  XNOR U25212 ( .A(n25259), .B(n25264), .Z(n25263) );
  NANDN U25213 ( .A(n25265), .B(n24853), .Z(n25264) );
  OR U25214 ( .A(n25266), .B(n25267), .Z(n25259) );
  XNOR U25215 ( .A(n24847), .B(n25268), .Z(n24884) );
  XNOR U25216 ( .A(n25269), .B(n25270), .Z(n25268) );
  NAND U25217 ( .A(n25271), .B(n25272), .Z(n25270) );
  XOR U25218 ( .A(n25273), .B(n25269), .Z(n24847) );
  NANDN U25219 ( .A(n25274), .B(n25275), .Z(n25269) );
  ANDN U25220 ( .B(n25276), .A(n25277), .Z(n25273) );
  XOR U25221 ( .A(n25278), .B(n25279), .Z(n24891) );
  XOR U25222 ( .A(n25280), .B(n25281), .Z(n25279) );
  NANDN U25223 ( .A(n25282), .B(n24858), .Z(n25281) );
  XOR U25224 ( .A(n23299), .B(n25283), .Z(n24984) );
  XOR U25225 ( .A(key[280]), .B(n24842), .Z(n25283) );
  IV U25226 ( .A(n21533), .Z(n24842) );
  XOR U25227 ( .A(n24854), .B(n24937), .Z(n21533) );
  XOR U25228 ( .A(n25278), .B(n25284), .Z(n24937) );
  XOR U25229 ( .A(n25285), .B(n24850), .Z(n25284) );
  OR U25230 ( .A(n25286), .B(n25266), .Z(n24850) );
  XNOR U25231 ( .A(n24853), .B(n25262), .Z(n25266) );
  ANDN U25232 ( .B(n25262), .A(n25287), .Z(n25285) );
  IV U25233 ( .A(n25288), .Z(n25278) );
  XNOR U25234 ( .A(n24848), .B(n25289), .Z(n24854) );
  XNOR U25235 ( .A(n25290), .B(n25280), .Z(n25289) );
  XNOR U25236 ( .A(n24890), .B(n24858), .Z(n24887) );
  ANDN U25237 ( .B(n25292), .A(n24890), .Z(n25290) );
  XOR U25238 ( .A(n25288), .B(n25293), .Z(n24848) );
  XNOR U25239 ( .A(n25294), .B(n25295), .Z(n25293) );
  NAND U25240 ( .A(n25272), .B(n25296), .Z(n25295) );
  XNOR U25241 ( .A(n25297), .B(n25294), .Z(n25288) );
  OR U25242 ( .A(n25298), .B(n25274), .Z(n25294) );
  XOR U25243 ( .A(n25277), .B(n25272), .Z(n25274) );
  XOR U25244 ( .A(n25262), .B(n24858), .Z(n25272) );
  XOR U25245 ( .A(n25299), .B(n25300), .Z(n24858) );
  NANDN U25246 ( .A(n25301), .B(n25302), .Z(n25300) );
  XOR U25247 ( .A(n25303), .B(n25304), .Z(n25262) );
  NANDN U25248 ( .A(n25301), .B(n25305), .Z(n25304) );
  NOR U25249 ( .A(n25277), .B(n25306), .Z(n25297) );
  XOR U25250 ( .A(n24890), .B(n24853), .Z(n25277) );
  XNOR U25251 ( .A(n25307), .B(n25303), .Z(n24853) );
  NANDN U25252 ( .A(n25308), .B(n25309), .Z(n25303) );
  XOR U25253 ( .A(n25305), .B(n25310), .Z(n25309) );
  ANDN U25254 ( .B(n25310), .A(n25311), .Z(n25307) );
  XOR U25255 ( .A(n25312), .B(n25299), .Z(n24890) );
  NANDN U25256 ( .A(n25308), .B(n25313), .Z(n25299) );
  XOR U25257 ( .A(n25314), .B(n25302), .Z(n25313) );
  XNOR U25258 ( .A(n25315), .B(n25316), .Z(n25301) );
  XOR U25259 ( .A(n25317), .B(n25318), .Z(n25316) );
  XNOR U25260 ( .A(n25319), .B(n25320), .Z(n25315) );
  XNOR U25261 ( .A(n25321), .B(n25322), .Z(n25320) );
  ANDN U25262 ( .B(n25314), .A(n25318), .Z(n25321) );
  ANDN U25263 ( .B(n25314), .A(n25311), .Z(n25312) );
  XNOR U25264 ( .A(n25317), .B(n25323), .Z(n25311) );
  XOR U25265 ( .A(n25324), .B(n25322), .Z(n25323) );
  NAND U25266 ( .A(n25325), .B(n25326), .Z(n25322) );
  XNOR U25267 ( .A(n25319), .B(n25302), .Z(n25326) );
  IV U25268 ( .A(n25314), .Z(n25319) );
  XNOR U25269 ( .A(n25305), .B(n25318), .Z(n25325) );
  IV U25270 ( .A(n25310), .Z(n25318) );
  XOR U25271 ( .A(n25327), .B(n25328), .Z(n25310) );
  XNOR U25272 ( .A(n25329), .B(n25330), .Z(n25328) );
  XNOR U25273 ( .A(n25331), .B(n25332), .Z(n25327) );
  ANDN U25274 ( .B(n25292), .A(n24889), .Z(n25331) );
  AND U25275 ( .A(n25302), .B(n25305), .Z(n25324) );
  XNOR U25276 ( .A(n25302), .B(n25305), .Z(n25317) );
  XNOR U25277 ( .A(n25333), .B(n25334), .Z(n25305) );
  XNOR U25278 ( .A(n25335), .B(n25330), .Z(n25334) );
  XOR U25279 ( .A(n25336), .B(n25337), .Z(n25333) );
  XNOR U25280 ( .A(n25338), .B(n25332), .Z(n25337) );
  OR U25281 ( .A(n24888), .B(n25291), .Z(n25332) );
  XNOR U25282 ( .A(n25292), .B(n25339), .Z(n25291) );
  XNOR U25283 ( .A(n24889), .B(n24859), .Z(n24888) );
  ANDN U25284 ( .B(n25340), .A(n25282), .Z(n25338) );
  XNOR U25285 ( .A(n25341), .B(n25342), .Z(n25302) );
  XNOR U25286 ( .A(n25330), .B(n25343), .Z(n25342) );
  XOR U25287 ( .A(n25265), .B(n25336), .Z(n25343) );
  XNOR U25288 ( .A(n25292), .B(n24889), .Z(n25330) );
  XOR U25289 ( .A(n24852), .B(n25344), .Z(n25341) );
  XNOR U25290 ( .A(n25345), .B(n25346), .Z(n25344) );
  ANDN U25291 ( .B(n25347), .A(n25287), .Z(n25345) );
  XNOR U25292 ( .A(n25348), .B(n25349), .Z(n25314) );
  XNOR U25293 ( .A(n25335), .B(n25350), .Z(n25349) );
  XNOR U25294 ( .A(n25261), .B(n25329), .Z(n25350) );
  XOR U25295 ( .A(n25336), .B(n25351), .Z(n25329) );
  XNOR U25296 ( .A(n25352), .B(n25353), .Z(n25351) );
  NAND U25297 ( .A(n25296), .B(n25271), .Z(n25353) );
  XNOR U25298 ( .A(n25354), .B(n25352), .Z(n25336) );
  NANDN U25299 ( .A(n25298), .B(n25275), .Z(n25352) );
  XOR U25300 ( .A(n25276), .B(n25271), .Z(n25275) );
  XNOR U25301 ( .A(n25347), .B(n24859), .Z(n25271) );
  XOR U25302 ( .A(n25306), .B(n25296), .Z(n25298) );
  XNOR U25303 ( .A(n25287), .B(n25339), .Z(n25296) );
  ANDN U25304 ( .B(n25276), .A(n25306), .Z(n25354) );
  XOR U25305 ( .A(n24852), .B(n25292), .Z(n25306) );
  XNOR U25306 ( .A(n25355), .B(n25356), .Z(n25292) );
  XNOR U25307 ( .A(n25357), .B(n25358), .Z(n25356) );
  XOR U25308 ( .A(n25339), .B(n25340), .Z(n25335) );
  IV U25309 ( .A(n24859), .Z(n25340) );
  XOR U25310 ( .A(n25360), .B(n25361), .Z(n24859) );
  XNOR U25311 ( .A(n25362), .B(n25358), .Z(n25361) );
  IV U25312 ( .A(n25282), .Z(n25339) );
  XOR U25313 ( .A(n25358), .B(n25363), .Z(n25282) );
  XNOR U25314 ( .A(n25364), .B(n25365), .Z(n25348) );
  XNOR U25315 ( .A(n25366), .B(n25346), .Z(n25365) );
  OR U25316 ( .A(n25267), .B(n25286), .Z(n25346) );
  XNOR U25317 ( .A(n24852), .B(n25287), .Z(n25286) );
  IV U25318 ( .A(n25364), .Z(n25287) );
  XOR U25319 ( .A(n25265), .B(n25347), .Z(n25267) );
  IV U25320 ( .A(n25261), .Z(n25347) );
  XOR U25321 ( .A(n25359), .B(n25367), .Z(n25261) );
  XNOR U25322 ( .A(n25362), .B(n25355), .Z(n25367) );
  XOR U25323 ( .A(n25368), .B(n25369), .Z(n25355) );
  XNOR U25324 ( .A(n25370), .B(n25371), .Z(n25369) );
  XNOR U25325 ( .A(key[242]), .B(n25372), .Z(n25368) );
  IV U25326 ( .A(n24889), .Z(n25359) );
  XOR U25327 ( .A(n25360), .B(n25373), .Z(n24889) );
  XOR U25328 ( .A(n25358), .B(n25374), .Z(n25373) );
  NOR U25329 ( .A(n25265), .B(n24852), .Z(n25366) );
  XOR U25330 ( .A(n25360), .B(n25375), .Z(n25265) );
  XOR U25331 ( .A(n25358), .B(n25376), .Z(n25375) );
  XOR U25332 ( .A(n25377), .B(n25378), .Z(n25358) );
  XOR U25333 ( .A(n24852), .B(n25379), .Z(n25378) );
  XNOR U25334 ( .A(n25380), .B(n25381), .Z(n25377) );
  XNOR U25335 ( .A(key[246]), .B(n24345), .Z(n25381) );
  XOR U25336 ( .A(n24355), .B(n25382), .Z(n24345) );
  IV U25337 ( .A(n25363), .Z(n25360) );
  XOR U25338 ( .A(n25383), .B(n25384), .Z(n25363) );
  XOR U25339 ( .A(n25385), .B(n25386), .Z(n25384) );
  XOR U25340 ( .A(key[245]), .B(n25387), .Z(n25383) );
  XOR U25341 ( .A(n25388), .B(n25389), .Z(n25364) );
  XNOR U25342 ( .A(n25376), .B(n25374), .Z(n25389) );
  XNOR U25343 ( .A(n25390), .B(n25391), .Z(n25374) );
  XOR U25344 ( .A(n25392), .B(n25393), .Z(n25391) );
  XNOR U25345 ( .A(key[247]), .B(n25394), .Z(n25390) );
  XNOR U25346 ( .A(n25395), .B(n25396), .Z(n25376) );
  XOR U25347 ( .A(n25397), .B(n25398), .Z(n25396) );
  XOR U25348 ( .A(n25399), .B(n25400), .Z(n25395) );
  XNOR U25349 ( .A(key[244]), .B(n24323), .Z(n25400) );
  XOR U25350 ( .A(n24355), .B(n25401), .Z(n24323) );
  XNOR U25351 ( .A(n24852), .B(n25357), .Z(n25388) );
  XOR U25352 ( .A(n25402), .B(n25403), .Z(n25357) );
  XNOR U25353 ( .A(n25404), .B(n25405), .Z(n25403) );
  XOR U25354 ( .A(n25362), .B(n25406), .Z(n25405) );
  XOR U25355 ( .A(n25407), .B(n25408), .Z(n25362) );
  XOR U25356 ( .A(n24375), .B(n25409), .Z(n25408) );
  XNOR U25357 ( .A(key[241]), .B(n25410), .Z(n25407) );
  XOR U25358 ( .A(n25411), .B(n25412), .Z(n25402) );
  XNOR U25359 ( .A(key[243]), .B(n24368), .Z(n25412) );
  XOR U25360 ( .A(n24355), .B(n25413), .Z(n24368) );
  XNOR U25361 ( .A(n25414), .B(n25415), .Z(n24852) );
  XNOR U25362 ( .A(n25416), .B(n24363), .Z(n25415) );
  XNOR U25363 ( .A(key[240]), .B(n24353), .Z(n25414) );
  IV U25364 ( .A(n22569), .Z(n23299) );
  XNOR U25365 ( .A(n24762), .B(n24763), .Z(n25417) );
  IV U25366 ( .A(n24775), .Z(n24763) );
  XOR U25367 ( .A(n24807), .B(n25418), .Z(n24775) );
  XNOR U25368 ( .A(n25419), .B(n25420), .Z(n25418) );
  OR U25369 ( .A(n24869), .B(n25421), .Z(n25420) );
  XNOR U25370 ( .A(n24871), .B(n25422), .Z(n24807) );
  XNOR U25371 ( .A(n25423), .B(n25424), .Z(n25422) );
  NAND U25372 ( .A(n25425), .B(n24948), .Z(n25424) );
  XOR U25373 ( .A(n24942), .B(n25427), .Z(n25426) );
  NAND U25374 ( .A(n25428), .B(n24874), .Z(n25427) );
  XNOR U25375 ( .A(n24812), .B(n24874), .Z(n24876) );
  XNOR U25376 ( .A(n24939), .B(n24760), .Z(n24773) );
  XOR U25377 ( .A(n24871), .B(n25430), .Z(n24760) );
  XNOR U25378 ( .A(n25419), .B(n25431), .Z(n25430) );
  NANDN U25379 ( .A(n25432), .B(n25433), .Z(n25431) );
  OR U25380 ( .A(n25434), .B(n25435), .Z(n25419) );
  XOR U25381 ( .A(n25436), .B(n25423), .Z(n24871) );
  NANDN U25382 ( .A(n25437), .B(n25438), .Z(n25423) );
  AND U25383 ( .A(n25439), .B(n25440), .Z(n25436) );
  XNOR U25384 ( .A(n24944), .B(n25441), .Z(n24939) );
  XOR U25385 ( .A(n25442), .B(n24867), .Z(n25441) );
  OR U25386 ( .A(n25443), .B(n25434), .Z(n24867) );
  XNOR U25387 ( .A(n24869), .B(n25432), .Z(n25434) );
  NOR U25388 ( .A(n25444), .B(n25432), .Z(n25442) );
  XNOR U25389 ( .A(n25445), .B(n24946), .Z(n24944) );
  OR U25390 ( .A(n25437), .B(n25446), .Z(n24946) );
  XNOR U25391 ( .A(n25439), .B(n24948), .Z(n25437) );
  XNOR U25392 ( .A(n25432), .B(n24874), .Z(n24948) );
  XOR U25393 ( .A(n25447), .B(n25448), .Z(n24874) );
  NANDN U25394 ( .A(n25449), .B(n25450), .Z(n25448) );
  XNOR U25395 ( .A(n25451), .B(n25452), .Z(n25432) );
  OR U25396 ( .A(n25449), .B(n25453), .Z(n25452) );
  ANDN U25397 ( .B(n25439), .A(n25454), .Z(n25445) );
  XOR U25398 ( .A(n24869), .B(n24812), .Z(n25439) );
  XOR U25399 ( .A(n25455), .B(n25447), .Z(n24812) );
  NANDN U25400 ( .A(n25456), .B(n25457), .Z(n25447) );
  ANDN U25401 ( .B(n25458), .A(n25459), .Z(n25455) );
  NANDN U25402 ( .A(n25456), .B(n25461), .Z(n25451) );
  XOR U25403 ( .A(n25462), .B(n25449), .Z(n25456) );
  XNOR U25404 ( .A(n25463), .B(n25464), .Z(n25449) );
  XOR U25405 ( .A(n25465), .B(n25458), .Z(n25464) );
  XNOR U25406 ( .A(n25466), .B(n25467), .Z(n25463) );
  XNOR U25407 ( .A(n25468), .B(n25469), .Z(n25467) );
  ANDN U25408 ( .B(n25458), .A(n25470), .Z(n25468) );
  IV U25409 ( .A(n25471), .Z(n25458) );
  ANDN U25410 ( .B(n25462), .A(n25470), .Z(n25460) );
  IV U25411 ( .A(n25466), .Z(n25470) );
  IV U25412 ( .A(n25459), .Z(n25462) );
  XNOR U25413 ( .A(n25465), .B(n25472), .Z(n25459) );
  XOR U25414 ( .A(n25473), .B(n25469), .Z(n25472) );
  NAND U25415 ( .A(n25461), .B(n25457), .Z(n25469) );
  XNOR U25416 ( .A(n25450), .B(n25471), .Z(n25457) );
  XOR U25417 ( .A(n25474), .B(n25475), .Z(n25471) );
  XOR U25418 ( .A(n25476), .B(n25477), .Z(n25475) );
  XNOR U25419 ( .A(n25433), .B(n25478), .Z(n25477) );
  XNOR U25420 ( .A(n25479), .B(n25480), .Z(n25474) );
  XNOR U25421 ( .A(n25481), .B(n25482), .Z(n25480) );
  ANDN U25422 ( .B(n25483), .A(n24870), .Z(n25481) );
  XNOR U25423 ( .A(n25466), .B(n25453), .Z(n25461) );
  XOR U25424 ( .A(n25484), .B(n25485), .Z(n25466) );
  XNOR U25425 ( .A(n25486), .B(n25478), .Z(n25485) );
  XOR U25426 ( .A(n25487), .B(n25488), .Z(n25478) );
  XNOR U25427 ( .A(n25489), .B(n25490), .Z(n25488) );
  NAND U25428 ( .A(n24949), .B(n25425), .Z(n25490) );
  XNOR U25429 ( .A(n25491), .B(n25492), .Z(n25484) );
  ANDN U25430 ( .B(n25493), .A(n24943), .Z(n25491) );
  ANDN U25431 ( .B(n25450), .A(n25453), .Z(n25473) );
  XOR U25432 ( .A(n25453), .B(n25450), .Z(n25465) );
  XNOR U25433 ( .A(n25494), .B(n25495), .Z(n25450) );
  XNOR U25434 ( .A(n25487), .B(n25496), .Z(n25495) );
  XOR U25435 ( .A(n25486), .B(n25421), .Z(n25496) );
  XOR U25436 ( .A(n24870), .B(n25497), .Z(n25494) );
  XNOR U25437 ( .A(n25498), .B(n25482), .Z(n25497) );
  OR U25438 ( .A(n25435), .B(n25443), .Z(n25482) );
  XNOR U25439 ( .A(n24870), .B(n25444), .Z(n25443) );
  XOR U25440 ( .A(n25421), .B(n25433), .Z(n25435) );
  ANDN U25441 ( .B(n25433), .A(n25444), .Z(n25498) );
  XOR U25442 ( .A(n25499), .B(n25500), .Z(n25453) );
  XOR U25443 ( .A(n25487), .B(n25476), .Z(n25500) );
  XOR U25444 ( .A(n25428), .B(n24875), .Z(n25476) );
  XOR U25445 ( .A(n25501), .B(n25489), .Z(n25487) );
  NANDN U25446 ( .A(n25446), .B(n25438), .Z(n25489) );
  XOR U25447 ( .A(n25440), .B(n25425), .Z(n25438) );
  XNOR U25448 ( .A(n25493), .B(n25502), .Z(n25433) );
  XOR U25449 ( .A(n25503), .B(n25504), .Z(n25502) );
  XOR U25450 ( .A(n25454), .B(n24949), .Z(n25446) );
  XNOR U25451 ( .A(n25444), .B(n25428), .Z(n24949) );
  IV U25452 ( .A(n25479), .Z(n25444) );
  XOR U25453 ( .A(n25505), .B(n25506), .Z(n25479) );
  XOR U25454 ( .A(n25507), .B(n25508), .Z(n25506) );
  XNOR U25455 ( .A(n24870), .B(n25509), .Z(n25505) );
  ANDN U25456 ( .B(n25440), .A(n25454), .Z(n25501) );
  XNOR U25457 ( .A(n24870), .B(n24943), .Z(n25454) );
  XOR U25458 ( .A(n25493), .B(n25483), .Z(n25440) );
  IV U25459 ( .A(n25421), .Z(n25483) );
  XOR U25460 ( .A(n25510), .B(n25511), .Z(n25421) );
  XOR U25461 ( .A(n25512), .B(n25508), .Z(n25511) );
  XNOR U25462 ( .A(n25513), .B(n25514), .Z(n25508) );
  XOR U25463 ( .A(n24492), .B(n25515), .Z(n25514) );
  XOR U25464 ( .A(n25516), .B(n25517), .Z(n24492) );
  XNOR U25465 ( .A(n24491), .B(n25518), .Z(n25513) );
  XOR U25466 ( .A(key[156]), .B(n25519), .Z(n25518) );
  XNOR U25467 ( .A(n25520), .B(n24481), .Z(n24491) );
  IV U25468 ( .A(n24811), .Z(n25493) );
  XOR U25469 ( .A(n25486), .B(n25521), .Z(n25499) );
  XNOR U25470 ( .A(n25522), .B(n25492), .Z(n25521) );
  OR U25471 ( .A(n24877), .B(n25429), .Z(n25492) );
  XNOR U25472 ( .A(n25523), .B(n25428), .Z(n25429) );
  XNOR U25473 ( .A(n24811), .B(n24875), .Z(n24877) );
  ANDN U25474 ( .B(n25428), .A(n24875), .Z(n25522) );
  XOR U25475 ( .A(n25510), .B(n25524), .Z(n24875) );
  XNOR U25476 ( .A(n25525), .B(n25512), .Z(n25524) );
  XOR U25477 ( .A(n25512), .B(n25510), .Z(n25428) );
  XNOR U25478 ( .A(n24943), .B(n24811), .Z(n25486) );
  XOR U25479 ( .A(n25510), .B(n25526), .Z(n24811) );
  XNOR U25480 ( .A(n25512), .B(n25507), .Z(n25526) );
  XOR U25481 ( .A(n25527), .B(n25528), .Z(n25507) );
  XNOR U25482 ( .A(n25529), .B(n24487), .Z(n25528) );
  XOR U25483 ( .A(n25530), .B(n25531), .Z(n24487) );
  XOR U25484 ( .A(key[159]), .B(n24512), .Z(n25527) );
  XNOR U25485 ( .A(n25532), .B(n25533), .Z(n25510) );
  XOR U25486 ( .A(n25534), .B(n24479), .Z(n25533) );
  XNOR U25487 ( .A(n25535), .B(n25536), .Z(n24479) );
  XOR U25488 ( .A(n24473), .B(n25537), .Z(n25532) );
  XNOR U25489 ( .A(key[157]), .B(n25538), .Z(n25537) );
  IV U25490 ( .A(n25523), .Z(n24943) );
  XNOR U25491 ( .A(n25504), .B(n25539), .Z(n25523) );
  XOR U25492 ( .A(n25540), .B(n25541), .Z(n25512) );
  XOR U25493 ( .A(n24870), .B(n25542), .Z(n25541) );
  XNOR U25494 ( .A(n25543), .B(n25544), .Z(n24870) );
  XNOR U25495 ( .A(n25545), .B(n25546), .Z(n25544) );
  XNOR U25496 ( .A(n25547), .B(n25548), .Z(n25543) );
  XNOR U25497 ( .A(key[152]), .B(n25549), .Z(n25548) );
  XOR U25498 ( .A(n25550), .B(n25551), .Z(n25540) );
  XNOR U25499 ( .A(key[158]), .B(n24475), .Z(n25551) );
  XNOR U25500 ( .A(n25552), .B(n24486), .Z(n24475) );
  XOR U25501 ( .A(n25553), .B(n25554), .Z(n24486) );
  XOR U25502 ( .A(n25555), .B(n25556), .Z(n25509) );
  XNOR U25503 ( .A(n25557), .B(n25558), .Z(n25556) );
  XOR U25504 ( .A(n25559), .B(n25525), .Z(n25558) );
  IV U25505 ( .A(n25503), .Z(n25525) );
  XNOR U25506 ( .A(n25560), .B(n25561), .Z(n25503) );
  XNOR U25507 ( .A(n24503), .B(n25562), .Z(n25561) );
  XOR U25508 ( .A(n24466), .B(n25563), .Z(n25560) );
  XOR U25509 ( .A(key[153]), .B(n25564), .Z(n25563) );
  XNOR U25510 ( .A(n25565), .B(n25566), .Z(n25555) );
  XNOR U25511 ( .A(key[155]), .B(n24500), .Z(n25566) );
  XOR U25512 ( .A(n25553), .B(n24495), .Z(n24500) );
  XOR U25513 ( .A(n25567), .B(n25568), .Z(n25504) );
  XOR U25514 ( .A(n25569), .B(n24465), .Z(n25568) );
  XOR U25515 ( .A(n24506), .B(n25570), .Z(n25567) );
  XNOR U25516 ( .A(key[154]), .B(n25571), .Z(n25570) );
  XNOR U25517 ( .A(n25572), .B(n25573), .Z(n20014) );
  XOR U25518 ( .A(n25574), .B(n23678), .Z(n25573) );
  XNOR U25519 ( .A(n25575), .B(n25576), .Z(n23678) );
  XNOR U25520 ( .A(n25577), .B(n25578), .Z(n25576) );
  NANDN U25521 ( .A(n25579), .B(n23706), .Z(n25578) );
  XNOR U25522 ( .A(n23602), .B(n25580), .Z(n25572) );
  XOR U25523 ( .A(n25581), .B(n25582), .Z(n25580) );
  ANDN U25524 ( .B(n23701), .A(n25583), .Z(n25582) );
  XNOR U25525 ( .A(n25575), .B(n25584), .Z(n23602) );
  XNOR U25526 ( .A(n25585), .B(n23698), .Z(n25584) );
  ANDN U25527 ( .B(n25588), .A(n25589), .Z(n25585) );
  XNOR U25528 ( .A(n23696), .B(n25590), .Z(n25575) );
  XNOR U25529 ( .A(n25591), .B(n25592), .Z(n25590) );
  NANDN U25530 ( .A(n25593), .B(n25594), .Z(n25592) );
  XOR U25531 ( .A(n19414), .B(n25595), .Z(n23735) );
  XNOR U25532 ( .A(key[397]), .B(n20011), .Z(n25595) );
  XOR U25533 ( .A(n23679), .B(n23580), .Z(n20011) );
  XNOR U25534 ( .A(n23707), .B(n25596), .Z(n23580) );
  XNOR U25535 ( .A(n25597), .B(n25581), .Z(n25596) );
  ANDN U25536 ( .B(n25587), .A(n25598), .Z(n25581) );
  XOR U25537 ( .A(n25599), .B(n23701), .Z(n25587) );
  ANDN U25538 ( .B(n25600), .A(n25589), .Z(n25597) );
  IV U25539 ( .A(n25599), .Z(n25589) );
  XOR U25540 ( .A(n25574), .B(n25601), .Z(n23707) );
  XNOR U25541 ( .A(n25602), .B(n25603), .Z(n25601) );
  NANDN U25542 ( .A(n25593), .B(n25604), .Z(n25603) );
  XOR U25543 ( .A(n23603), .B(n23581), .Z(n23679) );
  XNOR U25544 ( .A(n23703), .B(n25606), .Z(n25605) );
  NANDN U25545 ( .A(n25607), .B(n25608), .Z(n25606) );
  OR U25546 ( .A(n25609), .B(n25610), .Z(n23703) );
  XNOR U25547 ( .A(n25611), .B(n25602), .Z(n25574) );
  NANDN U25548 ( .A(n25612), .B(n25613), .Z(n25602) );
  ANDN U25549 ( .B(n25614), .A(n25615), .Z(n25611) );
  XNOR U25550 ( .A(n23696), .B(n25616), .Z(n23603) );
  XOR U25551 ( .A(n25617), .B(n25577), .Z(n25616) );
  OR U25552 ( .A(n25618), .B(n25609), .Z(n25577) );
  XNOR U25553 ( .A(n23706), .B(n25608), .Z(n25609) );
  ANDN U25554 ( .B(n25608), .A(n25619), .Z(n25617) );
  XOR U25555 ( .A(n25620), .B(n25591), .Z(n23696) );
  OR U25556 ( .A(n25612), .B(n25621), .Z(n25591) );
  XNOR U25557 ( .A(n25615), .B(n25593), .Z(n25612) );
  XNOR U25558 ( .A(n25608), .B(n23701), .Z(n25593) );
  XOR U25559 ( .A(n25622), .B(n25623), .Z(n23701) );
  NANDN U25560 ( .A(n25624), .B(n25625), .Z(n25623) );
  XOR U25561 ( .A(n25626), .B(n25627), .Z(n25608) );
  NANDN U25562 ( .A(n25624), .B(n25628), .Z(n25627) );
  NOR U25563 ( .A(n25615), .B(n25629), .Z(n25620) );
  XNOR U25564 ( .A(n25599), .B(n23706), .Z(n25615) );
  XNOR U25565 ( .A(n25630), .B(n25626), .Z(n23706) );
  NANDN U25566 ( .A(n25631), .B(n25632), .Z(n25626) );
  XOR U25567 ( .A(n25628), .B(n25633), .Z(n25632) );
  ANDN U25568 ( .B(n25633), .A(n25634), .Z(n25630) );
  XNOR U25569 ( .A(n25635), .B(n25622), .Z(n25599) );
  NANDN U25570 ( .A(n25631), .B(n25636), .Z(n25622) );
  XOR U25571 ( .A(n25637), .B(n25625), .Z(n25636) );
  XNOR U25572 ( .A(n25638), .B(n25639), .Z(n25624) );
  XOR U25573 ( .A(n25640), .B(n25641), .Z(n25639) );
  XNOR U25574 ( .A(n25642), .B(n25643), .Z(n25638) );
  XNOR U25575 ( .A(n25644), .B(n25645), .Z(n25643) );
  ANDN U25576 ( .B(n25637), .A(n25641), .Z(n25644) );
  ANDN U25577 ( .B(n25637), .A(n25634), .Z(n25635) );
  XNOR U25578 ( .A(n25640), .B(n25646), .Z(n25634) );
  XOR U25579 ( .A(n25647), .B(n25645), .Z(n25646) );
  NAND U25580 ( .A(n25648), .B(n25649), .Z(n25645) );
  XNOR U25581 ( .A(n25642), .B(n25625), .Z(n25649) );
  IV U25582 ( .A(n25637), .Z(n25642) );
  XNOR U25583 ( .A(n25628), .B(n25641), .Z(n25648) );
  IV U25584 ( .A(n25633), .Z(n25641) );
  XOR U25585 ( .A(n25650), .B(n25651), .Z(n25633) );
  XNOR U25586 ( .A(n25652), .B(n25653), .Z(n25651) );
  XNOR U25587 ( .A(n25654), .B(n25655), .Z(n25650) );
  ANDN U25588 ( .B(n25588), .A(n25656), .Z(n25654) );
  AND U25589 ( .A(n25625), .B(n25628), .Z(n25647) );
  XNOR U25590 ( .A(n25625), .B(n25628), .Z(n25640) );
  XNOR U25591 ( .A(n25657), .B(n25658), .Z(n25628) );
  XNOR U25592 ( .A(n25659), .B(n25653), .Z(n25658) );
  XOR U25593 ( .A(n25660), .B(n25661), .Z(n25657) );
  XNOR U25594 ( .A(n25662), .B(n25655), .Z(n25661) );
  OR U25595 ( .A(n25598), .B(n25586), .Z(n25655) );
  XNOR U25596 ( .A(n25588), .B(n25663), .Z(n25586) );
  XNOR U25597 ( .A(n25656), .B(n25583), .Z(n25598) );
  ANDN U25598 ( .B(n25664), .A(n23700), .Z(n25662) );
  XNOR U25599 ( .A(n25665), .B(n25666), .Z(n25625) );
  XNOR U25600 ( .A(n25653), .B(n25667), .Z(n25666) );
  XOR U25601 ( .A(n23705), .B(n25660), .Z(n25667) );
  XNOR U25602 ( .A(n25588), .B(n25656), .Z(n25653) );
  XOR U25603 ( .A(n25579), .B(n25668), .Z(n25665) );
  XNOR U25604 ( .A(n25669), .B(n25670), .Z(n25668) );
  ANDN U25605 ( .B(n25671), .A(n25619), .Z(n25669) );
  XNOR U25606 ( .A(n25672), .B(n25673), .Z(n25637) );
  XNOR U25607 ( .A(n25659), .B(n25674), .Z(n25673) );
  XNOR U25608 ( .A(n25607), .B(n25652), .Z(n25674) );
  XOR U25609 ( .A(n25660), .B(n25675), .Z(n25652) );
  XNOR U25610 ( .A(n25676), .B(n25677), .Z(n25675) );
  NAND U25611 ( .A(n25594), .B(n25604), .Z(n25677) );
  XNOR U25612 ( .A(n25678), .B(n25676), .Z(n25660) );
  NANDN U25613 ( .A(n25621), .B(n25613), .Z(n25676) );
  XOR U25614 ( .A(n25614), .B(n25604), .Z(n25613) );
  XNOR U25615 ( .A(n25671), .B(n25583), .Z(n25604) );
  XOR U25616 ( .A(n25629), .B(n25594), .Z(n25621) );
  XNOR U25617 ( .A(n25619), .B(n25663), .Z(n25594) );
  ANDN U25618 ( .B(n25614), .A(n25629), .Z(n25678) );
  XOR U25619 ( .A(n25579), .B(n25588), .Z(n25629) );
  XNOR U25620 ( .A(n25679), .B(n25680), .Z(n25588) );
  XNOR U25621 ( .A(n25681), .B(n25682), .Z(n25680) );
  XOR U25622 ( .A(n25663), .B(n25664), .Z(n25659) );
  IV U25623 ( .A(n25583), .Z(n25664) );
  XOR U25624 ( .A(n25683), .B(n25684), .Z(n25583) );
  XNOR U25625 ( .A(n25685), .B(n25682), .Z(n25684) );
  IV U25626 ( .A(n23700), .Z(n25663) );
  XOR U25627 ( .A(n25682), .B(n25686), .Z(n23700) );
  XNOR U25628 ( .A(n25687), .B(n25688), .Z(n25672) );
  XNOR U25629 ( .A(n25689), .B(n25670), .Z(n25688) );
  OR U25630 ( .A(n25610), .B(n25618), .Z(n25670) );
  XNOR U25631 ( .A(n25579), .B(n25619), .Z(n25618) );
  IV U25632 ( .A(n25687), .Z(n25619) );
  XOR U25633 ( .A(n23705), .B(n25671), .Z(n25610) );
  IV U25634 ( .A(n25607), .Z(n25671) );
  XOR U25635 ( .A(n25600), .B(n25690), .Z(n25607) );
  XNOR U25636 ( .A(n25685), .B(n25679), .Z(n25690) );
  XOR U25637 ( .A(n25691), .B(n25692), .Z(n25679) );
  XNOR U25638 ( .A(n22100), .B(n21637), .Z(n25692) );
  IV U25639 ( .A(n23435), .Z(n21637) );
  XOR U25640 ( .A(n21680), .B(n22104), .Z(n23435) );
  XOR U25641 ( .A(n21640), .B(n21676), .Z(n22100) );
  XOR U25642 ( .A(n25693), .B(n25694), .Z(n21676) );
  XOR U25643 ( .A(n25695), .B(n25696), .Z(n25694) );
  XOR U25644 ( .A(n25697), .B(n25698), .Z(n25693) );
  XNOR U25645 ( .A(key[290]), .B(n21681), .Z(n25691) );
  IV U25646 ( .A(n25656), .Z(n25600) );
  XOR U25647 ( .A(n25683), .B(n25699), .Z(n25656) );
  XOR U25648 ( .A(n25682), .B(n25700), .Z(n25699) );
  NOR U25649 ( .A(n23705), .B(n25579), .Z(n25689) );
  XOR U25650 ( .A(n25683), .B(n25701), .Z(n23705) );
  XOR U25651 ( .A(n25682), .B(n25702), .Z(n25701) );
  XOR U25652 ( .A(n25703), .B(n25704), .Z(n25682) );
  XNOR U25653 ( .A(n22079), .B(n21650), .Z(n25704) );
  XOR U25654 ( .A(n23416), .B(n25705), .Z(n21650) );
  XNOR U25655 ( .A(n21655), .B(n22085), .Z(n23416) );
  XOR U25656 ( .A(n25706), .B(n25707), .Z(n22085) );
  XNOR U25657 ( .A(n25708), .B(n25709), .Z(n21655) );
  XOR U25658 ( .A(n22111), .B(n21662), .Z(n22079) );
  XNOR U25659 ( .A(n25710), .B(n25711), .Z(n21662) );
  XNOR U25660 ( .A(n25712), .B(n25713), .Z(n25711) );
  XNOR U25661 ( .A(n25714), .B(n25698), .Z(n25710) );
  XOR U25662 ( .A(n21657), .B(n25715), .Z(n25703) );
  XOR U25663 ( .A(key[294]), .B(n25579), .Z(n25715) );
  IV U25664 ( .A(n25686), .Z(n25683) );
  XOR U25665 ( .A(n25716), .B(n25717), .Z(n25686) );
  XNOR U25666 ( .A(n23408), .B(n21654), .Z(n25717) );
  XOR U25667 ( .A(n25718), .B(n25719), .Z(n22082) );
  XNOR U25668 ( .A(n25720), .B(n25721), .Z(n25719) );
  XOR U25669 ( .A(n25722), .B(n25723), .Z(n25718) );
  XOR U25670 ( .A(n25724), .B(n25725), .Z(n25723) );
  ANDN U25671 ( .B(n25726), .A(n25727), .Z(n25725) );
  XOR U25672 ( .A(n25728), .B(n25729), .Z(n23414) );
  XNOR U25673 ( .A(n25730), .B(n25731), .Z(n25729) );
  XNOR U25674 ( .A(n25732), .B(n25733), .Z(n25728) );
  XNOR U25675 ( .A(n25734), .B(n25735), .Z(n25733) );
  ANDN U25676 ( .B(n25736), .A(n25737), .Z(n25735) );
  XNOR U25677 ( .A(n21657), .B(n21648), .Z(n23408) );
  XOR U25678 ( .A(n25712), .B(n25696), .Z(n21648) );
  XNOR U25679 ( .A(n25738), .B(n25739), .Z(n25696) );
  XNOR U25680 ( .A(n25740), .B(n25741), .Z(n25739) );
  ANDN U25681 ( .B(n25742), .A(n25743), .Z(n25740) );
  XNOR U25682 ( .A(n25744), .B(n25745), .Z(n21657) );
  XOR U25683 ( .A(key[293]), .B(n23415), .Z(n25716) );
  XOR U25684 ( .A(n25746), .B(n25747), .Z(n25687) );
  XNOR U25685 ( .A(n25702), .B(n25700), .Z(n25747) );
  XNOR U25686 ( .A(n25748), .B(n25749), .Z(n25700) );
  XOR U25687 ( .A(n25705), .B(n21663), .Z(n25749) );
  XOR U25688 ( .A(n23423), .B(n22091), .Z(n21663) );
  XNOR U25689 ( .A(n25750), .B(n25751), .Z(n22091) );
  XOR U25690 ( .A(n25752), .B(n25721), .Z(n25751) );
  XNOR U25691 ( .A(n25753), .B(n25754), .Z(n25721) );
  XNOR U25692 ( .A(n25755), .B(n25756), .Z(n25754) );
  NANDN U25693 ( .A(n25757), .B(n25758), .Z(n25756) );
  XOR U25694 ( .A(n25759), .B(n25708), .Z(n25750) );
  XOR U25695 ( .A(n25760), .B(n25761), .Z(n23423) );
  XNOR U25696 ( .A(n25706), .B(n25731), .Z(n25761) );
  XNOR U25697 ( .A(n25762), .B(n25763), .Z(n25731) );
  XNOR U25698 ( .A(n25764), .B(n25765), .Z(n25763) );
  OR U25699 ( .A(n25766), .B(n25767), .Z(n25765) );
  XNOR U25700 ( .A(n23440), .B(n23421), .Z(n25705) );
  XNOR U25701 ( .A(n25768), .B(n25769), .Z(n23421) );
  XOR U25702 ( .A(n25770), .B(n25771), .Z(n25769) );
  XOR U25703 ( .A(n25772), .B(n25744), .Z(n25768) );
  XNOR U25704 ( .A(key[295]), .B(n22111), .Z(n25748) );
  XNOR U25705 ( .A(n25773), .B(n25774), .Z(n25702) );
  XNOR U25706 ( .A(n21669), .B(n21667), .Z(n25774) );
  XOR U25707 ( .A(n23429), .B(n22094), .Z(n21667) );
  XNOR U25708 ( .A(n25775), .B(n21680), .Z(n22094) );
  XOR U25709 ( .A(n25776), .B(n25752), .Z(n21680) );
  XNOR U25710 ( .A(n25732), .B(n22104), .Z(n23429) );
  XOR U25711 ( .A(n25777), .B(n25778), .Z(n22104) );
  XNOR U25712 ( .A(n25779), .B(n23415), .Z(n21669) );
  XNOR U25713 ( .A(n25780), .B(n25781), .Z(n23415) );
  XNOR U25714 ( .A(n25782), .B(n25771), .Z(n25781) );
  XNOR U25715 ( .A(n25783), .B(n25784), .Z(n25771) );
  XNOR U25716 ( .A(n25785), .B(n25786), .Z(n25784) );
  NANDN U25717 ( .A(n25787), .B(n25788), .Z(n25786) );
  XNOR U25718 ( .A(n25789), .B(n25790), .Z(n25780) );
  XOR U25719 ( .A(n25791), .B(n25792), .Z(n25790) );
  ANDN U25720 ( .B(n25793), .A(n25794), .Z(n25792) );
  XNOR U25721 ( .A(n22096), .B(n25795), .Z(n25773) );
  XOR U25722 ( .A(key[292]), .B(n23427), .Z(n25795) );
  XOR U25723 ( .A(n25796), .B(n21653), .Z(n22096) );
  XOR U25724 ( .A(n25797), .B(n25798), .Z(n21653) );
  XNOR U25725 ( .A(n25799), .B(n25713), .Z(n25798) );
  XNOR U25726 ( .A(n25800), .B(n25801), .Z(n25713) );
  XNOR U25727 ( .A(n25802), .B(n25803), .Z(n25801) );
  NANDN U25728 ( .A(n25804), .B(n25805), .Z(n25803) );
  XNOR U25729 ( .A(n25806), .B(n25807), .Z(n25797) );
  XOR U25730 ( .A(n25741), .B(n25808), .Z(n25807) );
  ANDN U25731 ( .B(n25809), .A(n25810), .Z(n25808) );
  ANDN U25732 ( .B(n25811), .A(n25812), .Z(n25741) );
  XNOR U25733 ( .A(n25579), .B(n25681), .Z(n25746) );
  XOR U25734 ( .A(n25813), .B(n25814), .Z(n25681) );
  XNOR U25735 ( .A(n25685), .B(n21686), .Z(n25815) );
  XOR U25736 ( .A(n23440), .B(n23427), .Z(n21686) );
  XOR U25737 ( .A(n25789), .B(n21681), .Z(n23427) );
  IV U25738 ( .A(n25816), .Z(n21681) );
  IV U25739 ( .A(n25779), .Z(n23440) );
  XOR U25740 ( .A(n25817), .B(n25818), .Z(n25685) );
  XOR U25741 ( .A(n22070), .B(n21679), .Z(n25818) );
  XOR U25742 ( .A(n22112), .B(n21689), .Z(n21679) );
  XNOR U25743 ( .A(n25752), .B(n25819), .Z(n21689) );
  XNOR U25744 ( .A(n25759), .B(n25708), .Z(n25819) );
  XNOR U25745 ( .A(n25776), .B(n25820), .Z(n25708) );
  XOR U25746 ( .A(n25706), .B(n25821), .Z(n22112) );
  XNOR U25747 ( .A(n25778), .B(n25822), .Z(n25821) );
  XNOR U25748 ( .A(n25777), .B(n25823), .Z(n25706) );
  XNOR U25749 ( .A(n21638), .B(n25816), .Z(n22070) );
  XNOR U25750 ( .A(n25824), .B(n25770), .Z(n25816) );
  XNOR U25751 ( .A(key[289]), .B(n21691), .Z(n25817) );
  XOR U25752 ( .A(n22068), .B(n21636), .Z(n21684) );
  XNOR U25753 ( .A(n25825), .B(n25826), .Z(n21636) );
  XOR U25754 ( .A(n25752), .B(n25709), .Z(n25826) );
  XNOR U25755 ( .A(n25827), .B(n25828), .Z(n25709) );
  XNOR U25756 ( .A(n25829), .B(n25724), .Z(n25828) );
  ANDN U25757 ( .B(n25830), .A(n25831), .Z(n25724) );
  ANDN U25758 ( .B(n25832), .A(n25833), .Z(n25829) );
  XOR U25759 ( .A(n25834), .B(n25835), .Z(n25752) );
  XOR U25760 ( .A(n25836), .B(n25837), .Z(n25835) );
  NANDN U25761 ( .A(n25838), .B(n25726), .Z(n25837) );
  XOR U25762 ( .A(n25759), .B(n25820), .Z(n25825) );
  XOR U25763 ( .A(n25720), .B(n25839), .Z(n25820) );
  XNOR U25764 ( .A(n25840), .B(n25841), .Z(n25839) );
  NANDN U25765 ( .A(n25842), .B(n25843), .Z(n25841) );
  XNOR U25766 ( .A(n25840), .B(n25845), .Z(n25844) );
  NANDN U25767 ( .A(n25846), .B(n25758), .Z(n25845) );
  OR U25768 ( .A(n25847), .B(n25848), .Z(n25840) );
  XNOR U25769 ( .A(n25720), .B(n25849), .Z(n25827) );
  XNOR U25770 ( .A(n25850), .B(n25851), .Z(n25849) );
  NANDN U25771 ( .A(n25852), .B(n25853), .Z(n25851) );
  XOR U25772 ( .A(n25854), .B(n25850), .Z(n25720) );
  NANDN U25773 ( .A(n25855), .B(n25856), .Z(n25850) );
  ANDN U25774 ( .B(n25857), .A(n25858), .Z(n25854) );
  IV U25775 ( .A(n23437), .Z(n22068) );
  XNOR U25776 ( .A(n25760), .B(n25859), .Z(n23437) );
  XOR U25777 ( .A(n25823), .B(n25707), .Z(n25859) );
  XNOR U25778 ( .A(n25860), .B(n25861), .Z(n25707) );
  XOR U25779 ( .A(n25862), .B(n25734), .Z(n25861) );
  NANDN U25780 ( .A(n25863), .B(n25864), .Z(n25734) );
  ANDN U25781 ( .B(n25865), .A(n25866), .Z(n25862) );
  XOR U25782 ( .A(n25730), .B(n25867), .Z(n25823) );
  XNOR U25783 ( .A(n25868), .B(n25869), .Z(n25867) );
  NANDN U25784 ( .A(n25870), .B(n25871), .Z(n25869) );
  XOR U25785 ( .A(n25778), .B(n25822), .Z(n25760) );
  XOR U25786 ( .A(n25860), .B(n25872), .Z(n25822) );
  XNOR U25787 ( .A(n25868), .B(n25873), .Z(n25872) );
  OR U25788 ( .A(n25766), .B(n25874), .Z(n25873) );
  OR U25789 ( .A(n25875), .B(n25876), .Z(n25868) );
  XNOR U25790 ( .A(n25730), .B(n25877), .Z(n25860) );
  XNOR U25791 ( .A(n25878), .B(n25879), .Z(n25877) );
  NANDN U25792 ( .A(n25880), .B(n25881), .Z(n25879) );
  XOR U25793 ( .A(n25882), .B(n25878), .Z(n25730) );
  NANDN U25794 ( .A(n25883), .B(n25884), .Z(n25878) );
  ANDN U25795 ( .B(n25885), .A(n25886), .Z(n25882) );
  XOR U25796 ( .A(n25887), .B(n25888), .Z(n25778) );
  XNOR U25797 ( .A(n25889), .B(n25890), .Z(n25888) );
  NAND U25798 ( .A(n25891), .B(n25736), .Z(n25890) );
  XNOR U25799 ( .A(n22108), .B(n25892), .Z(n25813) );
  XNOR U25800 ( .A(key[291]), .B(n21640), .Z(n25892) );
  XOR U25801 ( .A(n25893), .B(n25894), .Z(n21640) );
  XOR U25802 ( .A(n25770), .B(n25745), .Z(n25894) );
  XNOR U25803 ( .A(n25895), .B(n25896), .Z(n25745) );
  XNOR U25804 ( .A(n25897), .B(n25791), .Z(n25896) );
  ANDN U25805 ( .B(n25898), .A(n25899), .Z(n25791) );
  NOR U25806 ( .A(n25900), .B(n25901), .Z(n25897) );
  XNOR U25807 ( .A(n25772), .B(n25902), .Z(n25893) );
  XOR U25808 ( .A(n25796), .B(n21671), .Z(n22108) );
  XOR U25809 ( .A(n25799), .B(n21638), .Z(n21671) );
  XNOR U25810 ( .A(n25697), .B(n25903), .Z(n21638) );
  IV U25811 ( .A(n22111), .Z(n25796) );
  XNOR U25812 ( .A(n25903), .B(n25799), .Z(n22111) );
  XNOR U25813 ( .A(n25800), .B(n25904), .Z(n25799) );
  XOR U25814 ( .A(n25905), .B(n25906), .Z(n25904) );
  ANDN U25815 ( .B(n25907), .A(n25743), .Z(n25905) );
  IV U25816 ( .A(n25908), .Z(n25743) );
  XNOR U25817 ( .A(n25909), .B(n25910), .Z(n25800) );
  XNOR U25818 ( .A(n25911), .B(n25912), .Z(n25910) );
  NANDN U25819 ( .A(n25913), .B(n25914), .Z(n25912) );
  XNOR U25820 ( .A(n25915), .B(n25916), .Z(n25579) );
  XOR U25821 ( .A(n23422), .B(n22106), .Z(n25916) );
  XNOR U25822 ( .A(n21683), .B(n21691), .Z(n22106) );
  XOR U25823 ( .A(n25770), .B(n25917), .Z(n21691) );
  XNOR U25824 ( .A(n25772), .B(n25744), .Z(n25917) );
  XOR U25825 ( .A(n25824), .B(n25902), .Z(n25744) );
  XNOR U25826 ( .A(n25782), .B(n25918), .Z(n25902) );
  XNOR U25827 ( .A(n25919), .B(n25920), .Z(n25918) );
  NANDN U25828 ( .A(n25921), .B(n25922), .Z(n25920) );
  XNOR U25829 ( .A(n25919), .B(n25924), .Z(n25923) );
  NANDN U25830 ( .A(n25925), .B(n25788), .Z(n25924) );
  OR U25831 ( .A(n25926), .B(n25927), .Z(n25919) );
  XNOR U25832 ( .A(n25782), .B(n25928), .Z(n25895) );
  XNOR U25833 ( .A(n25929), .B(n25930), .Z(n25928) );
  NAND U25834 ( .A(n25931), .B(n25932), .Z(n25930) );
  XOR U25835 ( .A(n25933), .B(n25929), .Z(n25782) );
  NANDN U25836 ( .A(n25934), .B(n25935), .Z(n25929) );
  ANDN U25837 ( .B(n25936), .A(n25937), .Z(n25933) );
  XOR U25838 ( .A(n25938), .B(n25939), .Z(n25770) );
  XOR U25839 ( .A(n25940), .B(n25941), .Z(n25939) );
  NANDN U25840 ( .A(n25942), .B(n25793), .Z(n25941) );
  XOR U25841 ( .A(n25712), .B(n25943), .Z(n21683) );
  XOR U25842 ( .A(n25714), .B(n25698), .Z(n25943) );
  XOR U25843 ( .A(n25738), .B(n25944), .Z(n25698) );
  XNOR U25844 ( .A(n25945), .B(n25946), .Z(n25944) );
  NANDN U25845 ( .A(n25947), .B(n25805), .Z(n25946) );
  XNOR U25846 ( .A(n25806), .B(n25948), .Z(n25738) );
  XNOR U25847 ( .A(n25949), .B(n25950), .Z(n25948) );
  NANDN U25848 ( .A(n25913), .B(n25951), .Z(n25950) );
  IV U25849 ( .A(n25697), .Z(n25714) );
  XOR U25850 ( .A(n25909), .B(n25952), .Z(n25697) );
  XNOR U25851 ( .A(n25906), .B(n25953), .Z(n25952) );
  NANDN U25852 ( .A(n25954), .B(n25809), .Z(n25953) );
  XOR U25853 ( .A(n25908), .B(n25809), .Z(n25811) );
  XOR U25854 ( .A(n25903), .B(n25695), .Z(n25712) );
  XOR U25855 ( .A(n25806), .B(n25956), .Z(n25695) );
  XNOR U25856 ( .A(n25945), .B(n25957), .Z(n25956) );
  NANDN U25857 ( .A(n25958), .B(n25959), .Z(n25957) );
  OR U25858 ( .A(n25960), .B(n25961), .Z(n25945) );
  XOR U25859 ( .A(n25962), .B(n25949), .Z(n25806) );
  NANDN U25860 ( .A(n25963), .B(n25964), .Z(n25949) );
  ANDN U25861 ( .B(n25965), .A(n25966), .Z(n25962) );
  XNOR U25862 ( .A(n25909), .B(n25967), .Z(n25903) );
  XOR U25863 ( .A(n25968), .B(n25802), .Z(n25967) );
  OR U25864 ( .A(n25969), .B(n25960), .Z(n25802) );
  XNOR U25865 ( .A(n25805), .B(n25959), .Z(n25960) );
  ANDN U25866 ( .B(n25959), .A(n25970), .Z(n25968) );
  XOR U25867 ( .A(n25971), .B(n25911), .Z(n25909) );
  OR U25868 ( .A(n25963), .B(n25972), .Z(n25911) );
  XNOR U25869 ( .A(n25966), .B(n25913), .Z(n25963) );
  XNOR U25870 ( .A(n25959), .B(n25809), .Z(n25913) );
  XOR U25871 ( .A(n25973), .B(n25974), .Z(n25809) );
  NANDN U25872 ( .A(n25975), .B(n25976), .Z(n25974) );
  XOR U25873 ( .A(n25977), .B(n25978), .Z(n25959) );
  NANDN U25874 ( .A(n25975), .B(n25979), .Z(n25978) );
  NOR U25875 ( .A(n25966), .B(n25980), .Z(n25971) );
  XNOR U25876 ( .A(n25908), .B(n25805), .Z(n25966) );
  XNOR U25877 ( .A(n25981), .B(n25977), .Z(n25805) );
  NANDN U25878 ( .A(n25982), .B(n25983), .Z(n25977) );
  XOR U25879 ( .A(n25979), .B(n25984), .Z(n25983) );
  ANDN U25880 ( .B(n25984), .A(n25985), .Z(n25981) );
  XNOR U25881 ( .A(n25986), .B(n25973), .Z(n25908) );
  NANDN U25882 ( .A(n25982), .B(n25987), .Z(n25973) );
  XOR U25883 ( .A(n25988), .B(n25976), .Z(n25987) );
  XNOR U25884 ( .A(n25989), .B(n25990), .Z(n25975) );
  XOR U25885 ( .A(n25991), .B(n25992), .Z(n25990) );
  XNOR U25886 ( .A(n25993), .B(n25994), .Z(n25989) );
  XNOR U25887 ( .A(n25995), .B(n25996), .Z(n25994) );
  ANDN U25888 ( .B(n25988), .A(n25992), .Z(n25995) );
  ANDN U25889 ( .B(n25988), .A(n25985), .Z(n25986) );
  XNOR U25890 ( .A(n25991), .B(n25997), .Z(n25985) );
  XOR U25891 ( .A(n25998), .B(n25996), .Z(n25997) );
  NAND U25892 ( .A(n25999), .B(n26000), .Z(n25996) );
  XNOR U25893 ( .A(n25993), .B(n25976), .Z(n26000) );
  IV U25894 ( .A(n25988), .Z(n25993) );
  XNOR U25895 ( .A(n25979), .B(n25992), .Z(n25999) );
  IV U25896 ( .A(n25984), .Z(n25992) );
  XOR U25897 ( .A(n26001), .B(n26002), .Z(n25984) );
  XNOR U25898 ( .A(n26003), .B(n26004), .Z(n26002) );
  XNOR U25899 ( .A(n26005), .B(n26006), .Z(n26001) );
  ANDN U25900 ( .B(n25907), .A(n26007), .Z(n26005) );
  AND U25901 ( .A(n25976), .B(n25979), .Z(n25998) );
  XNOR U25902 ( .A(n25976), .B(n25979), .Z(n25991) );
  XNOR U25903 ( .A(n26008), .B(n26009), .Z(n25979) );
  XNOR U25904 ( .A(n26010), .B(n26004), .Z(n26009) );
  XOR U25905 ( .A(n26011), .B(n26012), .Z(n26008) );
  XNOR U25906 ( .A(n26013), .B(n26006), .Z(n26012) );
  OR U25907 ( .A(n25812), .B(n25955), .Z(n26006) );
  XNOR U25908 ( .A(n25907), .B(n26014), .Z(n25955) );
  XNOR U25909 ( .A(n26007), .B(n25810), .Z(n25812) );
  ANDN U25910 ( .B(n26015), .A(n25954), .Z(n26013) );
  XNOR U25911 ( .A(n26016), .B(n26017), .Z(n25976) );
  XNOR U25912 ( .A(n26004), .B(n26018), .Z(n26017) );
  XOR U25913 ( .A(n25947), .B(n26011), .Z(n26018) );
  XNOR U25914 ( .A(n25907), .B(n26007), .Z(n26004) );
  XOR U25915 ( .A(n25804), .B(n26019), .Z(n26016) );
  XNOR U25916 ( .A(n26020), .B(n26021), .Z(n26019) );
  ANDN U25917 ( .B(n26022), .A(n25970), .Z(n26020) );
  XNOR U25918 ( .A(n26023), .B(n26024), .Z(n25988) );
  XNOR U25919 ( .A(n26010), .B(n26025), .Z(n26024) );
  XNOR U25920 ( .A(n25958), .B(n26003), .Z(n26025) );
  XOR U25921 ( .A(n26011), .B(n26026), .Z(n26003) );
  XNOR U25922 ( .A(n26027), .B(n26028), .Z(n26026) );
  NAND U25923 ( .A(n25914), .B(n25951), .Z(n26028) );
  XNOR U25924 ( .A(n26029), .B(n26027), .Z(n26011) );
  NANDN U25925 ( .A(n25972), .B(n25964), .Z(n26027) );
  XOR U25926 ( .A(n25965), .B(n25951), .Z(n25964) );
  XNOR U25927 ( .A(n26022), .B(n25810), .Z(n25951) );
  XOR U25928 ( .A(n25980), .B(n25914), .Z(n25972) );
  XNOR U25929 ( .A(n25970), .B(n26014), .Z(n25914) );
  ANDN U25930 ( .B(n25965), .A(n25980), .Z(n26029) );
  XOR U25931 ( .A(n25804), .B(n25907), .Z(n25980) );
  XNOR U25932 ( .A(n26030), .B(n26031), .Z(n25907) );
  XNOR U25933 ( .A(n26032), .B(n26033), .Z(n26031) );
  XOR U25934 ( .A(n26014), .B(n26015), .Z(n26010) );
  IV U25935 ( .A(n25810), .Z(n26015) );
  XOR U25936 ( .A(n26034), .B(n26035), .Z(n25810) );
  XOR U25937 ( .A(n26036), .B(n26033), .Z(n26035) );
  IV U25938 ( .A(n25954), .Z(n26014) );
  XOR U25939 ( .A(n26033), .B(n26037), .Z(n25954) );
  XNOR U25940 ( .A(n26038), .B(n26039), .Z(n26023) );
  XNOR U25941 ( .A(n26040), .B(n26021), .Z(n26039) );
  OR U25942 ( .A(n25961), .B(n25969), .Z(n26021) );
  XNOR U25943 ( .A(n25804), .B(n25970), .Z(n25969) );
  IV U25944 ( .A(n26038), .Z(n25970) );
  XOR U25945 ( .A(n25947), .B(n26022), .Z(n25961) );
  IV U25946 ( .A(n25958), .Z(n26022) );
  XOR U25947 ( .A(n25742), .B(n26041), .Z(n25958) );
  XNOR U25948 ( .A(n26042), .B(n26030), .Z(n26041) );
  XOR U25949 ( .A(n26043), .B(n26044), .Z(n26030) );
  XNOR U25950 ( .A(n24227), .B(n26045), .Z(n26044) );
  XOR U25951 ( .A(key[194]), .B(n25250), .Z(n26043) );
  XOR U25952 ( .A(n26046), .B(n25204), .Z(n25250) );
  IV U25953 ( .A(n26007), .Z(n25742) );
  XOR U25954 ( .A(n26034), .B(n26047), .Z(n26007) );
  XOR U25955 ( .A(n26033), .B(n26048), .Z(n26047) );
  NOR U25956 ( .A(n25947), .B(n25804), .Z(n26040) );
  XOR U25957 ( .A(n26034), .B(n26049), .Z(n25947) );
  XOR U25958 ( .A(n26033), .B(n26050), .Z(n26049) );
  XOR U25959 ( .A(n26051), .B(n26052), .Z(n26033) );
  XNOR U25960 ( .A(n25804), .B(n26053), .Z(n26052) );
  XOR U25961 ( .A(n25211), .B(n26054), .Z(n26051) );
  XNOR U25962 ( .A(key[198]), .B(n26055), .Z(n26054) );
  XOR U25963 ( .A(n26056), .B(n25230), .Z(n25211) );
  IV U25964 ( .A(n26057), .Z(n25230) );
  IV U25965 ( .A(n26037), .Z(n26034) );
  XOR U25966 ( .A(n26058), .B(n26059), .Z(n26037) );
  XNOR U25967 ( .A(n25221), .B(n26060), .Z(n26059) );
  XNOR U25968 ( .A(key[197]), .B(n25214), .Z(n26058) );
  XOR U25969 ( .A(n25224), .B(n26055), .Z(n25214) );
  XOR U25970 ( .A(n26061), .B(n26062), .Z(n26038) );
  XNOR U25971 ( .A(n26050), .B(n26048), .Z(n26062) );
  XNOR U25972 ( .A(n26063), .B(n26064), .Z(n26048) );
  XOR U25973 ( .A(n26065), .B(n26066), .Z(n26064) );
  XOR U25974 ( .A(key[199]), .B(n26056), .Z(n26063) );
  XNOR U25975 ( .A(n26067), .B(n26068), .Z(n26050) );
  XNOR U25976 ( .A(n25234), .B(n26069), .Z(n26067) );
  XOR U25977 ( .A(key[196]), .B(n25235), .Z(n26069) );
  XNOR U25978 ( .A(n26056), .B(n25220), .Z(n25234) );
  XNOR U25979 ( .A(n25804), .B(n26032), .Z(n26061) );
  XOR U25980 ( .A(n26070), .B(n26071), .Z(n26032) );
  XOR U25981 ( .A(n26072), .B(n26073), .Z(n26071) );
  XNOR U25982 ( .A(n25241), .B(n26042), .Z(n26073) );
  IV U25983 ( .A(n26036), .Z(n26042) );
  XNOR U25984 ( .A(n26074), .B(n26075), .Z(n26036) );
  XOR U25985 ( .A(n26076), .B(n24187), .Z(n26075) );
  XOR U25986 ( .A(n26045), .B(n25246), .Z(n24187) );
  XOR U25987 ( .A(key[193]), .B(n24235), .Z(n26074) );
  XNOR U25988 ( .A(n25255), .B(n25236), .Z(n25241) );
  IV U25989 ( .A(n26056), .Z(n25255) );
  XOR U25990 ( .A(n26077), .B(n26078), .Z(n26070) );
  XNOR U25991 ( .A(key[195]), .B(n26046), .Z(n26078) );
  XNOR U25992 ( .A(n26079), .B(n26080), .Z(n25804) );
  XNOR U25993 ( .A(n24226), .B(n25254), .Z(n26080) );
  XOR U25994 ( .A(n26076), .B(n25253), .Z(n24226) );
  IV U25995 ( .A(n26081), .Z(n26076) );
  XNOR U25996 ( .A(key[192]), .B(n26082), .Z(n26079) );
  XOR U25997 ( .A(n25777), .B(n25732), .Z(n23422) );
  XNOR U25998 ( .A(n25762), .B(n26083), .Z(n25732) );
  XOR U25999 ( .A(n26084), .B(n25889), .Z(n26083) );
  NANDN U26000 ( .A(n26085), .B(n25864), .Z(n25889) );
  XOR U26001 ( .A(n25865), .B(n25736), .Z(n25864) );
  ANDN U26002 ( .B(n25865), .A(n26086), .Z(n26084) );
  XNOR U26003 ( .A(n25887), .B(n26087), .Z(n25762) );
  XNOR U26004 ( .A(n26088), .B(n26089), .Z(n26087) );
  NANDN U26005 ( .A(n25880), .B(n26090), .Z(n26089) );
  XOR U26006 ( .A(n25887), .B(n26091), .Z(n25777) );
  XOR U26007 ( .A(n26092), .B(n25764), .Z(n26091) );
  OR U26008 ( .A(n26093), .B(n25875), .Z(n25764) );
  XNOR U26009 ( .A(n25766), .B(n25870), .Z(n25875) );
  NOR U26010 ( .A(n26094), .B(n25870), .Z(n26092) );
  XOR U26011 ( .A(n26095), .B(n26088), .Z(n25887) );
  OR U26012 ( .A(n25883), .B(n26096), .Z(n26088) );
  XOR U26013 ( .A(n26097), .B(n25880), .Z(n25883) );
  XOR U26014 ( .A(n25870), .B(n25736), .Z(n25880) );
  XOR U26015 ( .A(n26098), .B(n26099), .Z(n25736) );
  NANDN U26016 ( .A(n26100), .B(n26101), .Z(n26099) );
  XNOR U26017 ( .A(n26102), .B(n26103), .Z(n25870) );
  OR U26018 ( .A(n26100), .B(n26104), .Z(n26103) );
  ANDN U26019 ( .B(n26097), .A(n26105), .Z(n26095) );
  IV U26020 ( .A(n25886), .Z(n26097) );
  XOR U26021 ( .A(n25766), .B(n25865), .Z(n25886) );
  XNOR U26022 ( .A(n26106), .B(n26098), .Z(n25865) );
  NANDN U26023 ( .A(n26107), .B(n26108), .Z(n26098) );
  ANDN U26024 ( .B(n26109), .A(n26110), .Z(n26106) );
  NANDN U26025 ( .A(n26107), .B(n26112), .Z(n26102) );
  XOR U26026 ( .A(n26113), .B(n26100), .Z(n26107) );
  XNOR U26027 ( .A(n26114), .B(n26115), .Z(n26100) );
  XOR U26028 ( .A(n26116), .B(n26109), .Z(n26115) );
  XNOR U26029 ( .A(n26117), .B(n26118), .Z(n26114) );
  XNOR U26030 ( .A(n26119), .B(n26120), .Z(n26118) );
  ANDN U26031 ( .B(n26109), .A(n26121), .Z(n26119) );
  IV U26032 ( .A(n26122), .Z(n26109) );
  ANDN U26033 ( .B(n26113), .A(n26121), .Z(n26111) );
  IV U26034 ( .A(n26117), .Z(n26121) );
  IV U26035 ( .A(n26110), .Z(n26113) );
  XNOR U26036 ( .A(n26116), .B(n26123), .Z(n26110) );
  XOR U26037 ( .A(n26124), .B(n26120), .Z(n26123) );
  NAND U26038 ( .A(n26112), .B(n26108), .Z(n26120) );
  XNOR U26039 ( .A(n26101), .B(n26122), .Z(n26108) );
  XOR U26040 ( .A(n26125), .B(n26126), .Z(n26122) );
  XOR U26041 ( .A(n26127), .B(n26128), .Z(n26126) );
  XNOR U26042 ( .A(n25871), .B(n26129), .Z(n26128) );
  XNOR U26043 ( .A(n26130), .B(n26131), .Z(n26125) );
  XNOR U26044 ( .A(n26132), .B(n26133), .Z(n26131) );
  ANDN U26045 ( .B(n26134), .A(n25767), .Z(n26132) );
  XNOR U26046 ( .A(n26117), .B(n26104), .Z(n26112) );
  XOR U26047 ( .A(n26135), .B(n26136), .Z(n26117) );
  XNOR U26048 ( .A(n26137), .B(n26129), .Z(n26136) );
  XOR U26049 ( .A(n26138), .B(n26139), .Z(n26129) );
  XNOR U26050 ( .A(n26140), .B(n26141), .Z(n26139) );
  NAND U26051 ( .A(n26090), .B(n25881), .Z(n26141) );
  XNOR U26052 ( .A(n26142), .B(n26143), .Z(n26135) );
  ANDN U26053 ( .B(n26144), .A(n26086), .Z(n26142) );
  ANDN U26054 ( .B(n26101), .A(n26104), .Z(n26124) );
  XOR U26055 ( .A(n26104), .B(n26101), .Z(n26116) );
  XNOR U26056 ( .A(n26145), .B(n26146), .Z(n26101) );
  XNOR U26057 ( .A(n26138), .B(n26147), .Z(n26146) );
  XOR U26058 ( .A(n26137), .B(n25874), .Z(n26147) );
  XOR U26059 ( .A(n25767), .B(n26148), .Z(n26145) );
  XNOR U26060 ( .A(n26149), .B(n26133), .Z(n26148) );
  OR U26061 ( .A(n25876), .B(n26093), .Z(n26133) );
  XNOR U26062 ( .A(n25767), .B(n26094), .Z(n26093) );
  XOR U26063 ( .A(n25874), .B(n25871), .Z(n25876) );
  ANDN U26064 ( .B(n25871), .A(n26094), .Z(n26149) );
  XOR U26065 ( .A(n26150), .B(n26151), .Z(n26104) );
  XOR U26066 ( .A(n26138), .B(n26127), .Z(n26151) );
  XOR U26067 ( .A(n25891), .B(n25737), .Z(n26127) );
  XOR U26068 ( .A(n26152), .B(n26140), .Z(n26138) );
  NANDN U26069 ( .A(n26096), .B(n25884), .Z(n26140) );
  XOR U26070 ( .A(n25885), .B(n25881), .Z(n25884) );
  XNOR U26071 ( .A(n26144), .B(n26153), .Z(n25871) );
  XOR U26072 ( .A(n26154), .B(n26155), .Z(n26153) );
  XOR U26073 ( .A(n26105), .B(n26090), .Z(n26096) );
  XNOR U26074 ( .A(n26094), .B(n25891), .Z(n26090) );
  IV U26075 ( .A(n26130), .Z(n26094) );
  XOR U26076 ( .A(n26156), .B(n26157), .Z(n26130) );
  XOR U26077 ( .A(n26158), .B(n26159), .Z(n26157) );
  XNOR U26078 ( .A(n25767), .B(n26160), .Z(n26156) );
  ANDN U26079 ( .B(n25885), .A(n26105), .Z(n26152) );
  XNOR U26080 ( .A(n25767), .B(n26086), .Z(n26105) );
  XOR U26081 ( .A(n26144), .B(n26134), .Z(n25885) );
  IV U26082 ( .A(n25874), .Z(n26134) );
  XOR U26083 ( .A(n26161), .B(n26162), .Z(n25874) );
  XOR U26084 ( .A(n26163), .B(n26159), .Z(n26162) );
  XNOR U26085 ( .A(n26164), .B(n26165), .Z(n26159) );
  XNOR U26086 ( .A(n25398), .B(n26166), .Z(n26165) );
  XNOR U26087 ( .A(n26167), .B(n24319), .Z(n25398) );
  XNOR U26088 ( .A(n25397), .B(n26168), .Z(n26164) );
  XNOR U26089 ( .A(key[236]), .B(n25413), .Z(n26168) );
  XNOR U26090 ( .A(n26169), .B(n25385), .Z(n25397) );
  IV U26091 ( .A(n25866), .Z(n26144) );
  XOR U26092 ( .A(n26137), .B(n26170), .Z(n26150) );
  XNOR U26093 ( .A(n26171), .B(n26143), .Z(n26170) );
  OR U26094 ( .A(n25863), .B(n26085), .Z(n26143) );
  XNOR U26095 ( .A(n26172), .B(n25891), .Z(n26085) );
  XNOR U26096 ( .A(n25866), .B(n25737), .Z(n25863) );
  ANDN U26097 ( .B(n25891), .A(n25737), .Z(n26171) );
  XOR U26098 ( .A(n26161), .B(n26173), .Z(n25737) );
  XOR U26099 ( .A(n26163), .B(n26161), .Z(n25891) );
  XNOR U26100 ( .A(n26086), .B(n25866), .Z(n26137) );
  XOR U26101 ( .A(n26161), .B(n26174), .Z(n25866) );
  XNOR U26102 ( .A(n26163), .B(n26158), .Z(n26174) );
  XOR U26103 ( .A(n26175), .B(n26176), .Z(n26158) );
  XOR U26104 ( .A(n25382), .B(n25393), .Z(n26176) );
  XNOR U26105 ( .A(n26177), .B(n26178), .Z(n25393) );
  XOR U26106 ( .A(n26179), .B(n26180), .Z(n24353) );
  XNOR U26107 ( .A(n26181), .B(n26182), .Z(n26161) );
  XNOR U26108 ( .A(n26183), .B(n25386), .Z(n26182) );
  XOR U26109 ( .A(n26184), .B(n24339), .Z(n25386) );
  XOR U26110 ( .A(key[237]), .B(n24347), .Z(n26185) );
  IV U26111 ( .A(n26172), .Z(n26086) );
  XNOR U26112 ( .A(n26155), .B(n26186), .Z(n26172) );
  XOR U26113 ( .A(n26187), .B(n26188), .Z(n26163) );
  XOR U26114 ( .A(n25767), .B(n26189), .Z(n26188) );
  XNOR U26115 ( .A(n26190), .B(n26191), .Z(n25767) );
  XNOR U26116 ( .A(n24364), .B(n26192), .Z(n26191) );
  XOR U26117 ( .A(n26193), .B(n26194), .Z(n26190) );
  XNOR U26118 ( .A(key[232]), .B(n26180), .Z(n26194) );
  XNOR U26119 ( .A(n25379), .B(n26195), .Z(n26187) );
  XNOR U26120 ( .A(key[238]), .B(n24341), .Z(n26195) );
  XNOR U26121 ( .A(n26196), .B(n25392), .Z(n25379) );
  XOR U26122 ( .A(n26169), .B(n26197), .Z(n25392) );
  XOR U26123 ( .A(n26198), .B(n26199), .Z(n26160) );
  XOR U26124 ( .A(n26200), .B(n26201), .Z(n26199) );
  XOR U26125 ( .A(n25404), .B(n26154), .Z(n26201) );
  XNOR U26126 ( .A(n26202), .B(n26203), .Z(n26154) );
  XOR U26127 ( .A(n24374), .B(n25409), .Z(n26203) );
  XNOR U26128 ( .A(n25370), .B(n26204), .Z(n26202) );
  XOR U26129 ( .A(key[233]), .B(n26205), .Z(n26204) );
  XOR U26130 ( .A(n25406), .B(n26206), .Z(n26198) );
  XNOR U26131 ( .A(key[235]), .B(n24377), .Z(n26206) );
  XOR U26132 ( .A(n26179), .B(n25399), .Z(n25406) );
  XOR U26133 ( .A(n26207), .B(n26208), .Z(n26155) );
  XOR U26134 ( .A(n25411), .B(n25371), .Z(n26208) );
  XOR U26135 ( .A(n24360), .B(n26209), .Z(n26207) );
  XOR U26136 ( .A(key[234]), .B(n26210), .Z(n26209) );
  XNOR U26137 ( .A(n21693), .B(n25779), .Z(n21664) );
  XOR U26138 ( .A(n25789), .B(n25824), .Z(n25779) );
  XNOR U26139 ( .A(n25938), .B(n26211), .Z(n25824) );
  XOR U26140 ( .A(n26212), .B(n25785), .Z(n26211) );
  OR U26141 ( .A(n26213), .B(n25926), .Z(n25785) );
  XNOR U26142 ( .A(n25788), .B(n25922), .Z(n25926) );
  ANDN U26143 ( .B(n25922), .A(n26214), .Z(n26212) );
  IV U26144 ( .A(n26215), .Z(n25938) );
  XNOR U26145 ( .A(n25783), .B(n26216), .Z(n25789) );
  XNOR U26146 ( .A(n26217), .B(n25940), .Z(n26216) );
  XNOR U26147 ( .A(n25901), .B(n25793), .Z(n25898) );
  ANDN U26148 ( .B(n26219), .A(n25901), .Z(n26217) );
  XOR U26149 ( .A(n26215), .B(n26220), .Z(n25783) );
  XNOR U26150 ( .A(n26221), .B(n26222), .Z(n26220) );
  NAND U26151 ( .A(n25932), .B(n26223), .Z(n26222) );
  XNOR U26152 ( .A(n26224), .B(n26221), .Z(n26215) );
  OR U26153 ( .A(n25934), .B(n26225), .Z(n26221) );
  XNOR U26154 ( .A(n26226), .B(n25932), .Z(n25934) );
  XOR U26155 ( .A(n25922), .B(n25793), .Z(n25932) );
  XOR U26156 ( .A(n26227), .B(n26228), .Z(n25793) );
  NANDN U26157 ( .A(n26229), .B(n26230), .Z(n26228) );
  XOR U26158 ( .A(n26231), .B(n26232), .Z(n25922) );
  NANDN U26159 ( .A(n26229), .B(n26233), .Z(n26232) );
  ANDN U26160 ( .B(n26226), .A(n26234), .Z(n26224) );
  IV U26161 ( .A(n25937), .Z(n26226) );
  XOR U26162 ( .A(n25901), .B(n25788), .Z(n25937) );
  XNOR U26163 ( .A(n26235), .B(n26231), .Z(n25788) );
  NANDN U26164 ( .A(n26236), .B(n26237), .Z(n26231) );
  XOR U26165 ( .A(n26233), .B(n26238), .Z(n26237) );
  ANDN U26166 ( .B(n26238), .A(n26239), .Z(n26235) );
  XOR U26167 ( .A(n26240), .B(n26227), .Z(n25901) );
  NANDN U26168 ( .A(n26236), .B(n26241), .Z(n26227) );
  XOR U26169 ( .A(n26242), .B(n26230), .Z(n26241) );
  XNOR U26170 ( .A(n26243), .B(n26244), .Z(n26229) );
  XOR U26171 ( .A(n26245), .B(n26246), .Z(n26244) );
  XNOR U26172 ( .A(n26247), .B(n26248), .Z(n26243) );
  XNOR U26173 ( .A(n26249), .B(n26250), .Z(n26248) );
  ANDN U26174 ( .B(n26242), .A(n26246), .Z(n26249) );
  ANDN U26175 ( .B(n26242), .A(n26239), .Z(n26240) );
  XNOR U26176 ( .A(n26245), .B(n26251), .Z(n26239) );
  XOR U26177 ( .A(n26252), .B(n26250), .Z(n26251) );
  NAND U26178 ( .A(n26253), .B(n26254), .Z(n26250) );
  XNOR U26179 ( .A(n26247), .B(n26230), .Z(n26254) );
  IV U26180 ( .A(n26242), .Z(n26247) );
  XNOR U26181 ( .A(n26233), .B(n26246), .Z(n26253) );
  IV U26182 ( .A(n26238), .Z(n26246) );
  XOR U26183 ( .A(n26255), .B(n26256), .Z(n26238) );
  XNOR U26184 ( .A(n26257), .B(n26258), .Z(n26256) );
  XNOR U26185 ( .A(n26259), .B(n26260), .Z(n26255) );
  ANDN U26186 ( .B(n26219), .A(n25900), .Z(n26259) );
  AND U26187 ( .A(n26230), .B(n26233), .Z(n26252) );
  XNOR U26188 ( .A(n26230), .B(n26233), .Z(n26245) );
  XNOR U26189 ( .A(n26261), .B(n26262), .Z(n26233) );
  XNOR U26190 ( .A(n26263), .B(n26258), .Z(n26262) );
  XOR U26191 ( .A(n26264), .B(n26265), .Z(n26261) );
  XNOR U26192 ( .A(n26266), .B(n26260), .Z(n26265) );
  OR U26193 ( .A(n25899), .B(n26218), .Z(n26260) );
  XNOR U26194 ( .A(n26219), .B(n26267), .Z(n26218) );
  XNOR U26195 ( .A(n25900), .B(n25794), .Z(n25899) );
  ANDN U26196 ( .B(n26268), .A(n25942), .Z(n26266) );
  XNOR U26197 ( .A(n26269), .B(n26270), .Z(n26230) );
  XNOR U26198 ( .A(n26258), .B(n26271), .Z(n26270) );
  XOR U26199 ( .A(n25925), .B(n26264), .Z(n26271) );
  XNOR U26200 ( .A(n26219), .B(n25900), .Z(n26258) );
  XOR U26201 ( .A(n25787), .B(n26272), .Z(n26269) );
  XNOR U26202 ( .A(n26273), .B(n26274), .Z(n26272) );
  ANDN U26203 ( .B(n26275), .A(n26214), .Z(n26273) );
  XNOR U26204 ( .A(n26276), .B(n26277), .Z(n26242) );
  XNOR U26205 ( .A(n26263), .B(n26278), .Z(n26277) );
  XNOR U26206 ( .A(n25921), .B(n26257), .Z(n26278) );
  XOR U26207 ( .A(n26264), .B(n26279), .Z(n26257) );
  XNOR U26208 ( .A(n26280), .B(n26281), .Z(n26279) );
  NAND U26209 ( .A(n26223), .B(n25931), .Z(n26281) );
  XNOR U26210 ( .A(n26282), .B(n26280), .Z(n26264) );
  NANDN U26211 ( .A(n26225), .B(n25935), .Z(n26280) );
  XOR U26212 ( .A(n25936), .B(n25931), .Z(n25935) );
  XNOR U26213 ( .A(n26275), .B(n25794), .Z(n25931) );
  XOR U26214 ( .A(n26234), .B(n26223), .Z(n26225) );
  XNOR U26215 ( .A(n26214), .B(n26267), .Z(n26223) );
  ANDN U26216 ( .B(n25936), .A(n26234), .Z(n26282) );
  XOR U26217 ( .A(n25787), .B(n26219), .Z(n26234) );
  XNOR U26218 ( .A(n26283), .B(n26284), .Z(n26219) );
  XNOR U26219 ( .A(n26285), .B(n26286), .Z(n26284) );
  XOR U26220 ( .A(n26267), .B(n26268), .Z(n26263) );
  IV U26221 ( .A(n25794), .Z(n26268) );
  XOR U26222 ( .A(n26288), .B(n26289), .Z(n25794) );
  XOR U26223 ( .A(n26290), .B(n26286), .Z(n26289) );
  IV U26224 ( .A(n25942), .Z(n26267) );
  XOR U26225 ( .A(n26286), .B(n26291), .Z(n25942) );
  XNOR U26226 ( .A(n26292), .B(n26293), .Z(n26276) );
  XNOR U26227 ( .A(n26294), .B(n26274), .Z(n26293) );
  OR U26228 ( .A(n25927), .B(n26213), .Z(n26274) );
  XNOR U26229 ( .A(n25787), .B(n26214), .Z(n26213) );
  IV U26230 ( .A(n26292), .Z(n26214) );
  XOR U26231 ( .A(n25925), .B(n26275), .Z(n25927) );
  IV U26232 ( .A(n25921), .Z(n26275) );
  XOR U26233 ( .A(n26287), .B(n26295), .Z(n25921) );
  XOR U26234 ( .A(n26296), .B(n26297), .Z(n26283) );
  XNOR U26235 ( .A(n25108), .B(n26298), .Z(n26296) );
  XOR U26236 ( .A(key[186]), .B(n26299), .Z(n26298) );
  IV U26237 ( .A(n25900), .Z(n26287) );
  XOR U26238 ( .A(n26288), .B(n26300), .Z(n25900) );
  XOR U26239 ( .A(n26286), .B(n26301), .Z(n26300) );
  NOR U26240 ( .A(n25925), .B(n25787), .Z(n26294) );
  XOR U26241 ( .A(n26288), .B(n26302), .Z(n25925) );
  XOR U26242 ( .A(n26286), .B(n26303), .Z(n26302) );
  XOR U26243 ( .A(n26304), .B(n26305), .Z(n26286) );
  XOR U26244 ( .A(n25787), .B(n26306), .Z(n26305) );
  XNOR U26245 ( .A(n25092), .B(n26307), .Z(n26304) );
  XOR U26246 ( .A(key[190]), .B(n24621), .Z(n26307) );
  XNOR U26247 ( .A(n26308), .B(n25082), .Z(n25092) );
  XNOR U26248 ( .A(n26309), .B(n26310), .Z(n25082) );
  IV U26249 ( .A(n26291), .Z(n26288) );
  XOR U26250 ( .A(n26311), .B(n26312), .Z(n26291) );
  XOR U26251 ( .A(n25073), .B(n25087), .Z(n26312) );
  XOR U26252 ( .A(n26313), .B(n24618), .Z(n25087) );
  XOR U26253 ( .A(n25096), .B(n26314), .Z(n26311) );
  XOR U26254 ( .A(key[189]), .B(n24612), .Z(n26314) );
  XOR U26255 ( .A(n26315), .B(n26316), .Z(n26292) );
  XNOR U26256 ( .A(n26303), .B(n26301), .Z(n26316) );
  XNOR U26257 ( .A(n26317), .B(n26318), .Z(n26301) );
  XOR U26258 ( .A(n25098), .B(n25083), .Z(n26318) );
  XOR U26259 ( .A(n26319), .B(n24627), .Z(n25083) );
  XOR U26260 ( .A(key[191]), .B(n24657), .Z(n26317) );
  XOR U26261 ( .A(n26320), .B(n26309), .Z(n24657) );
  XNOR U26262 ( .A(n26321), .B(n26322), .Z(n26303) );
  XNOR U26263 ( .A(n25069), .B(n26323), .Z(n26322) );
  XNOR U26264 ( .A(n26324), .B(n24631), .Z(n25069) );
  XNOR U26265 ( .A(n25068), .B(n26325), .Z(n26321) );
  XNOR U26266 ( .A(key[188]), .B(n25110), .Z(n26325) );
  XNOR U26267 ( .A(n26309), .B(n26326), .Z(n25068) );
  XNOR U26268 ( .A(n25787), .B(n26285), .Z(n26315) );
  XOR U26269 ( .A(n26327), .B(n26328), .Z(n26285) );
  XOR U26270 ( .A(n26329), .B(n26330), .Z(n26328) );
  XOR U26271 ( .A(n25101), .B(n26290), .Z(n26330) );
  XNOR U26272 ( .A(n26331), .B(n26332), .Z(n26290) );
  XOR U26273 ( .A(n24600), .B(n25106), .Z(n26332) );
  XOR U26274 ( .A(n25113), .B(n26333), .Z(n26331) );
  XNOR U26275 ( .A(key[185]), .B(n24653), .Z(n26333) );
  XOR U26276 ( .A(n25103), .B(n26334), .Z(n26327) );
  XNOR U26277 ( .A(key[187]), .B(n24604), .Z(n26334) );
  XOR U26278 ( .A(n26309), .B(n25070), .Z(n25103) );
  XNOR U26279 ( .A(n26335), .B(n26336), .Z(n25787) );
  XOR U26280 ( .A(n25107), .B(n26337), .Z(n26335) );
  XOR U26281 ( .A(key[184]), .B(n26320), .Z(n26337) );
  IV U26282 ( .A(n23411), .Z(n21693) );
  XOR U26283 ( .A(n25722), .B(n25776), .Z(n23411) );
  XNOR U26284 ( .A(n25834), .B(n26338), .Z(n25776) );
  XOR U26285 ( .A(n26339), .B(n25755), .Z(n26338) );
  OR U26286 ( .A(n26340), .B(n25847), .Z(n25755) );
  XNOR U26287 ( .A(n25758), .B(n25843), .Z(n25847) );
  ANDN U26288 ( .B(n25843), .A(n26341), .Z(n26339) );
  IV U26289 ( .A(n25775), .Z(n25722) );
  XNOR U26290 ( .A(n26343), .B(n25836), .Z(n26342) );
  XOR U26291 ( .A(n26345), .B(n25726), .Z(n25830) );
  ANDN U26292 ( .B(n26346), .A(n25833), .Z(n26343) );
  IV U26293 ( .A(n26345), .Z(n25833) );
  XNOR U26294 ( .A(n25834), .B(n26347), .Z(n25753) );
  XNOR U26295 ( .A(n26348), .B(n26349), .Z(n26347) );
  NANDN U26296 ( .A(n25852), .B(n26350), .Z(n26349) );
  XOR U26297 ( .A(n26351), .B(n26348), .Z(n25834) );
  OR U26298 ( .A(n25855), .B(n26352), .Z(n26348) );
  XNOR U26299 ( .A(n25858), .B(n25852), .Z(n25855) );
  XNOR U26300 ( .A(n25843), .B(n25726), .Z(n25852) );
  XOR U26301 ( .A(n26353), .B(n26354), .Z(n25726) );
  NANDN U26302 ( .A(n26355), .B(n26356), .Z(n26354) );
  XOR U26303 ( .A(n26357), .B(n26358), .Z(n25843) );
  NANDN U26304 ( .A(n26355), .B(n26359), .Z(n26358) );
  NOR U26305 ( .A(n25858), .B(n26360), .Z(n26351) );
  XNOR U26306 ( .A(n26345), .B(n25758), .Z(n25858) );
  XNOR U26307 ( .A(n26361), .B(n26357), .Z(n25758) );
  NANDN U26308 ( .A(n26362), .B(n26363), .Z(n26357) );
  XOR U26309 ( .A(n26359), .B(n26364), .Z(n26363) );
  ANDN U26310 ( .B(n26364), .A(n26365), .Z(n26361) );
  XNOR U26311 ( .A(n26366), .B(n26353), .Z(n26345) );
  NANDN U26312 ( .A(n26362), .B(n26367), .Z(n26353) );
  XOR U26313 ( .A(n26368), .B(n26356), .Z(n26367) );
  XNOR U26314 ( .A(n26369), .B(n26370), .Z(n26355) );
  XOR U26315 ( .A(n26371), .B(n26372), .Z(n26370) );
  XNOR U26316 ( .A(n26373), .B(n26374), .Z(n26369) );
  XNOR U26317 ( .A(n26375), .B(n26376), .Z(n26374) );
  ANDN U26318 ( .B(n26368), .A(n26372), .Z(n26375) );
  ANDN U26319 ( .B(n26368), .A(n26365), .Z(n26366) );
  XNOR U26320 ( .A(n26371), .B(n26377), .Z(n26365) );
  XOR U26321 ( .A(n26378), .B(n26376), .Z(n26377) );
  NAND U26322 ( .A(n26379), .B(n26380), .Z(n26376) );
  XNOR U26323 ( .A(n26373), .B(n26356), .Z(n26380) );
  IV U26324 ( .A(n26368), .Z(n26373) );
  XNOR U26325 ( .A(n26359), .B(n26372), .Z(n26379) );
  IV U26326 ( .A(n26364), .Z(n26372) );
  XOR U26327 ( .A(n26381), .B(n26382), .Z(n26364) );
  XNOR U26328 ( .A(n26383), .B(n26384), .Z(n26382) );
  XNOR U26329 ( .A(n26385), .B(n26386), .Z(n26381) );
  ANDN U26330 ( .B(n26346), .A(n26387), .Z(n26385) );
  AND U26331 ( .A(n26356), .B(n26359), .Z(n26378) );
  XNOR U26332 ( .A(n26356), .B(n26359), .Z(n26371) );
  XNOR U26333 ( .A(n26388), .B(n26389), .Z(n26359) );
  XNOR U26334 ( .A(n26390), .B(n26384), .Z(n26389) );
  XOR U26335 ( .A(n26391), .B(n26392), .Z(n26388) );
  XNOR U26336 ( .A(n26393), .B(n26386), .Z(n26392) );
  OR U26337 ( .A(n25831), .B(n26344), .Z(n26386) );
  XNOR U26338 ( .A(n26346), .B(n26394), .Z(n26344) );
  XNOR U26339 ( .A(n26387), .B(n25727), .Z(n25831) );
  ANDN U26340 ( .B(n26395), .A(n25838), .Z(n26393) );
  XNOR U26341 ( .A(n26396), .B(n26397), .Z(n26356) );
  XNOR U26342 ( .A(n26384), .B(n26398), .Z(n26397) );
  XOR U26343 ( .A(n25846), .B(n26391), .Z(n26398) );
  XNOR U26344 ( .A(n26346), .B(n26387), .Z(n26384) );
  XOR U26345 ( .A(n25757), .B(n26399), .Z(n26396) );
  XNOR U26346 ( .A(n26400), .B(n26401), .Z(n26399) );
  ANDN U26347 ( .B(n26402), .A(n26341), .Z(n26400) );
  XNOR U26348 ( .A(n26403), .B(n26404), .Z(n26368) );
  XNOR U26349 ( .A(n26390), .B(n26405), .Z(n26404) );
  XNOR U26350 ( .A(n25842), .B(n26383), .Z(n26405) );
  XOR U26351 ( .A(n26391), .B(n26406), .Z(n26383) );
  XNOR U26352 ( .A(n26407), .B(n26408), .Z(n26406) );
  NAND U26353 ( .A(n26350), .B(n25853), .Z(n26408) );
  XNOR U26354 ( .A(n26409), .B(n26407), .Z(n26391) );
  NANDN U26355 ( .A(n26352), .B(n25856), .Z(n26407) );
  XOR U26356 ( .A(n25857), .B(n25853), .Z(n25856) );
  XNOR U26357 ( .A(n26402), .B(n25727), .Z(n25853) );
  XOR U26358 ( .A(n26360), .B(n26350), .Z(n26352) );
  XNOR U26359 ( .A(n26341), .B(n26394), .Z(n26350) );
  ANDN U26360 ( .B(n25857), .A(n26360), .Z(n26409) );
  XOR U26361 ( .A(n25757), .B(n26346), .Z(n26360) );
  XNOR U26362 ( .A(n26410), .B(n26411), .Z(n26346) );
  XNOR U26363 ( .A(n26412), .B(n26413), .Z(n26411) );
  XOR U26364 ( .A(n26394), .B(n26395), .Z(n26390) );
  IV U26365 ( .A(n25727), .Z(n26395) );
  XOR U26366 ( .A(n26414), .B(n26415), .Z(n25727) );
  XOR U26367 ( .A(n26416), .B(n26413), .Z(n26415) );
  IV U26368 ( .A(n25838), .Z(n26394) );
  XOR U26369 ( .A(n26413), .B(n26417), .Z(n25838) );
  XNOR U26370 ( .A(n26418), .B(n26419), .Z(n26403) );
  XNOR U26371 ( .A(n26420), .B(n26401), .Z(n26419) );
  OR U26372 ( .A(n25848), .B(n26340), .Z(n26401) );
  XNOR U26373 ( .A(n25757), .B(n26341), .Z(n26340) );
  IV U26374 ( .A(n26418), .Z(n26341) );
  XOR U26375 ( .A(n25846), .B(n26402), .Z(n25848) );
  IV U26376 ( .A(n25842), .Z(n26402) );
  XOR U26377 ( .A(n25832), .B(n26421), .Z(n25842) );
  XNOR U26378 ( .A(n26422), .B(n26410), .Z(n26421) );
  XOR U26379 ( .A(n26423), .B(n26424), .Z(n26410) );
  XNOR U26380 ( .A(n24498), .B(n26425), .Z(n26424) );
  IV U26381 ( .A(n25565), .Z(n24498) );
  XOR U26382 ( .A(n26426), .B(n25569), .Z(n25565) );
  XOR U26383 ( .A(key[146]), .B(n24504), .Z(n26423) );
  IV U26384 ( .A(n26387), .Z(n25832) );
  XOR U26385 ( .A(n26414), .B(n26427), .Z(n26387) );
  XOR U26386 ( .A(n26413), .B(n26428), .Z(n26427) );
  NOR U26387 ( .A(n25846), .B(n25757), .Z(n26420) );
  XOR U26388 ( .A(n26414), .B(n26429), .Z(n25846) );
  XOR U26389 ( .A(n26413), .B(n26430), .Z(n26429) );
  XOR U26390 ( .A(n26431), .B(n26432), .Z(n26413) );
  XNOR U26391 ( .A(n25757), .B(n26433), .Z(n26432) );
  XNOR U26392 ( .A(n25542), .B(n26434), .Z(n26431) );
  XNOR U26393 ( .A(key[150]), .B(n26435), .Z(n26434) );
  XNOR U26394 ( .A(n26436), .B(n25531), .Z(n25542) );
  IV U26395 ( .A(n26417), .Z(n26414) );
  XOR U26396 ( .A(n26437), .B(n26438), .Z(n26417) );
  XOR U26397 ( .A(n26439), .B(n26440), .Z(n26438) );
  XNOR U26398 ( .A(key[149]), .B(n25552), .Z(n26437) );
  XNOR U26399 ( .A(n25538), .B(n26435), .Z(n25552) );
  XOR U26400 ( .A(n26441), .B(n26442), .Z(n26418) );
  XNOR U26401 ( .A(n26430), .B(n26428), .Z(n26442) );
  XNOR U26402 ( .A(n26443), .B(n26444), .Z(n26428) );
  XOR U26403 ( .A(n26445), .B(n26446), .Z(n26444) );
  XOR U26404 ( .A(key[151]), .B(n26436), .Z(n26443) );
  XNOR U26405 ( .A(n26447), .B(n26448), .Z(n26430) );
  XNOR U26406 ( .A(n25515), .B(n26449), .Z(n26448) );
  XNOR U26407 ( .A(n25547), .B(n25536), .Z(n25515) );
  XOR U26408 ( .A(key[148]), .B(n25516), .Z(n26447) );
  XNOR U26409 ( .A(n25757), .B(n26412), .Z(n26441) );
  XOR U26410 ( .A(n26450), .B(n26451), .Z(n26412) );
  XNOR U26411 ( .A(n26452), .B(n26453), .Z(n26451) );
  XNOR U26412 ( .A(n25557), .B(n26422), .Z(n26453) );
  IV U26413 ( .A(n26416), .Z(n26422) );
  XNOR U26414 ( .A(n26454), .B(n26455), .Z(n26416) );
  XNOR U26415 ( .A(n26456), .B(n24465), .Z(n26455) );
  XOR U26416 ( .A(n25562), .B(n26425), .Z(n24465) );
  XNOR U26417 ( .A(key[145]), .B(n24511), .Z(n26454) );
  XNOR U26418 ( .A(n25547), .B(n25517), .Z(n25557) );
  IV U26419 ( .A(n26436), .Z(n25547) );
  XOR U26420 ( .A(n26457), .B(n26458), .Z(n26450) );
  XNOR U26421 ( .A(key[147]), .B(n26426), .Z(n26458) );
  XNOR U26422 ( .A(n26459), .B(n26460), .Z(n25757) );
  XNOR U26423 ( .A(n24503), .B(n25546), .Z(n26460) );
  XNOR U26424 ( .A(n26461), .B(n26462), .Z(n24503) );
  XNOR U26425 ( .A(key[144]), .B(n25520), .Z(n26459) );
  IV U26426 ( .A(n25553), .Z(n25520) );
  XOR U26427 ( .A(n23656), .B(n23575), .Z(n19414) );
  XNOR U26428 ( .A(n23685), .B(n26463), .Z(n23575) );
  XNOR U26429 ( .A(n26464), .B(n23597), .Z(n26463) );
  ANDN U26430 ( .B(n23694), .A(n26465), .Z(n23597) );
  XOR U26431 ( .A(n26466), .B(n23599), .Z(n23694) );
  ANDN U26432 ( .B(n26467), .A(n23669), .Z(n26464) );
  IV U26433 ( .A(n26466), .Z(n23669) );
  XNOR U26434 ( .A(n23595), .B(n26468), .Z(n23685) );
  XNOR U26435 ( .A(n26469), .B(n26470), .Z(n26468) );
  NANDN U26436 ( .A(n23674), .B(n26471), .Z(n26470) );
  XOR U26437 ( .A(n23569), .B(n23574), .Z(n23656) );
  XNOR U26438 ( .A(n23595), .B(n26472), .Z(n23574) );
  XNOR U26439 ( .A(n23687), .B(n26473), .Z(n26472) );
  NANDN U26440 ( .A(n26474), .B(n26475), .Z(n26473) );
  OR U26441 ( .A(n26476), .B(n26477), .Z(n23687) );
  XOR U26442 ( .A(n26478), .B(n26469), .Z(n23595) );
  NANDN U26443 ( .A(n26479), .B(n26480), .Z(n26469) );
  ANDN U26444 ( .B(n26481), .A(n26482), .Z(n26478) );
  XOR U26445 ( .A(n23670), .B(n26483), .Z(n23569) );
  XOR U26446 ( .A(n26484), .B(n23659), .Z(n26483) );
  OR U26447 ( .A(n26485), .B(n26476), .Z(n23659) );
  XNOR U26448 ( .A(n23662), .B(n26475), .Z(n26476) );
  ANDN U26449 ( .B(n26475), .A(n26486), .Z(n26484) );
  XOR U26450 ( .A(n26487), .B(n23672), .Z(n23670) );
  OR U26451 ( .A(n26479), .B(n26488), .Z(n23672) );
  XNOR U26452 ( .A(n26482), .B(n23674), .Z(n26479) );
  XNOR U26453 ( .A(n26475), .B(n23599), .Z(n23674) );
  XOR U26454 ( .A(n26489), .B(n26490), .Z(n23599) );
  NANDN U26455 ( .A(n26491), .B(n26492), .Z(n26490) );
  XOR U26456 ( .A(n26493), .B(n26494), .Z(n26475) );
  NANDN U26457 ( .A(n26491), .B(n26495), .Z(n26494) );
  NOR U26458 ( .A(n26482), .B(n26496), .Z(n26487) );
  XNOR U26459 ( .A(n26466), .B(n23662), .Z(n26482) );
  XNOR U26460 ( .A(n26497), .B(n26493), .Z(n23662) );
  NANDN U26461 ( .A(n26498), .B(n26499), .Z(n26493) );
  XOR U26462 ( .A(n26495), .B(n26500), .Z(n26499) );
  ANDN U26463 ( .B(n26500), .A(n26501), .Z(n26497) );
  XNOR U26464 ( .A(n26502), .B(n26489), .Z(n26466) );
  NANDN U26465 ( .A(n26498), .B(n26503), .Z(n26489) );
  XOR U26466 ( .A(n26504), .B(n26492), .Z(n26503) );
  XNOR U26467 ( .A(n26505), .B(n26506), .Z(n26491) );
  XOR U26468 ( .A(n26507), .B(n26508), .Z(n26506) );
  XNOR U26469 ( .A(n26509), .B(n26510), .Z(n26505) );
  XNOR U26470 ( .A(n26511), .B(n26512), .Z(n26510) );
  ANDN U26471 ( .B(n26504), .A(n26508), .Z(n26511) );
  ANDN U26472 ( .B(n26504), .A(n26501), .Z(n26502) );
  XNOR U26473 ( .A(n26507), .B(n26513), .Z(n26501) );
  XOR U26474 ( .A(n26514), .B(n26512), .Z(n26513) );
  NAND U26475 ( .A(n26515), .B(n26516), .Z(n26512) );
  XNOR U26476 ( .A(n26509), .B(n26492), .Z(n26516) );
  IV U26477 ( .A(n26504), .Z(n26509) );
  XNOR U26478 ( .A(n26495), .B(n26508), .Z(n26515) );
  IV U26479 ( .A(n26500), .Z(n26508) );
  XOR U26480 ( .A(n26517), .B(n26518), .Z(n26500) );
  XNOR U26481 ( .A(n26519), .B(n26520), .Z(n26518) );
  XNOR U26482 ( .A(n26521), .B(n26522), .Z(n26517) );
  ANDN U26483 ( .B(n23668), .A(n26523), .Z(n26521) );
  AND U26484 ( .A(n26492), .B(n26495), .Z(n26514) );
  XNOR U26485 ( .A(n26492), .B(n26495), .Z(n26507) );
  XNOR U26486 ( .A(n26524), .B(n26525), .Z(n26495) );
  XNOR U26487 ( .A(n26526), .B(n26520), .Z(n26525) );
  XOR U26488 ( .A(n26527), .B(n26528), .Z(n26524) );
  XNOR U26489 ( .A(n26529), .B(n26522), .Z(n26528) );
  OR U26490 ( .A(n26465), .B(n23693), .Z(n26522) );
  XNOR U26491 ( .A(n23668), .B(n26530), .Z(n23693) );
  XNOR U26492 ( .A(n26523), .B(n23600), .Z(n26465) );
  ANDN U26493 ( .B(n26531), .A(n23692), .Z(n26529) );
  XNOR U26494 ( .A(n26532), .B(n26533), .Z(n26492) );
  XNOR U26495 ( .A(n26520), .B(n26534), .Z(n26533) );
  XOR U26496 ( .A(n23689), .B(n26527), .Z(n26534) );
  XNOR U26497 ( .A(n23668), .B(n26523), .Z(n26520) );
  XOR U26498 ( .A(n23661), .B(n26535), .Z(n26532) );
  XNOR U26499 ( .A(n26536), .B(n26537), .Z(n26535) );
  ANDN U26500 ( .B(n26538), .A(n26486), .Z(n26536) );
  XNOR U26501 ( .A(n26539), .B(n26540), .Z(n26504) );
  XNOR U26502 ( .A(n26526), .B(n26541), .Z(n26540) );
  XNOR U26503 ( .A(n26474), .B(n26519), .Z(n26541) );
  XOR U26504 ( .A(n26527), .B(n26542), .Z(n26519) );
  XNOR U26505 ( .A(n26543), .B(n26544), .Z(n26542) );
  NAND U26506 ( .A(n23675), .B(n26471), .Z(n26544) );
  XNOR U26507 ( .A(n26545), .B(n26543), .Z(n26527) );
  NANDN U26508 ( .A(n26488), .B(n26480), .Z(n26543) );
  XOR U26509 ( .A(n26481), .B(n26471), .Z(n26480) );
  XNOR U26510 ( .A(n26538), .B(n23600), .Z(n26471) );
  XOR U26511 ( .A(n26496), .B(n23675), .Z(n26488) );
  XNOR U26512 ( .A(n26486), .B(n26530), .Z(n23675) );
  ANDN U26513 ( .B(n26481), .A(n26496), .Z(n26545) );
  XOR U26514 ( .A(n23661), .B(n23668), .Z(n26496) );
  XNOR U26515 ( .A(n26546), .B(n26547), .Z(n23668) );
  XNOR U26516 ( .A(n26548), .B(n26549), .Z(n26547) );
  XOR U26517 ( .A(n26530), .B(n26531), .Z(n26526) );
  IV U26518 ( .A(n23600), .Z(n26531) );
  XOR U26519 ( .A(n26550), .B(n26551), .Z(n23600) );
  XNOR U26520 ( .A(n26552), .B(n26549), .Z(n26551) );
  IV U26521 ( .A(n23692), .Z(n26530) );
  XOR U26522 ( .A(n26549), .B(n26553), .Z(n23692) );
  XNOR U26523 ( .A(n26554), .B(n26555), .Z(n26539) );
  XNOR U26524 ( .A(n26556), .B(n26537), .Z(n26555) );
  OR U26525 ( .A(n26477), .B(n26485), .Z(n26537) );
  XNOR U26526 ( .A(n23661), .B(n26486), .Z(n26485) );
  IV U26527 ( .A(n26554), .Z(n26486) );
  XOR U26528 ( .A(n23689), .B(n26538), .Z(n26477) );
  IV U26529 ( .A(n26474), .Z(n26538) );
  XOR U26530 ( .A(n26467), .B(n26557), .Z(n26474) );
  XNOR U26531 ( .A(n26552), .B(n26546), .Z(n26557) );
  XOR U26532 ( .A(n26558), .B(n26559), .Z(n26546) );
  XNOR U26533 ( .A(n26560), .B(n21194), .Z(n21233) );
  XOR U26534 ( .A(n22235), .B(n26561), .Z(n26558) );
  XNOR U26535 ( .A(key[330]), .B(n23038), .Z(n26561) );
  XNOR U26536 ( .A(n26562), .B(n26563), .Z(n22235) );
  XNOR U26537 ( .A(n26564), .B(n26565), .Z(n26563) );
  IV U26538 ( .A(n26523), .Z(n26467) );
  XOR U26539 ( .A(n26550), .B(n26566), .Z(n26523) );
  XOR U26540 ( .A(n26549), .B(n26567), .Z(n26566) );
  NOR U26541 ( .A(n23689), .B(n23661), .Z(n26556) );
  XOR U26542 ( .A(n26550), .B(n26568), .Z(n23689) );
  XOR U26543 ( .A(n26549), .B(n26569), .Z(n26568) );
  XOR U26544 ( .A(n26570), .B(n26571), .Z(n26549) );
  XNOR U26545 ( .A(n22212), .B(n21204), .Z(n26571) );
  XOR U26546 ( .A(n21218), .B(n23008), .Z(n21204) );
  XNOR U26547 ( .A(n21211), .B(n22222), .Z(n22212) );
  XOR U26548 ( .A(n21242), .B(n23009), .Z(n22222) );
  XOR U26549 ( .A(n26562), .B(n26572), .Z(n23009) );
  XNOR U26550 ( .A(n26573), .B(n26574), .Z(n26572) );
  XNOR U26551 ( .A(n26575), .B(n26576), .Z(n26562) );
  XNOR U26552 ( .A(n23025), .B(n21206), .Z(n21211) );
  XNOR U26553 ( .A(n26577), .B(n26578), .Z(n21206) );
  XNOR U26554 ( .A(n23015), .B(n26579), .Z(n26570) );
  XOR U26555 ( .A(key[334]), .B(n23661), .Z(n26579) );
  XNOR U26556 ( .A(n26580), .B(n26581), .Z(n23015) );
  IV U26557 ( .A(n26553), .Z(n26550) );
  XOR U26558 ( .A(n26582), .B(n26583), .Z(n26553) );
  XOR U26559 ( .A(n22996), .B(n22215), .Z(n26583) );
  XNOR U26560 ( .A(n23013), .B(n21209), .Z(n22215) );
  XNOR U26561 ( .A(n26584), .B(n26585), .Z(n21209) );
  XNOR U26562 ( .A(n26586), .B(n26587), .Z(n26585) );
  XNOR U26563 ( .A(n26588), .B(n26589), .Z(n26584) );
  XOR U26564 ( .A(n26590), .B(n26591), .Z(n26589) );
  ANDN U26565 ( .B(n26592), .A(n26593), .Z(n26591) );
  XNOR U26566 ( .A(n26594), .B(n26595), .Z(n22996) );
  XNOR U26567 ( .A(n26596), .B(n26597), .Z(n26595) );
  XNOR U26568 ( .A(n26598), .B(n26599), .Z(n26594) );
  XNOR U26569 ( .A(n26600), .B(n26601), .Z(n26599) );
  ANDN U26570 ( .B(n26602), .A(n26603), .Z(n26601) );
  XNOR U26571 ( .A(n22210), .B(n26604), .Z(n26582) );
  XNOR U26572 ( .A(key[333]), .B(n23025), .Z(n26604) );
  XOR U26573 ( .A(n26605), .B(n26606), .Z(n23025) );
  XNOR U26574 ( .A(n26565), .B(n26573), .Z(n22210) );
  XNOR U26575 ( .A(n26609), .B(n26610), .Z(n26565) );
  XNOR U26576 ( .A(n26611), .B(n26612), .Z(n26610) );
  NOR U26577 ( .A(n26613), .B(n26614), .Z(n26611) );
  XOR U26578 ( .A(n26615), .B(n26616), .Z(n26554) );
  XNOR U26579 ( .A(n26569), .B(n26567), .Z(n26616) );
  XNOR U26580 ( .A(n26617), .B(n26618), .Z(n26567) );
  XOR U26581 ( .A(n23010), .B(n22223), .Z(n26618) );
  XNOR U26582 ( .A(n23008), .B(n23026), .Z(n22223) );
  XNOR U26583 ( .A(n26619), .B(n26620), .Z(n23026) );
  XOR U26584 ( .A(n26621), .B(n26587), .Z(n26620) );
  XNOR U26585 ( .A(n26622), .B(n26623), .Z(n26587) );
  XNOR U26586 ( .A(n26624), .B(n26625), .Z(n26623) );
  NANDN U26587 ( .A(n26626), .B(n26627), .Z(n26625) );
  XNOR U26588 ( .A(n26628), .B(n26629), .Z(n26619) );
  XNOR U26589 ( .A(n26630), .B(n26631), .Z(n23008) );
  XOR U26590 ( .A(n26632), .B(n26633), .Z(n26631) );
  XNOR U26591 ( .A(n26634), .B(n26635), .Z(n26630) );
  XNOR U26592 ( .A(n26636), .B(n26637), .Z(n23010) );
  XNOR U26593 ( .A(n26581), .B(n26597), .Z(n26637) );
  XNOR U26594 ( .A(n26638), .B(n26639), .Z(n26597) );
  XNOR U26595 ( .A(n26640), .B(n26641), .Z(n26639) );
  OR U26596 ( .A(n26642), .B(n26643), .Z(n26641) );
  XNOR U26597 ( .A(n26644), .B(n26645), .Z(n26636) );
  XOR U26598 ( .A(key[335]), .B(n22245), .Z(n26617) );
  XOR U26599 ( .A(n26646), .B(n21242), .Z(n22245) );
  XNOR U26600 ( .A(n26647), .B(n26648), .Z(n26569) );
  XNOR U26601 ( .A(n22227), .B(n21223), .Z(n26648) );
  XOR U26602 ( .A(n21218), .B(n23013), .Z(n21223) );
  XNOR U26603 ( .A(n26649), .B(n26650), .Z(n23013) );
  XNOR U26604 ( .A(n26651), .B(n26633), .Z(n26650) );
  XNOR U26605 ( .A(n26652), .B(n26653), .Z(n26633) );
  XNOR U26606 ( .A(n26654), .B(n26655), .Z(n26653) );
  OR U26607 ( .A(n26656), .B(n26657), .Z(n26655) );
  XNOR U26608 ( .A(n26658), .B(n26659), .Z(n26649) );
  XNOR U26609 ( .A(n26660), .B(n26661), .Z(n26659) );
  ANDN U26610 ( .B(n26662), .A(n26663), .Z(n26660) );
  XNOR U26611 ( .A(n22999), .B(n21225), .Z(n22227) );
  XNOR U26612 ( .A(n26588), .B(n23034), .Z(n21225) );
  IV U26613 ( .A(n21194), .Z(n23034) );
  XNOR U26614 ( .A(n26664), .B(n26628), .Z(n21194) );
  XNOR U26615 ( .A(n22997), .B(n26665), .Z(n26647) );
  XNOR U26616 ( .A(key[332]), .B(n22229), .Z(n26665) );
  XOR U26617 ( .A(n21242), .B(n22217), .Z(n22229) );
  XOR U26618 ( .A(n26666), .B(n26667), .Z(n22217) );
  XOR U26619 ( .A(n26668), .B(n26574), .Z(n26667) );
  XNOR U26620 ( .A(n26669), .B(n26670), .Z(n26574) );
  XNOR U26621 ( .A(n26671), .B(n26672), .Z(n26670) );
  OR U26622 ( .A(n26673), .B(n26674), .Z(n26672) );
  XNOR U26623 ( .A(n26675), .B(n26676), .Z(n26666) );
  XOR U26624 ( .A(n26612), .B(n26677), .Z(n26676) );
  ANDN U26625 ( .B(n26678), .A(n26679), .Z(n26677) );
  NOR U26626 ( .A(n26680), .B(n26681), .Z(n26612) );
  XOR U26627 ( .A(n26598), .B(n23032), .Z(n22997) );
  XOR U26628 ( .A(n26682), .B(n26645), .Z(n23032) );
  XNOR U26629 ( .A(n23661), .B(n26548), .Z(n26615) );
  XOR U26630 ( .A(n26683), .B(n26684), .Z(n26548) );
  XNOR U26631 ( .A(n21236), .B(n26685), .Z(n26684) );
  XNOR U26632 ( .A(n26552), .B(n22240), .Z(n26685) );
  XOR U26633 ( .A(n21242), .B(n22231), .Z(n22240) );
  XOR U26634 ( .A(n22202), .B(n26668), .Z(n22231) );
  XOR U26635 ( .A(n26686), .B(n26668), .Z(n21242) );
  XOR U26636 ( .A(n26669), .B(n26687), .Z(n26668) );
  XNOR U26637 ( .A(n26688), .B(n26689), .Z(n26687) );
  OR U26638 ( .A(n26614), .B(n26690), .Z(n26689) );
  XNOR U26639 ( .A(n26691), .B(n26692), .Z(n26669) );
  XNOR U26640 ( .A(n26693), .B(n26694), .Z(n26692) );
  NAND U26641 ( .A(n26695), .B(n26696), .Z(n26694) );
  XOR U26642 ( .A(n26697), .B(n26698), .Z(n26552) );
  XOR U26643 ( .A(n23036), .B(n21235), .Z(n21241) );
  IV U26644 ( .A(n23021), .Z(n21235) );
  XOR U26645 ( .A(n26621), .B(n26699), .Z(n23021) );
  XOR U26646 ( .A(n26628), .B(n26629), .Z(n26699) );
  IV U26647 ( .A(n26700), .Z(n26629) );
  IV U26648 ( .A(n26578), .Z(n26621) );
  XOR U26649 ( .A(n26664), .B(n26701), .Z(n26578) );
  XOR U26650 ( .A(n26575), .B(n26686), .Z(n22202) );
  IV U26651 ( .A(n26702), .Z(n26686) );
  XOR U26652 ( .A(n23033), .B(n26703), .Z(n26697) );
  XOR U26653 ( .A(key[329]), .B(n26560), .Z(n26703) );
  IV U26654 ( .A(n23022), .Z(n23033) );
  XOR U26655 ( .A(n26644), .B(n26645), .Z(n26704) );
  XNOR U26656 ( .A(n26682), .B(n26705), .Z(n26581) );
  XNOR U26657 ( .A(n21218), .B(n22999), .Z(n21236) );
  XOR U26658 ( .A(n26658), .B(n26560), .Z(n22999) );
  IV U26659 ( .A(n23042), .Z(n26560) );
  XOR U26660 ( .A(n26607), .B(n26635), .Z(n23042) );
  IV U26661 ( .A(n26646), .Z(n21218) );
  XNOR U26662 ( .A(n23039), .B(n26706), .Z(n26683) );
  XOR U26663 ( .A(key[331]), .B(n22242), .Z(n26706) );
  XOR U26664 ( .A(n21238), .B(n23038), .Z(n22242) );
  XOR U26665 ( .A(n26707), .B(n26708), .Z(n23038) );
  XOR U26666 ( .A(n26709), .B(n26605), .Z(n26708) );
  XOR U26667 ( .A(n26710), .B(n26711), .Z(n26605) );
  XNOR U26668 ( .A(n26661), .B(n26712), .Z(n26711) );
  OR U26669 ( .A(n26713), .B(n26714), .Z(n26712) );
  NANDN U26670 ( .A(n26715), .B(n26716), .Z(n26661) );
  XNOR U26671 ( .A(n26608), .B(n26635), .Z(n26707) );
  XOR U26672 ( .A(n26717), .B(n26718), .Z(n21238) );
  XNOR U26673 ( .A(n26628), .B(n26700), .Z(n26718) );
  XOR U26674 ( .A(n26719), .B(n26720), .Z(n26700) );
  XNOR U26675 ( .A(n26721), .B(n26722), .Z(n26720) );
  NANDN U26676 ( .A(n26723), .B(n26627), .Z(n26722) );
  XOR U26677 ( .A(n26724), .B(n26725), .Z(n26628) );
  XOR U26678 ( .A(n26726), .B(n26727), .Z(n26725) );
  NANDN U26679 ( .A(n26728), .B(n26592), .Z(n26727) );
  XNOR U26680 ( .A(n26701), .B(n26577), .Z(n26717) );
  XNOR U26681 ( .A(n26719), .B(n26729), .Z(n26577) );
  XNOR U26682 ( .A(n26730), .B(n26590), .Z(n26729) );
  ANDN U26683 ( .B(n26731), .A(n26732), .Z(n26590) );
  ANDN U26684 ( .B(n26733), .A(n26734), .Z(n26730) );
  XNOR U26685 ( .A(n26586), .B(n26735), .Z(n26719) );
  XNOR U26686 ( .A(n26736), .B(n26737), .Z(n26735) );
  NANDN U26687 ( .A(n26738), .B(n26739), .Z(n26737) );
  XOR U26688 ( .A(n26586), .B(n26740), .Z(n26701) );
  XNOR U26689 ( .A(n26721), .B(n26741), .Z(n26740) );
  NANDN U26690 ( .A(n26742), .B(n26743), .Z(n26741) );
  OR U26691 ( .A(n26744), .B(n26745), .Z(n26721) );
  XOR U26692 ( .A(n26746), .B(n26736), .Z(n26586) );
  NANDN U26693 ( .A(n26747), .B(n26748), .Z(n26736) );
  ANDN U26694 ( .B(n26749), .A(n26750), .Z(n26746) );
  XOR U26695 ( .A(n26751), .B(n26752), .Z(n23039) );
  XOR U26696 ( .A(n26645), .B(n26580), .Z(n26752) );
  XNOR U26697 ( .A(n26753), .B(n26754), .Z(n26580) );
  XOR U26698 ( .A(n26755), .B(n26600), .Z(n26754) );
  NANDN U26699 ( .A(n26756), .B(n26757), .Z(n26600) );
  ANDN U26700 ( .B(n26758), .A(n26759), .Z(n26755) );
  XOR U26701 ( .A(n26760), .B(n26761), .Z(n26645) );
  XNOR U26702 ( .A(n26762), .B(n26763), .Z(n26761) );
  NAND U26703 ( .A(n26764), .B(n26602), .Z(n26763) );
  XNOR U26704 ( .A(n26644), .B(n26705), .Z(n26751) );
  XOR U26705 ( .A(n26596), .B(n26765), .Z(n26705) );
  XNOR U26706 ( .A(n26766), .B(n26767), .Z(n26765) );
  NANDN U26707 ( .A(n26768), .B(n26769), .Z(n26767) );
  XNOR U26708 ( .A(n26753), .B(n26770), .Z(n26644) );
  XNOR U26709 ( .A(n26766), .B(n26771), .Z(n26770) );
  NANDN U26710 ( .A(n26642), .B(n26772), .Z(n26771) );
  OR U26711 ( .A(n26773), .B(n26774), .Z(n26766) );
  XNOR U26712 ( .A(n26596), .B(n26775), .Z(n26753) );
  XNOR U26713 ( .A(n26776), .B(n26777), .Z(n26775) );
  NANDN U26714 ( .A(n26778), .B(n26779), .Z(n26777) );
  XOR U26715 ( .A(n26780), .B(n26776), .Z(n26596) );
  NANDN U26716 ( .A(n26781), .B(n26782), .Z(n26776) );
  ANDN U26717 ( .B(n26783), .A(n26784), .Z(n26780) );
  XNOR U26718 ( .A(n26785), .B(n26786), .Z(n23661) );
  XOR U26719 ( .A(n23036), .B(n21243), .Z(n26786) );
  XOR U26720 ( .A(n22246), .B(n22224), .Z(n21243) );
  XOR U26721 ( .A(n26682), .B(n26598), .Z(n22224) );
  XNOR U26722 ( .A(n26638), .B(n26787), .Z(n26598) );
  XOR U26723 ( .A(n26788), .B(n26762), .Z(n26787) );
  NANDN U26724 ( .A(n26789), .B(n26757), .Z(n26762) );
  XOR U26725 ( .A(n26758), .B(n26602), .Z(n26757) );
  ANDN U26726 ( .B(n26758), .A(n26790), .Z(n26788) );
  XNOR U26727 ( .A(n26760), .B(n26791), .Z(n26638) );
  XNOR U26728 ( .A(n26792), .B(n26793), .Z(n26791) );
  NANDN U26729 ( .A(n26778), .B(n26794), .Z(n26793) );
  XOR U26730 ( .A(n26760), .B(n26795), .Z(n26682) );
  XOR U26731 ( .A(n26796), .B(n26640), .Z(n26795) );
  OR U26732 ( .A(n26797), .B(n26773), .Z(n26640) );
  XNOR U26733 ( .A(n26642), .B(n26768), .Z(n26773) );
  NOR U26734 ( .A(n26798), .B(n26768), .Z(n26796) );
  XOR U26735 ( .A(n26799), .B(n26792), .Z(n26760) );
  OR U26736 ( .A(n26781), .B(n26800), .Z(n26792) );
  XOR U26737 ( .A(n26801), .B(n26778), .Z(n26781) );
  XOR U26738 ( .A(n26768), .B(n26602), .Z(n26778) );
  XOR U26739 ( .A(n26802), .B(n26803), .Z(n26602) );
  NANDN U26740 ( .A(n26804), .B(n26805), .Z(n26803) );
  XNOR U26741 ( .A(n26806), .B(n26807), .Z(n26768) );
  OR U26742 ( .A(n26804), .B(n26808), .Z(n26807) );
  ANDN U26743 ( .B(n26801), .A(n26809), .Z(n26799) );
  IV U26744 ( .A(n26784), .Z(n26801) );
  XOR U26745 ( .A(n26642), .B(n26758), .Z(n26784) );
  XNOR U26746 ( .A(n26810), .B(n26802), .Z(n26758) );
  NANDN U26747 ( .A(n26811), .B(n26812), .Z(n26802) );
  ANDN U26748 ( .B(n26813), .A(n26814), .Z(n26810) );
  NANDN U26749 ( .A(n26811), .B(n26816), .Z(n26806) );
  XOR U26750 ( .A(n26817), .B(n26804), .Z(n26811) );
  XNOR U26751 ( .A(n26818), .B(n26819), .Z(n26804) );
  XOR U26752 ( .A(n26820), .B(n26813), .Z(n26819) );
  XNOR U26753 ( .A(n26821), .B(n26822), .Z(n26818) );
  XNOR U26754 ( .A(n26823), .B(n26824), .Z(n26822) );
  ANDN U26755 ( .B(n26813), .A(n26825), .Z(n26823) );
  IV U26756 ( .A(n26826), .Z(n26813) );
  ANDN U26757 ( .B(n26817), .A(n26825), .Z(n26815) );
  IV U26758 ( .A(n26821), .Z(n26825) );
  IV U26759 ( .A(n26814), .Z(n26817) );
  XNOR U26760 ( .A(n26820), .B(n26827), .Z(n26814) );
  XOR U26761 ( .A(n26828), .B(n26824), .Z(n26827) );
  NAND U26762 ( .A(n26816), .B(n26812), .Z(n26824) );
  XNOR U26763 ( .A(n26805), .B(n26826), .Z(n26812) );
  XOR U26764 ( .A(n26829), .B(n26830), .Z(n26826) );
  XOR U26765 ( .A(n26831), .B(n26832), .Z(n26830) );
  XNOR U26766 ( .A(n26769), .B(n26833), .Z(n26832) );
  XNOR U26767 ( .A(n26834), .B(n26835), .Z(n26829) );
  XNOR U26768 ( .A(n26836), .B(n26837), .Z(n26835) );
  ANDN U26769 ( .B(n26772), .A(n26643), .Z(n26836) );
  XNOR U26770 ( .A(n26821), .B(n26808), .Z(n26816) );
  XOR U26771 ( .A(n26838), .B(n26839), .Z(n26821) );
  XNOR U26772 ( .A(n26840), .B(n26833), .Z(n26839) );
  XOR U26773 ( .A(n26841), .B(n26842), .Z(n26833) );
  XNOR U26774 ( .A(n26843), .B(n26844), .Z(n26842) );
  NAND U26775 ( .A(n26794), .B(n26779), .Z(n26844) );
  XNOR U26776 ( .A(n26845), .B(n26846), .Z(n26838) );
  ANDN U26777 ( .B(n26847), .A(n26790), .Z(n26845) );
  ANDN U26778 ( .B(n26805), .A(n26808), .Z(n26828) );
  XOR U26779 ( .A(n26808), .B(n26805), .Z(n26820) );
  XNOR U26780 ( .A(n26848), .B(n26849), .Z(n26805) );
  XNOR U26781 ( .A(n26841), .B(n26850), .Z(n26849) );
  XNOR U26782 ( .A(n26840), .B(n26772), .Z(n26850) );
  XNOR U26783 ( .A(n26851), .B(n26852), .Z(n26848) );
  XNOR U26784 ( .A(n26853), .B(n26837), .Z(n26852) );
  OR U26785 ( .A(n26774), .B(n26797), .Z(n26837) );
  XNOR U26786 ( .A(n26851), .B(n26834), .Z(n26797) );
  XNOR U26787 ( .A(n26772), .B(n26769), .Z(n26774) );
  ANDN U26788 ( .B(n26769), .A(n26798), .Z(n26853) );
  XOR U26789 ( .A(n26854), .B(n26855), .Z(n26808) );
  XOR U26790 ( .A(n26841), .B(n26831), .Z(n26855) );
  XOR U26791 ( .A(n26764), .B(n26603), .Z(n26831) );
  XOR U26792 ( .A(n26856), .B(n26843), .Z(n26841) );
  NANDN U26793 ( .A(n26800), .B(n26782), .Z(n26843) );
  XOR U26794 ( .A(n26783), .B(n26779), .Z(n26782) );
  XNOR U26795 ( .A(n26847), .B(n26857), .Z(n26769) );
  XNOR U26796 ( .A(n26858), .B(n26859), .Z(n26857) );
  XOR U26797 ( .A(n26809), .B(n26794), .Z(n26800) );
  XNOR U26798 ( .A(n26798), .B(n26764), .Z(n26794) );
  IV U26799 ( .A(n26834), .Z(n26798) );
  XOR U26800 ( .A(n26860), .B(n26861), .Z(n26834) );
  XOR U26801 ( .A(n26862), .B(n26863), .Z(n26861) );
  XOR U26802 ( .A(n26851), .B(n26864), .Z(n26860) );
  ANDN U26803 ( .B(n26783), .A(n26809), .Z(n26856) );
  XNOR U26804 ( .A(n26851), .B(n26865), .Z(n26809) );
  XOR U26805 ( .A(n26847), .B(n26772), .Z(n26783) );
  XNOR U26806 ( .A(n26866), .B(n26867), .Z(n26772) );
  XOR U26807 ( .A(n26868), .B(n26863), .Z(n26867) );
  XNOR U26808 ( .A(n26869), .B(n26870), .Z(n26863) );
  XNOR U26809 ( .A(n24632), .B(n26323), .Z(n26870) );
  XOR U26810 ( .A(n26320), .B(n24618), .Z(n26323) );
  XNOR U26811 ( .A(n26871), .B(n26872), .Z(n24618) );
  XNOR U26812 ( .A(n26873), .B(n26874), .Z(n26872) );
  XNOR U26813 ( .A(n26875), .B(n26876), .Z(n26871) );
  XOR U26814 ( .A(n26877), .B(n26878), .Z(n26876) );
  ANDN U26815 ( .B(n26879), .A(n26880), .Z(n26878) );
  XNOR U26816 ( .A(n25110), .B(n25070), .Z(n24632) );
  XNOR U26817 ( .A(n26881), .B(n25113), .Z(n25070) );
  XNOR U26818 ( .A(n26882), .B(n24645), .Z(n25110) );
  IV U26819 ( .A(n26299), .Z(n24645) );
  XNOR U26820 ( .A(n24635), .B(n26883), .Z(n26869) );
  XNOR U26821 ( .A(key[180]), .B(n26324), .Z(n26883) );
  XNOR U26822 ( .A(n25095), .B(n26313), .Z(n24635) );
  IV U26823 ( .A(n26759), .Z(n26847) );
  XOR U26824 ( .A(n26840), .B(n26884), .Z(n26854) );
  XNOR U26825 ( .A(n26885), .B(n26846), .Z(n26884) );
  OR U26826 ( .A(n26756), .B(n26789), .Z(n26846) );
  XNOR U26827 ( .A(n26865), .B(n26764), .Z(n26789) );
  XNOR U26828 ( .A(n26759), .B(n26603), .Z(n26756) );
  ANDN U26829 ( .B(n26764), .A(n26603), .Z(n26885) );
  XOR U26830 ( .A(n26866), .B(n26886), .Z(n26603) );
  XOR U26831 ( .A(n26858), .B(n26887), .Z(n26886) );
  XOR U26832 ( .A(n26868), .B(n26866), .Z(n26764) );
  XNOR U26833 ( .A(n26790), .B(n26759), .Z(n26840) );
  XOR U26834 ( .A(n26866), .B(n26888), .Z(n26759) );
  XNOR U26835 ( .A(n26868), .B(n26862), .Z(n26888) );
  XOR U26836 ( .A(n26889), .B(n26890), .Z(n26862) );
  XNOR U26837 ( .A(n26891), .B(n24628), .Z(n26890) );
  XOR U26838 ( .A(n25098), .B(n26310), .Z(n24628) );
  XNOR U26839 ( .A(n26892), .B(n26893), .Z(n26310) );
  XNOR U26840 ( .A(n26894), .B(n26895), .Z(n26893) );
  XOR U26841 ( .A(n26896), .B(n26897), .Z(n26892) );
  XOR U26842 ( .A(n26898), .B(n26899), .Z(n25098) );
  XOR U26843 ( .A(n26900), .B(n26901), .Z(n26899) );
  XNOR U26844 ( .A(key[183]), .B(n26902), .Z(n26889) );
  XNOR U26845 ( .A(n26903), .B(n26904), .Z(n26866) );
  XNOR U26846 ( .A(n24619), .B(n26308), .Z(n26904) );
  XOR U26847 ( .A(n24612), .B(n24617), .Z(n26308) );
  IV U26848 ( .A(n26905), .Z(n24617) );
  XNOR U26849 ( .A(n26906), .B(n26907), .Z(n24612) );
  XOR U26850 ( .A(n25073), .B(n26326), .Z(n24619) );
  IV U26851 ( .A(n25086), .Z(n26326) );
  XOR U26852 ( .A(n26908), .B(n26909), .Z(n25086) );
  XNOR U26853 ( .A(n26910), .B(n26895), .Z(n26909) );
  XNOR U26854 ( .A(n26911), .B(n26912), .Z(n26895) );
  XNOR U26855 ( .A(n26913), .B(n26914), .Z(n26912) );
  OR U26856 ( .A(n26915), .B(n26916), .Z(n26914) );
  XNOR U26857 ( .A(n26881), .B(n26917), .Z(n26908) );
  XOR U26858 ( .A(n26918), .B(n26919), .Z(n26917) );
  ANDN U26859 ( .B(n26920), .A(n26921), .Z(n26919) );
  XOR U26860 ( .A(n26922), .B(n26923), .Z(n25073) );
  XOR U26861 ( .A(n26924), .B(n26901), .Z(n26923) );
  XNOR U26862 ( .A(n26925), .B(n26926), .Z(n26901) );
  XNOR U26863 ( .A(n26927), .B(n26928), .Z(n26926) );
  OR U26864 ( .A(n26929), .B(n26930), .Z(n26928) );
  XNOR U26865 ( .A(n26882), .B(n26931), .Z(n26922) );
  XOR U26866 ( .A(n26932), .B(n26933), .Z(n26931) );
  ANDN U26867 ( .B(n26934), .A(n26935), .Z(n26933) );
  XOR U26868 ( .A(key[181]), .B(n26313), .Z(n26903) );
  XNOR U26869 ( .A(n26936), .B(n26937), .Z(n26313) );
  XOR U26870 ( .A(n26938), .B(n26939), .Z(n26937) );
  XOR U26871 ( .A(n26940), .B(n26941), .Z(n26936) );
  XOR U26872 ( .A(n26942), .B(n26943), .Z(n26941) );
  ANDN U26873 ( .B(n26944), .A(n26945), .Z(n26943) );
  IV U26874 ( .A(n26865), .Z(n26790) );
  XNOR U26875 ( .A(n26859), .B(n26946), .Z(n26865) );
  XOR U26876 ( .A(n26864), .B(n26887), .Z(n26946) );
  IV U26877 ( .A(n26868), .Z(n26887) );
  XOR U26878 ( .A(n26947), .B(n26948), .Z(n26868) );
  XOR U26879 ( .A(n26306), .B(n26643), .Z(n26948) );
  IV U26880 ( .A(n26851), .Z(n26643) );
  XOR U26881 ( .A(n26949), .B(n26950), .Z(n26851) );
  XNOR U26882 ( .A(n24626), .B(n25106), .Z(n26950) );
  XNOR U26883 ( .A(n24654), .B(n24644), .Z(n25106) );
  XOR U26884 ( .A(n26951), .B(n26952), .Z(n24644) );
  XNOR U26885 ( .A(n26953), .B(n26906), .Z(n26952) );
  XOR U26886 ( .A(n24655), .B(n25095), .Z(n24626) );
  XOR U26887 ( .A(n26882), .B(n26954), .Z(n24655) );
  XNOR U26888 ( .A(n26925), .B(n26955), .Z(n26882) );
  XOR U26889 ( .A(n26956), .B(n26957), .Z(n26955) );
  XOR U26890 ( .A(n26960), .B(n26961), .Z(n26925) );
  XNOR U26891 ( .A(n26962), .B(n26963), .Z(n26961) );
  NANDN U26892 ( .A(n26964), .B(n26965), .Z(n26963) );
  XOR U26893 ( .A(key[176]), .B(n26309), .Z(n26949) );
  XNOR U26894 ( .A(n26911), .B(n26967), .Z(n26881) );
  XOR U26895 ( .A(n26968), .B(n26969), .Z(n26967) );
  XOR U26896 ( .A(n26972), .B(n26973), .Z(n26911) );
  XNOR U26897 ( .A(n26974), .B(n26975), .Z(n26973) );
  NANDN U26898 ( .A(n26976), .B(n26977), .Z(n26975) );
  XNOR U26899 ( .A(n26320), .B(n24627), .Z(n26306) );
  XNOR U26900 ( .A(n26978), .B(n26979), .Z(n24627) );
  XOR U26901 ( .A(n26980), .B(n26874), .Z(n26979) );
  XNOR U26902 ( .A(n26981), .B(n26982), .Z(n26874) );
  XNOR U26903 ( .A(n26983), .B(n26984), .Z(n26982) );
  OR U26904 ( .A(n26985), .B(n26986), .Z(n26984) );
  XOR U26905 ( .A(n26953), .B(n26906), .Z(n26978) );
  XOR U26906 ( .A(n26987), .B(n26988), .Z(n26906) );
  XOR U26907 ( .A(n26905), .B(n26989), .Z(n26947) );
  XOR U26908 ( .A(key[182]), .B(n24611), .Z(n26989) );
  XOR U26909 ( .A(n25088), .B(n26891), .Z(n24611) );
  XNOR U26910 ( .A(n25095), .B(n26319), .Z(n26891) );
  XNOR U26911 ( .A(n26990), .B(n26991), .Z(n26319) );
  XOR U26912 ( .A(n26992), .B(n26939), .Z(n26991) );
  XNOR U26913 ( .A(n26993), .B(n26994), .Z(n26939) );
  XNOR U26914 ( .A(n26995), .B(n26996), .Z(n26994) );
  NANDN U26915 ( .A(n26997), .B(n26998), .Z(n26996) );
  XOR U26916 ( .A(n26999), .B(n27000), .Z(n26990) );
  XNOR U26917 ( .A(n24621), .B(n25096), .Z(n25088) );
  XNOR U26918 ( .A(n26897), .B(n27001), .Z(n25096) );
  XNOR U26919 ( .A(n26900), .B(n27002), .Z(n24621) );
  XOR U26920 ( .A(n27004), .B(n27005), .Z(n26864) );
  XNOR U26921 ( .A(n26858), .B(n27006), .Z(n27005) );
  XNOR U26922 ( .A(n24601), .B(n26329), .Z(n27006) );
  XOR U26923 ( .A(n26320), .B(n24631), .Z(n26329) );
  XNOR U26924 ( .A(n26875), .B(n24600), .Z(n24631) );
  IV U26925 ( .A(n26902), .Z(n26320) );
  XOR U26926 ( .A(n26875), .B(n26987), .Z(n26902) );
  XNOR U26927 ( .A(n26981), .B(n27007), .Z(n26875) );
  XOR U26928 ( .A(n27008), .B(n27009), .Z(n27007) );
  XNOR U26929 ( .A(n27012), .B(n27013), .Z(n26981) );
  XNOR U26930 ( .A(n27014), .B(n27015), .Z(n27013) );
  NANDN U26931 ( .A(n27016), .B(n27017), .Z(n27015) );
  XOR U26932 ( .A(n27018), .B(n27019), .Z(n26858) );
  XNOR U26933 ( .A(n24643), .B(n25114), .Z(n27019) );
  XOR U26934 ( .A(n27020), .B(n24600), .Z(n25114) );
  XOR U26935 ( .A(n26987), .B(n26980), .Z(n24600) );
  XOR U26936 ( .A(n27012), .B(n27021), .Z(n26987) );
  XOR U26937 ( .A(n27022), .B(n26983), .Z(n27021) );
  OR U26938 ( .A(n27023), .B(n27024), .Z(n26983) );
  ANDN U26939 ( .B(n27025), .A(n27026), .Z(n27022) );
  XNOR U26940 ( .A(n24653), .B(n25107), .Z(n24643) );
  XNOR U26941 ( .A(n27027), .B(n27028), .Z(n25107) );
  XNOR U26942 ( .A(n26896), .B(n26897), .Z(n27028) );
  XOR U26943 ( .A(n26966), .B(n27029), .Z(n26897) );
  XOR U26944 ( .A(n26900), .B(n27030), .Z(n24653) );
  XNOR U26945 ( .A(n27031), .B(n27032), .Z(n27030) );
  XOR U26946 ( .A(n26954), .B(n27033), .Z(n26900) );
  XOR U26947 ( .A(key[177]), .B(n24654), .Z(n27018) );
  XNOR U26948 ( .A(n26992), .B(n27034), .Z(n24654) );
  XOR U26949 ( .A(n27035), .B(n27000), .Z(n27034) );
  XOR U26950 ( .A(n27036), .B(n27037), .Z(n26992) );
  XOR U26951 ( .A(n24640), .B(n27038), .Z(n27004) );
  XNOR U26952 ( .A(key[179]), .B(n24650), .Z(n27038) );
  XOR U26953 ( .A(n25095), .B(n26324), .Z(n24650) );
  XOR U26954 ( .A(n26938), .B(n24647), .Z(n26324) );
  XOR U26955 ( .A(n27036), .B(n26938), .Z(n25095) );
  XOR U26956 ( .A(n26993), .B(n27039), .Z(n26938) );
  XOR U26957 ( .A(n27040), .B(n27041), .Z(n27039) );
  ANDN U26958 ( .B(n27042), .A(n27043), .Z(n27040) );
  XOR U26959 ( .A(n27044), .B(n27045), .Z(n26993) );
  XNOR U26960 ( .A(n27046), .B(n27047), .Z(n27045) );
  NAND U26961 ( .A(n27048), .B(n27049), .Z(n27047) );
  XOR U26962 ( .A(n24604), .B(n25108), .Z(n24640) );
  XOR U26963 ( .A(n27050), .B(n27051), .Z(n25108) );
  XNOR U26964 ( .A(n26894), .B(n27001), .Z(n27051) );
  XNOR U26965 ( .A(n27052), .B(n27053), .Z(n27001) );
  XNOR U26966 ( .A(n27054), .B(n26918), .Z(n27053) );
  NOR U26967 ( .A(n27055), .B(n27056), .Z(n26918) );
  ANDN U26968 ( .B(n26971), .A(n27057), .Z(n27054) );
  XOR U26969 ( .A(n26896), .B(n27029), .Z(n27050) );
  XOR U26970 ( .A(n26910), .B(n27058), .Z(n27029) );
  XNOR U26971 ( .A(n27059), .B(n27060), .Z(n27058) );
  NANDN U26972 ( .A(n27061), .B(n27062), .Z(n27060) );
  XNOR U26973 ( .A(n27059), .B(n27064), .Z(n27063) );
  OR U26974 ( .A(n26915), .B(n27065), .Z(n27064) );
  OR U26975 ( .A(n27066), .B(n27067), .Z(n27059) );
  XNOR U26976 ( .A(n26910), .B(n27068), .Z(n27052) );
  XNOR U26977 ( .A(n27069), .B(n27070), .Z(n27068) );
  OR U26978 ( .A(n26976), .B(n27071), .Z(n27070) );
  XOR U26979 ( .A(n27072), .B(n27069), .Z(n26910) );
  NANDN U26980 ( .A(n27073), .B(n27074), .Z(n27069) );
  ANDN U26981 ( .B(n27075), .A(n27076), .Z(n27072) );
  XOR U26982 ( .A(n26898), .B(n27077), .Z(n24604) );
  XOR U26983 ( .A(n27033), .B(n27002), .Z(n27077) );
  XNOR U26984 ( .A(n27078), .B(n27079), .Z(n27002) );
  XNOR U26985 ( .A(n27080), .B(n26932), .Z(n27079) );
  NOR U26986 ( .A(n27081), .B(n27082), .Z(n26932) );
  ANDN U26987 ( .B(n26959), .A(n27083), .Z(n27080) );
  XNOR U26988 ( .A(n26924), .B(n27084), .Z(n27033) );
  XNOR U26989 ( .A(n27085), .B(n27086), .Z(n27084) );
  NANDN U26990 ( .A(n27087), .B(n27088), .Z(n27086) );
  XOR U26991 ( .A(n27031), .B(n27032), .Z(n26898) );
  XNOR U26992 ( .A(n27085), .B(n27090), .Z(n27089) );
  OR U26993 ( .A(n26929), .B(n27091), .Z(n27090) );
  OR U26994 ( .A(n27092), .B(n27093), .Z(n27085) );
  XOR U26995 ( .A(n26924), .B(n27094), .Z(n27078) );
  XNOR U26996 ( .A(n27095), .B(n27096), .Z(n27094) );
  OR U26997 ( .A(n26964), .B(n27097), .Z(n27096) );
  XNOR U26998 ( .A(n27098), .B(n27095), .Z(n26924) );
  NANDN U26999 ( .A(n27099), .B(n27100), .Z(n27095) );
  ANDN U27000 ( .B(n27101), .A(n27102), .Z(n27098) );
  XOR U27001 ( .A(n27103), .B(n27104), .Z(n26859) );
  XOR U27002 ( .A(n24602), .B(n25101), .Z(n27104) );
  XOR U27003 ( .A(n24638), .B(n24601), .Z(n25101) );
  XNOR U27004 ( .A(n27105), .B(n27106), .Z(n24601) );
  XOR U27005 ( .A(n27037), .B(n27003), .Z(n27106) );
  XNOR U27006 ( .A(n27107), .B(n27108), .Z(n27003) );
  XNOR U27007 ( .A(n27109), .B(n26942), .Z(n27108) );
  NOR U27008 ( .A(n27110), .B(n27111), .Z(n26942) );
  ANDN U27009 ( .B(n27042), .A(n27112), .Z(n27109) );
  XNOR U27010 ( .A(n26940), .B(n27113), .Z(n27037) );
  XNOR U27011 ( .A(n27114), .B(n27115), .Z(n27113) );
  OR U27012 ( .A(n27116), .B(n27117), .Z(n27115) );
  XNOR U27013 ( .A(n27035), .B(n27000), .Z(n27105) );
  XNOR U27014 ( .A(n27114), .B(n27119), .Z(n27118) );
  NANDN U27015 ( .A(n26997), .B(n27120), .Z(n27119) );
  OR U27016 ( .A(n27121), .B(n27122), .Z(n27114) );
  XOR U27017 ( .A(n26940), .B(n27123), .Z(n27107) );
  XNOR U27018 ( .A(n27124), .B(n27125), .Z(n27123) );
  NAND U27019 ( .A(n27048), .B(n27126), .Z(n27125) );
  XNOR U27020 ( .A(n27127), .B(n27124), .Z(n26940) );
  NANDN U27021 ( .A(n27128), .B(n27129), .Z(n27124) );
  ANDN U27022 ( .B(n27130), .A(n27131), .Z(n27127) );
  XOR U27023 ( .A(n27132), .B(n27133), .Z(n24638) );
  XNOR U27024 ( .A(n26951), .B(n26907), .Z(n27133) );
  XNOR U27025 ( .A(n27134), .B(n27135), .Z(n26907) );
  XNOR U27026 ( .A(n27136), .B(n26877), .Z(n27135) );
  NOR U27027 ( .A(n27137), .B(n27138), .Z(n26877) );
  ANDN U27028 ( .B(n27011), .A(n27139), .Z(n27136) );
  IV U27029 ( .A(n26980), .Z(n26951) );
  XOR U27030 ( .A(n27012), .B(n27140), .Z(n26980) );
  XNOR U27031 ( .A(n27009), .B(n27141), .Z(n27140) );
  NANDN U27032 ( .A(n27142), .B(n27143), .Z(n27141) );
  OR U27033 ( .A(n27144), .B(n27137), .Z(n27009) );
  XNOR U27034 ( .A(n27011), .B(n27143), .Z(n27137) );
  XOR U27035 ( .A(n27145), .B(n27014), .Z(n27012) );
  OR U27036 ( .A(n27146), .B(n27147), .Z(n27014) );
  ANDN U27037 ( .B(n27148), .A(n27149), .Z(n27145) );
  XOR U27038 ( .A(n26953), .B(n26988), .Z(n27132) );
  XOR U27039 ( .A(n26873), .B(n27150), .Z(n26988) );
  XNOR U27040 ( .A(n27151), .B(n27152), .Z(n27150) );
  NANDN U27041 ( .A(n27026), .B(n27153), .Z(n27152) );
  XNOR U27042 ( .A(n27151), .B(n27155), .Z(n27154) );
  OR U27043 ( .A(n26985), .B(n27156), .Z(n27155) );
  OR U27044 ( .A(n27024), .B(n27157), .Z(n27151) );
  XOR U27045 ( .A(n26985), .B(n27158), .Z(n27024) );
  XNOR U27046 ( .A(n26873), .B(n27159), .Z(n27134) );
  XNOR U27047 ( .A(n27160), .B(n27161), .Z(n27159) );
  OR U27048 ( .A(n27016), .B(n27162), .Z(n27161) );
  XOR U27049 ( .A(n27163), .B(n27160), .Z(n26873) );
  NANDN U27050 ( .A(n27146), .B(n27164), .Z(n27160) );
  XOR U27051 ( .A(n27148), .B(n27016), .Z(n27146) );
  XOR U27052 ( .A(n27158), .B(n26880), .Z(n27016) );
  IV U27053 ( .A(n27143), .Z(n26880) );
  XOR U27054 ( .A(n27165), .B(n27166), .Z(n27143) );
  NANDN U27055 ( .A(n27167), .B(n27168), .Z(n27166) );
  IV U27056 ( .A(n27026), .Z(n27158) );
  XNOR U27057 ( .A(n27169), .B(n27170), .Z(n27026) );
  NANDN U27058 ( .A(n27167), .B(n27171), .Z(n27170) );
  IV U27059 ( .A(n27172), .Z(n27148) );
  ANDN U27060 ( .B(n27173), .A(n27172), .Z(n27163) );
  XOR U27061 ( .A(n27011), .B(n26985), .Z(n27172) );
  XOR U27062 ( .A(n27174), .B(n27169), .Z(n26985) );
  NANDN U27063 ( .A(n27175), .B(n27176), .Z(n27169) );
  NANDN U27064 ( .A(n27175), .B(n27180), .Z(n27165) );
  XOR U27065 ( .A(n27181), .B(n27182), .Z(n27167) );
  XOR U27066 ( .A(n27183), .B(n27178), .Z(n27182) );
  XNOR U27067 ( .A(n27184), .B(n27185), .Z(n27181) );
  XNOR U27068 ( .A(n27186), .B(n27187), .Z(n27185) );
  ANDN U27069 ( .B(n27183), .A(n27178), .Z(n27186) );
  ANDN U27070 ( .B(n27183), .A(n27177), .Z(n27179) );
  XNOR U27071 ( .A(n27184), .B(n27188), .Z(n27177) );
  XOR U27072 ( .A(n27189), .B(n27187), .Z(n27188) );
  NAND U27073 ( .A(n27176), .B(n27180), .Z(n27187) );
  XNOR U27074 ( .A(n27171), .B(n27178), .Z(n27176) );
  XOR U27075 ( .A(n27190), .B(n27191), .Z(n27178) );
  XOR U27076 ( .A(n27192), .B(n27193), .Z(n27191) );
  XNOR U27077 ( .A(n27194), .B(n27195), .Z(n27190) );
  ANDN U27078 ( .B(n27010), .A(n27139), .Z(n27194) );
  AND U27079 ( .A(n27168), .B(n27171), .Z(n27189) );
  XNOR U27080 ( .A(n27168), .B(n27171), .Z(n27184) );
  XNOR U27081 ( .A(n27196), .B(n27197), .Z(n27171) );
  XNOR U27082 ( .A(n27198), .B(n27199), .Z(n27197) );
  XOR U27083 ( .A(n27192), .B(n27200), .Z(n27196) );
  XNOR U27084 ( .A(n27201), .B(n27195), .Z(n27200) );
  OR U27085 ( .A(n27138), .B(n27144), .Z(n27195) );
  XNOR U27086 ( .A(n27202), .B(n27142), .Z(n27144) );
  XNOR U27087 ( .A(n27139), .B(n27203), .Z(n27138) );
  NOR U27088 ( .A(n27203), .B(n27142), .Z(n27201) );
  XNOR U27089 ( .A(n27204), .B(n27205), .Z(n27168) );
  XNOR U27090 ( .A(n27206), .B(n27207), .Z(n27205) );
  XOR U27091 ( .A(n27156), .B(n27192), .Z(n27207) );
  XOR U27092 ( .A(n27010), .B(n27208), .Z(n27192) );
  XNOR U27093 ( .A(n26986), .B(n27209), .Z(n27204) );
  XNOR U27094 ( .A(n27210), .B(n27211), .Z(n27209) );
  ANDN U27095 ( .B(n27153), .A(n27212), .Z(n27210) );
  XNOR U27096 ( .A(n27213), .B(n27214), .Z(n27183) );
  XNOR U27097 ( .A(n27193), .B(n27215), .Z(n27214) );
  XNOR U27098 ( .A(n27153), .B(n27199), .Z(n27215) );
  XOR U27099 ( .A(n27142), .B(n27203), .Z(n27199) );
  XNOR U27100 ( .A(n27206), .B(n27216), .Z(n27193) );
  XNOR U27101 ( .A(n27217), .B(n27218), .Z(n27216) );
  NANDN U27102 ( .A(n27162), .B(n27017), .Z(n27218) );
  IV U27103 ( .A(n27198), .Z(n27206) );
  XNOR U27104 ( .A(n27219), .B(n27217), .Z(n27198) );
  NANDN U27105 ( .A(n27147), .B(n27164), .Z(n27217) );
  XOR U27106 ( .A(n27153), .B(n27203), .Z(n27162) );
  IV U27107 ( .A(n26879), .Z(n27203) );
  XOR U27108 ( .A(n27220), .B(n27221), .Z(n26879) );
  XNOR U27109 ( .A(n27222), .B(n27223), .Z(n27221) );
  XOR U27110 ( .A(n27149), .B(n27017), .Z(n27147) );
  XNOR U27111 ( .A(n27025), .B(n27142), .Z(n27017) );
  XNOR U27112 ( .A(n27223), .B(n27220), .Z(n27142) );
  ANDN U27113 ( .B(n27173), .A(n27149), .Z(n27219) );
  XNOR U27114 ( .A(n27224), .B(n27010), .Z(n27149) );
  IV U27115 ( .A(n27202), .Z(n27010) );
  XNOR U27116 ( .A(n27225), .B(n27226), .Z(n27202) );
  XNOR U27117 ( .A(n27227), .B(n27223), .Z(n27226) );
  XNOR U27118 ( .A(n27212), .B(n27228), .Z(n27213) );
  XNOR U27119 ( .A(n27229), .B(n27211), .Z(n27228) );
  OR U27120 ( .A(n27157), .B(n27023), .Z(n27211) );
  XOR U27121 ( .A(n26986), .B(n27025), .Z(n27023) );
  IV U27122 ( .A(n27212), .Z(n27025) );
  XOR U27123 ( .A(n27156), .B(n27153), .Z(n27157) );
  XNOR U27124 ( .A(n27208), .B(n27230), .Z(n27153) );
  XNOR U27125 ( .A(n27222), .B(n27225), .Z(n27230) );
  XNOR U27126 ( .A(msg[18]), .B(key[18]), .Z(n27225) );
  IV U27127 ( .A(n27231), .Z(n27156) );
  ANDN U27128 ( .B(n27231), .A(n26986), .Z(n27229) );
  XOR U27129 ( .A(n27232), .B(n27233), .Z(n27212) );
  XOR U27130 ( .A(n27234), .B(n27235), .Z(n27233) );
  XOR U27131 ( .A(n26986), .B(n27227), .Z(n27232) );
  XNOR U27132 ( .A(n27222), .B(n27236), .Z(n27227) );
  XNOR U27133 ( .A(msg[19]), .B(key[19]), .Z(n27236) );
  XNOR U27134 ( .A(msg[17]), .B(key[17]), .Z(n27222) );
  IV U27135 ( .A(n27224), .Z(n26986) );
  XOR U27136 ( .A(n27231), .B(n27208), .Z(n27173) );
  IV U27137 ( .A(n27139), .Z(n27208) );
  XOR U27138 ( .A(n27237), .B(n27238), .Z(n27139) );
  XOR U27139 ( .A(n27223), .B(n27235), .Z(n27238) );
  XOR U27140 ( .A(msg[23]), .B(key[23]), .Z(n27235) );
  XOR U27141 ( .A(n27220), .B(n27239), .Z(n27231) );
  XNOR U27142 ( .A(n27223), .B(n27234), .Z(n27239) );
  XNOR U27143 ( .A(msg[20]), .B(key[20]), .Z(n27234) );
  XOR U27144 ( .A(n27224), .B(n27240), .Z(n27223) );
  XNOR U27145 ( .A(msg[22]), .B(key[22]), .Z(n27240) );
  XOR U27146 ( .A(msg[16]), .B(key[16]), .Z(n27224) );
  IV U27147 ( .A(n27237), .Z(n27220) );
  XOR U27148 ( .A(msg[21]), .B(key[21]), .Z(n27237) );
  XOR U27149 ( .A(n26299), .B(n25113), .Z(n24602) );
  XOR U27150 ( .A(n26966), .B(n27027), .Z(n25113) );
  IV U27151 ( .A(n26894), .Z(n27027) );
  XOR U27152 ( .A(n26972), .B(n27241), .Z(n26894) );
  XNOR U27153 ( .A(n26969), .B(n27242), .Z(n27241) );
  NANDN U27154 ( .A(n27243), .B(n27244), .Z(n27242) );
  OR U27155 ( .A(n27245), .B(n27055), .Z(n26969) );
  XNOR U27156 ( .A(n26971), .B(n27244), .Z(n27055) );
  XOR U27157 ( .A(n27247), .B(n26913), .Z(n27246) );
  OR U27158 ( .A(n27066), .B(n27248), .Z(n26913) );
  XOR U27159 ( .A(n26915), .B(n27249), .Z(n27066) );
  ANDN U27160 ( .B(n27250), .A(n27061), .Z(n27247) );
  XNOR U27161 ( .A(n27251), .B(n26974), .Z(n26972) );
  OR U27162 ( .A(n27073), .B(n27252), .Z(n26974) );
  XOR U27163 ( .A(n27253), .B(n26976), .Z(n27073) );
  XOR U27164 ( .A(n27249), .B(n26921), .Z(n26976) );
  IV U27165 ( .A(n27244), .Z(n26921) );
  XOR U27166 ( .A(n27254), .B(n27255), .Z(n27244) );
  NANDN U27167 ( .A(n27256), .B(n27257), .Z(n27255) );
  IV U27168 ( .A(n27061), .Z(n27249) );
  XNOR U27169 ( .A(n27258), .B(n27259), .Z(n27061) );
  NANDN U27170 ( .A(n27256), .B(n27260), .Z(n27259) );
  ANDN U27171 ( .B(n27253), .A(n27261), .Z(n27251) );
  IV U27172 ( .A(n27076), .Z(n27253) );
  XOR U27173 ( .A(n26971), .B(n26915), .Z(n27076) );
  XOR U27174 ( .A(n27262), .B(n27258), .Z(n26915) );
  NANDN U27175 ( .A(n27263), .B(n27264), .Z(n27258) );
  NANDN U27176 ( .A(n27263), .B(n27268), .Z(n27254) );
  XOR U27177 ( .A(n27269), .B(n27270), .Z(n27256) );
  XOR U27178 ( .A(n27271), .B(n27266), .Z(n27270) );
  XNOR U27179 ( .A(n27272), .B(n27273), .Z(n27269) );
  XNOR U27180 ( .A(n27274), .B(n27275), .Z(n27273) );
  ANDN U27181 ( .B(n27271), .A(n27266), .Z(n27274) );
  ANDN U27182 ( .B(n27271), .A(n27265), .Z(n27267) );
  XNOR U27183 ( .A(n27272), .B(n27276), .Z(n27265) );
  XOR U27184 ( .A(n27277), .B(n27275), .Z(n27276) );
  NAND U27185 ( .A(n27264), .B(n27268), .Z(n27275) );
  XNOR U27186 ( .A(n27260), .B(n27266), .Z(n27264) );
  XOR U27187 ( .A(n27278), .B(n27279), .Z(n27266) );
  XOR U27188 ( .A(n27280), .B(n27281), .Z(n27279) );
  XNOR U27189 ( .A(n27282), .B(n27283), .Z(n27278) );
  ANDN U27190 ( .B(n26970), .A(n27057), .Z(n27282) );
  AND U27191 ( .A(n27257), .B(n27260), .Z(n27277) );
  XNOR U27192 ( .A(n27257), .B(n27260), .Z(n27272) );
  XNOR U27193 ( .A(n27284), .B(n27285), .Z(n27260) );
  XNOR U27194 ( .A(n27286), .B(n27287), .Z(n27285) );
  XOR U27195 ( .A(n27280), .B(n27288), .Z(n27284) );
  XNOR U27196 ( .A(n27289), .B(n27283), .Z(n27288) );
  OR U27197 ( .A(n27056), .B(n27245), .Z(n27283) );
  XNOR U27198 ( .A(n27290), .B(n27243), .Z(n27245) );
  XNOR U27199 ( .A(n27057), .B(n27291), .Z(n27056) );
  NOR U27200 ( .A(n27291), .B(n27243), .Z(n27289) );
  XNOR U27201 ( .A(n27292), .B(n27293), .Z(n27257) );
  XNOR U27202 ( .A(n27294), .B(n27295), .Z(n27293) );
  XOR U27203 ( .A(n27065), .B(n27280), .Z(n27295) );
  XOR U27204 ( .A(n26970), .B(n27296), .Z(n27280) );
  XNOR U27205 ( .A(n26916), .B(n27297), .Z(n27292) );
  XNOR U27206 ( .A(n27298), .B(n27299), .Z(n27297) );
  ANDN U27207 ( .B(n27062), .A(n27300), .Z(n27298) );
  XNOR U27208 ( .A(n27301), .B(n27302), .Z(n27271) );
  XNOR U27209 ( .A(n27281), .B(n27303), .Z(n27302) );
  XNOR U27210 ( .A(n27062), .B(n27287), .Z(n27303) );
  XOR U27211 ( .A(n27243), .B(n27291), .Z(n27287) );
  XNOR U27212 ( .A(n27294), .B(n27304), .Z(n27281) );
  XNOR U27213 ( .A(n27305), .B(n27306), .Z(n27304) );
  NANDN U27214 ( .A(n27071), .B(n26977), .Z(n27306) );
  IV U27215 ( .A(n27286), .Z(n27294) );
  XNOR U27216 ( .A(n27307), .B(n27305), .Z(n27286) );
  NANDN U27217 ( .A(n27252), .B(n27074), .Z(n27305) );
  XOR U27218 ( .A(n27062), .B(n27291), .Z(n27071) );
  IV U27219 ( .A(n26920), .Z(n27291) );
  XOR U27220 ( .A(n27308), .B(n27309), .Z(n26920) );
  XNOR U27221 ( .A(n27310), .B(n27311), .Z(n27309) );
  XOR U27222 ( .A(n27261), .B(n26977), .Z(n27252) );
  XNOR U27223 ( .A(n27250), .B(n27243), .Z(n26977) );
  XNOR U27224 ( .A(n27311), .B(n27308), .Z(n27243) );
  ANDN U27225 ( .B(n27075), .A(n27261), .Z(n27307) );
  XNOR U27226 ( .A(n27312), .B(n26970), .Z(n27261) );
  IV U27227 ( .A(n27290), .Z(n26970) );
  XNOR U27228 ( .A(n27313), .B(n27314), .Z(n27290) );
  XNOR U27229 ( .A(n27315), .B(n27311), .Z(n27314) );
  XOR U27230 ( .A(n27316), .B(n27296), .Z(n27075) );
  XNOR U27231 ( .A(n27300), .B(n27317), .Z(n27301) );
  XNOR U27232 ( .A(n27318), .B(n27299), .Z(n27317) );
  OR U27233 ( .A(n27067), .B(n27248), .Z(n27299) );
  XOR U27234 ( .A(n26916), .B(n27250), .Z(n27248) );
  IV U27235 ( .A(n27300), .Z(n27250) );
  XOR U27236 ( .A(n27065), .B(n27062), .Z(n27067) );
  XNOR U27237 ( .A(n27296), .B(n27319), .Z(n27062) );
  XNOR U27238 ( .A(n27310), .B(n27313), .Z(n27319) );
  XNOR U27239 ( .A(msg[58]), .B(key[58]), .Z(n27313) );
  IV U27240 ( .A(n27057), .Z(n27296) );
  XOR U27241 ( .A(n27320), .B(n27321), .Z(n27057) );
  XOR U27242 ( .A(n27311), .B(n27322), .Z(n27321) );
  IV U27243 ( .A(n27316), .Z(n27065) );
  ANDN U27244 ( .B(n27316), .A(n26916), .Z(n27318) );
  XOR U27245 ( .A(n27308), .B(n27323), .Z(n27316) );
  XNOR U27246 ( .A(n27311), .B(n27324), .Z(n27323) );
  XOR U27247 ( .A(n27312), .B(n27325), .Z(n27311) );
  XNOR U27248 ( .A(msg[62]), .B(key[62]), .Z(n27325) );
  IV U27249 ( .A(n27320), .Z(n27308) );
  XOR U27250 ( .A(msg[61]), .B(key[61]), .Z(n27320) );
  XOR U27251 ( .A(n27326), .B(n27327), .Z(n27300) );
  XOR U27252 ( .A(n27324), .B(n27322), .Z(n27327) );
  XOR U27253 ( .A(msg[63]), .B(key[63]), .Z(n27322) );
  XNOR U27254 ( .A(msg[60]), .B(key[60]), .Z(n27324) );
  XOR U27255 ( .A(n26916), .B(n27315), .Z(n27326) );
  XNOR U27256 ( .A(n27310), .B(n27328), .Z(n27315) );
  XNOR U27257 ( .A(msg[59]), .B(key[59]), .Z(n27328) );
  XNOR U27258 ( .A(msg[57]), .B(key[57]), .Z(n27310) );
  IV U27259 ( .A(n27312), .Z(n26916) );
  XOR U27260 ( .A(msg[56]), .B(key[56]), .Z(n27312) );
  XOR U27261 ( .A(n26954), .B(n27031), .Z(n26299) );
  XNOR U27262 ( .A(n26960), .B(n27329), .Z(n27031) );
  XNOR U27263 ( .A(n26957), .B(n27330), .Z(n27329) );
  NANDN U27264 ( .A(n27331), .B(n27332), .Z(n27330) );
  OR U27265 ( .A(n27333), .B(n27081), .Z(n26957) );
  XNOR U27266 ( .A(n26959), .B(n27332), .Z(n27081) );
  XOR U27267 ( .A(n27335), .B(n26927), .Z(n27334) );
  OR U27268 ( .A(n27092), .B(n27336), .Z(n26927) );
  XOR U27269 ( .A(n26929), .B(n27337), .Z(n27092) );
  ANDN U27270 ( .B(n27338), .A(n27087), .Z(n27335) );
  XNOR U27271 ( .A(n27339), .B(n26962), .Z(n26960) );
  OR U27272 ( .A(n27099), .B(n27340), .Z(n26962) );
  XOR U27273 ( .A(n27341), .B(n26964), .Z(n27099) );
  XOR U27274 ( .A(n27337), .B(n26935), .Z(n26964) );
  IV U27275 ( .A(n27332), .Z(n26935) );
  XOR U27276 ( .A(n27342), .B(n27343), .Z(n27332) );
  NANDN U27277 ( .A(n27344), .B(n27345), .Z(n27343) );
  IV U27278 ( .A(n27087), .Z(n27337) );
  XNOR U27279 ( .A(n27346), .B(n27347), .Z(n27087) );
  NANDN U27280 ( .A(n27344), .B(n27348), .Z(n27347) );
  ANDN U27281 ( .B(n27341), .A(n27349), .Z(n27339) );
  IV U27282 ( .A(n27102), .Z(n27341) );
  XOR U27283 ( .A(n26959), .B(n26929), .Z(n27102) );
  XOR U27284 ( .A(n27350), .B(n27346), .Z(n26929) );
  NANDN U27285 ( .A(n27351), .B(n27352), .Z(n27346) );
  NANDN U27286 ( .A(n27351), .B(n27356), .Z(n27342) );
  XOR U27287 ( .A(n27357), .B(n27358), .Z(n27344) );
  XOR U27288 ( .A(n27359), .B(n27354), .Z(n27358) );
  XNOR U27289 ( .A(n27360), .B(n27361), .Z(n27357) );
  XNOR U27290 ( .A(n27362), .B(n27363), .Z(n27361) );
  ANDN U27291 ( .B(n27359), .A(n27354), .Z(n27362) );
  ANDN U27292 ( .B(n27359), .A(n27353), .Z(n27355) );
  XNOR U27293 ( .A(n27360), .B(n27364), .Z(n27353) );
  XOR U27294 ( .A(n27365), .B(n27363), .Z(n27364) );
  NAND U27295 ( .A(n27352), .B(n27356), .Z(n27363) );
  XNOR U27296 ( .A(n27348), .B(n27354), .Z(n27352) );
  XOR U27297 ( .A(n27366), .B(n27367), .Z(n27354) );
  XOR U27298 ( .A(n27368), .B(n27369), .Z(n27367) );
  XNOR U27299 ( .A(n27370), .B(n27371), .Z(n27366) );
  ANDN U27300 ( .B(n26958), .A(n27083), .Z(n27370) );
  AND U27301 ( .A(n27345), .B(n27348), .Z(n27365) );
  XNOR U27302 ( .A(n27345), .B(n27348), .Z(n27360) );
  XNOR U27303 ( .A(n27372), .B(n27373), .Z(n27348) );
  XNOR U27304 ( .A(n27374), .B(n27375), .Z(n27373) );
  XOR U27305 ( .A(n27368), .B(n27376), .Z(n27372) );
  XNOR U27306 ( .A(n27377), .B(n27371), .Z(n27376) );
  OR U27307 ( .A(n27082), .B(n27333), .Z(n27371) );
  XNOR U27308 ( .A(n27378), .B(n27331), .Z(n27333) );
  XNOR U27309 ( .A(n27083), .B(n27379), .Z(n27082) );
  NOR U27310 ( .A(n27379), .B(n27331), .Z(n27377) );
  XNOR U27311 ( .A(n27380), .B(n27381), .Z(n27345) );
  XNOR U27312 ( .A(n27382), .B(n27383), .Z(n27381) );
  XOR U27313 ( .A(n27091), .B(n27368), .Z(n27383) );
  XOR U27314 ( .A(n26958), .B(n27384), .Z(n27368) );
  XNOR U27315 ( .A(n26930), .B(n27385), .Z(n27380) );
  XNOR U27316 ( .A(n27386), .B(n27387), .Z(n27385) );
  ANDN U27317 ( .B(n27088), .A(n27388), .Z(n27386) );
  XNOR U27318 ( .A(n27389), .B(n27390), .Z(n27359) );
  XNOR U27319 ( .A(n27369), .B(n27391), .Z(n27390) );
  XNOR U27320 ( .A(n27088), .B(n27375), .Z(n27391) );
  XOR U27321 ( .A(n27331), .B(n27379), .Z(n27375) );
  XNOR U27322 ( .A(n27382), .B(n27392), .Z(n27369) );
  XNOR U27323 ( .A(n27393), .B(n27394), .Z(n27392) );
  NANDN U27324 ( .A(n27097), .B(n26965), .Z(n27394) );
  IV U27325 ( .A(n27374), .Z(n27382) );
  XNOR U27326 ( .A(n27395), .B(n27393), .Z(n27374) );
  NANDN U27327 ( .A(n27340), .B(n27100), .Z(n27393) );
  XOR U27328 ( .A(n27088), .B(n27379), .Z(n27097) );
  IV U27329 ( .A(n26934), .Z(n27379) );
  XOR U27330 ( .A(n27396), .B(n27397), .Z(n26934) );
  XNOR U27331 ( .A(n27398), .B(n27399), .Z(n27397) );
  XOR U27332 ( .A(n27349), .B(n26965), .Z(n27340) );
  XNOR U27333 ( .A(n27338), .B(n27331), .Z(n26965) );
  XNOR U27334 ( .A(n27399), .B(n27396), .Z(n27331) );
  ANDN U27335 ( .B(n27101), .A(n27349), .Z(n27395) );
  XNOR U27336 ( .A(n27400), .B(n26958), .Z(n27349) );
  IV U27337 ( .A(n27378), .Z(n26958) );
  XNOR U27338 ( .A(n27401), .B(n27402), .Z(n27378) );
  XNOR U27339 ( .A(n27403), .B(n27399), .Z(n27402) );
  XOR U27340 ( .A(n27404), .B(n27384), .Z(n27101) );
  XNOR U27341 ( .A(n27388), .B(n27405), .Z(n27389) );
  XNOR U27342 ( .A(n27406), .B(n27387), .Z(n27405) );
  OR U27343 ( .A(n27093), .B(n27336), .Z(n27387) );
  XOR U27344 ( .A(n26930), .B(n27338), .Z(n27336) );
  IV U27345 ( .A(n27388), .Z(n27338) );
  XOR U27346 ( .A(n27091), .B(n27088), .Z(n27093) );
  XNOR U27347 ( .A(n27384), .B(n27407), .Z(n27088) );
  XNOR U27348 ( .A(n27398), .B(n27401), .Z(n27407) );
  XNOR U27349 ( .A(msg[66]), .B(key[66]), .Z(n27401) );
  IV U27350 ( .A(n27083), .Z(n27384) );
  XOR U27351 ( .A(n27408), .B(n27409), .Z(n27083) );
  XOR U27352 ( .A(n27399), .B(n27410), .Z(n27409) );
  IV U27353 ( .A(n27404), .Z(n27091) );
  ANDN U27354 ( .B(n27404), .A(n26930), .Z(n27406) );
  XOR U27355 ( .A(n27396), .B(n27411), .Z(n27404) );
  XNOR U27356 ( .A(n27399), .B(n27412), .Z(n27411) );
  XOR U27357 ( .A(n27400), .B(n27413), .Z(n27399) );
  XNOR U27358 ( .A(msg[70]), .B(key[70]), .Z(n27413) );
  IV U27359 ( .A(n27408), .Z(n27396) );
  XOR U27360 ( .A(msg[69]), .B(key[69]), .Z(n27408) );
  XOR U27361 ( .A(n27414), .B(n27415), .Z(n27388) );
  XOR U27362 ( .A(n27412), .B(n27410), .Z(n27415) );
  XOR U27363 ( .A(msg[71]), .B(key[71]), .Z(n27410) );
  XNOR U27364 ( .A(msg[68]), .B(key[68]), .Z(n27412) );
  XOR U27365 ( .A(n26930), .B(n27403), .Z(n27414) );
  XNOR U27366 ( .A(n27398), .B(n27416), .Z(n27403) );
  XNOR U27367 ( .A(msg[67]), .B(key[67]), .Z(n27416) );
  XNOR U27368 ( .A(msg[65]), .B(key[65]), .Z(n27398) );
  IV U27369 ( .A(n27400), .Z(n26930) );
  XOR U27370 ( .A(msg[64]), .B(key[64]), .Z(n27400) );
  XNOR U27371 ( .A(key[178]), .B(n24647), .Z(n27103) );
  IV U27372 ( .A(n27020), .Z(n24647) );
  XOR U27373 ( .A(n26999), .B(n27036), .Z(n27020) );
  XOR U27374 ( .A(n27418), .B(n26995), .Z(n27417) );
  OR U27375 ( .A(n27419), .B(n27121), .Z(n26995) );
  XNOR U27376 ( .A(n26997), .B(n27116), .Z(n27121) );
  NOR U27377 ( .A(n27420), .B(n27116), .Z(n27418) );
  IV U27378 ( .A(n27035), .Z(n26999) );
  XOR U27379 ( .A(n27044), .B(n27421), .Z(n27035) );
  XNOR U27380 ( .A(n27041), .B(n27422), .Z(n27421) );
  NANDN U27381 ( .A(n27423), .B(n27424), .Z(n27422) );
  OR U27382 ( .A(n27425), .B(n27110), .Z(n27041) );
  XNOR U27383 ( .A(n27042), .B(n27424), .Z(n27110) );
  XNOR U27384 ( .A(n27426), .B(n27046), .Z(n27044) );
  OR U27385 ( .A(n27128), .B(n27427), .Z(n27046) );
  XNOR U27386 ( .A(n27428), .B(n27048), .Z(n27128) );
  XNOR U27387 ( .A(n27116), .B(n27424), .Z(n27048) );
  IV U27388 ( .A(n26945), .Z(n27424) );
  XNOR U27389 ( .A(n27429), .B(n27430), .Z(n26945) );
  NANDN U27390 ( .A(n27431), .B(n27432), .Z(n27430) );
  XNOR U27391 ( .A(n27433), .B(n27434), .Z(n27116) );
  NANDN U27392 ( .A(n27431), .B(n27435), .Z(n27434) );
  ANDN U27393 ( .B(n27428), .A(n27436), .Z(n27426) );
  IV U27394 ( .A(n27131), .Z(n27428) );
  XOR U27395 ( .A(n26997), .B(n27042), .Z(n27131) );
  XNOR U27396 ( .A(n27437), .B(n27429), .Z(n27042) );
  NANDN U27397 ( .A(n27438), .B(n27439), .Z(n27429) );
  XOR U27398 ( .A(n27432), .B(n27440), .Z(n27439) );
  ANDN U27399 ( .B(n27440), .A(n27441), .Z(n27437) );
  NANDN U27400 ( .A(n27438), .B(n27443), .Z(n27433) );
  XOR U27401 ( .A(n27444), .B(n27445), .Z(n27431) );
  XOR U27402 ( .A(n27446), .B(n27447), .Z(n27445) );
  XNOR U27403 ( .A(n27448), .B(n27449), .Z(n27444) );
  XNOR U27404 ( .A(n27450), .B(n27451), .Z(n27449) );
  ANDN U27405 ( .B(n27447), .A(n27446), .Z(n27450) );
  ANDN U27406 ( .B(n27447), .A(n27441), .Z(n27442) );
  XNOR U27407 ( .A(n27448), .B(n27452), .Z(n27441) );
  XOR U27408 ( .A(n27453), .B(n27451), .Z(n27452) );
  NAND U27409 ( .A(n27443), .B(n27454), .Z(n27451) );
  XNOR U27410 ( .A(n27432), .B(n27446), .Z(n27454) );
  IV U27411 ( .A(n27440), .Z(n27446) );
  XNOR U27412 ( .A(n27455), .B(n27456), .Z(n27440) );
  XNOR U27413 ( .A(n27457), .B(n27458), .Z(n27456) );
  XOR U27414 ( .A(n27117), .B(n27459), .Z(n27458) );
  XNOR U27415 ( .A(n27420), .B(n27460), .Z(n27455) );
  XNOR U27416 ( .A(n27461), .B(n27462), .Z(n27460) );
  AND U27417 ( .A(n27120), .B(n26998), .Z(n27461) );
  XOR U27418 ( .A(n27435), .B(n27447), .Z(n27443) );
  AND U27419 ( .A(n27432), .B(n27435), .Z(n27453) );
  XNOR U27420 ( .A(n27432), .B(n27435), .Z(n27448) );
  XNOR U27421 ( .A(n27463), .B(n27464), .Z(n27435) );
  XNOR U27422 ( .A(n27465), .B(n27459), .Z(n27464) );
  XOR U27423 ( .A(n27466), .B(n27467), .Z(n27463) );
  XNOR U27424 ( .A(n27468), .B(n27469), .Z(n27467) );
  ANDN U27425 ( .B(n26944), .A(n27423), .Z(n27468) );
  XNOR U27426 ( .A(n27470), .B(n27471), .Z(n27432) );
  XNOR U27427 ( .A(n27120), .B(n27466), .Z(n27472) );
  XOR U27428 ( .A(n26998), .B(n27473), .Z(n27470) );
  XNOR U27429 ( .A(n27474), .B(n27462), .Z(n27473) );
  OR U27430 ( .A(n27122), .B(n27419), .Z(n27462) );
  XOR U27431 ( .A(n26998), .B(n27420), .Z(n27419) );
  XNOR U27432 ( .A(n27120), .B(n27475), .Z(n27122) );
  ANDN U27433 ( .B(n27476), .A(n27117), .Z(n27474) );
  XNOR U27434 ( .A(n27477), .B(n27478), .Z(n27447) );
  XOR U27435 ( .A(n27465), .B(n27457), .Z(n27478) );
  XOR U27436 ( .A(n27466), .B(n27479), .Z(n27457) );
  XNOR U27437 ( .A(n27480), .B(n27481), .Z(n27479) );
  NAND U27438 ( .A(n27049), .B(n27126), .Z(n27481) );
  XNOR U27439 ( .A(n27482), .B(n27480), .Z(n27466) );
  NANDN U27440 ( .A(n27427), .B(n27129), .Z(n27480) );
  XOR U27441 ( .A(n27130), .B(n27126), .Z(n27129) );
  XOR U27442 ( .A(n27475), .B(n26944), .Z(n27126) );
  IV U27443 ( .A(n27117), .Z(n27475) );
  XOR U27444 ( .A(n27483), .B(n27484), .Z(n27117) );
  XNOR U27445 ( .A(n27485), .B(n27486), .Z(n27484) );
  XOR U27446 ( .A(n27436), .B(n27049), .Z(n27427) );
  XNOR U27447 ( .A(n27476), .B(n27423), .Z(n27049) );
  IV U27448 ( .A(n27420), .Z(n27476) );
  XOR U27449 ( .A(n27487), .B(n27488), .Z(n27420) );
  XOR U27450 ( .A(n27489), .B(n27490), .Z(n27488) );
  XNOR U27451 ( .A(n26998), .B(n27491), .Z(n27487) );
  ANDN U27452 ( .B(n27130), .A(n27436), .Z(n27482) );
  XNOR U27453 ( .A(n26998), .B(n27492), .Z(n27436) );
  XOR U27454 ( .A(n27120), .B(n27483), .Z(n27130) );
  XOR U27455 ( .A(n27493), .B(n27494), .Z(n27120) );
  XOR U27456 ( .A(n27495), .B(n27490), .Z(n27494) );
  XOR U27457 ( .A(msg[108]), .B(key[108]), .Z(n27490) );
  XNOR U27458 ( .A(n27492), .B(n27112), .Z(n27465) );
  XNOR U27459 ( .A(n27496), .B(n27469), .Z(n27477) );
  OR U27460 ( .A(n27111), .B(n27425), .Z(n27469) );
  XNOR U27461 ( .A(n27043), .B(n27423), .Z(n27425) );
  XOR U27462 ( .A(n27497), .B(n27493), .Z(n27423) );
  XNOR U27463 ( .A(n27483), .B(n26944), .Z(n27111) );
  XOR U27464 ( .A(n27493), .B(n27498), .Z(n26944) );
  XOR U27465 ( .A(n27485), .B(n27497), .Z(n27498) );
  IV U27466 ( .A(n27112), .Z(n27483) );
  ANDN U27467 ( .B(n27492), .A(n27112), .Z(n27496) );
  XNOR U27468 ( .A(n27493), .B(n27499), .Z(n27112) );
  XNOR U27469 ( .A(n27495), .B(n27489), .Z(n27499) );
  XNOR U27470 ( .A(msg[111]), .B(key[111]), .Z(n27489) );
  XNOR U27471 ( .A(msg[109]), .B(key[109]), .Z(n27493) );
  IV U27472 ( .A(n27043), .Z(n27492) );
  XNOR U27473 ( .A(n27486), .B(n27500), .Z(n27043) );
  XOR U27474 ( .A(n27491), .B(n27497), .Z(n27500) );
  IV U27475 ( .A(n27495), .Z(n27497) );
  XOR U27476 ( .A(n26998), .B(n27501), .Z(n27495) );
  XNOR U27477 ( .A(msg[110]), .B(key[110]), .Z(n27501) );
  XOR U27478 ( .A(msg[104]), .B(key[104]), .Z(n26998) );
  XNOR U27479 ( .A(n27485), .B(n27502), .Z(n27491) );
  XNOR U27480 ( .A(msg[107]), .B(key[107]), .Z(n27502) );
  XNOR U27481 ( .A(msg[105]), .B(key[105]), .Z(n27485) );
  XNOR U27482 ( .A(msg[106]), .B(key[106]), .Z(n27486) );
  XNOR U27483 ( .A(n26588), .B(n26664), .Z(n22246) );
  XNOR U27484 ( .A(n26724), .B(n27503), .Z(n26664) );
  XOR U27485 ( .A(n27504), .B(n26624), .Z(n27503) );
  OR U27486 ( .A(n27505), .B(n26744), .Z(n26624) );
  XNOR U27487 ( .A(n26627), .B(n26743), .Z(n26744) );
  ANDN U27488 ( .B(n27506), .A(n27507), .Z(n27504) );
  XNOR U27489 ( .A(n26622), .B(n27508), .Z(n26588) );
  XNOR U27490 ( .A(n27509), .B(n26726), .Z(n27508) );
  XOR U27491 ( .A(n27511), .B(n26592), .Z(n26731) );
  ANDN U27492 ( .B(n27512), .A(n26734), .Z(n27509) );
  IV U27493 ( .A(n27511), .Z(n26734) );
  XNOR U27494 ( .A(n26724), .B(n27513), .Z(n26622) );
  XNOR U27495 ( .A(n27514), .B(n27515), .Z(n27513) );
  NANDN U27496 ( .A(n26738), .B(n27516), .Z(n27515) );
  XOR U27497 ( .A(n27517), .B(n27514), .Z(n26724) );
  OR U27498 ( .A(n26747), .B(n27518), .Z(n27514) );
  XNOR U27499 ( .A(n26750), .B(n26738), .Z(n26747) );
  XNOR U27500 ( .A(n26743), .B(n26592), .Z(n26738) );
  XOR U27501 ( .A(n27519), .B(n27520), .Z(n26592) );
  NANDN U27502 ( .A(n27521), .B(n27522), .Z(n27520) );
  IV U27503 ( .A(n27507), .Z(n26743) );
  XNOR U27504 ( .A(n27523), .B(n27524), .Z(n27507) );
  NANDN U27505 ( .A(n27521), .B(n27525), .Z(n27524) );
  NOR U27506 ( .A(n26750), .B(n27526), .Z(n27517) );
  XNOR U27507 ( .A(n27511), .B(n26627), .Z(n26750) );
  XNOR U27508 ( .A(n27527), .B(n27523), .Z(n26627) );
  NANDN U27509 ( .A(n27528), .B(n27529), .Z(n27523) );
  XOR U27510 ( .A(n27525), .B(n27530), .Z(n27529) );
  ANDN U27511 ( .B(n27530), .A(n27531), .Z(n27527) );
  XNOR U27512 ( .A(n27532), .B(n27519), .Z(n27511) );
  NANDN U27513 ( .A(n27528), .B(n27533), .Z(n27519) );
  XOR U27514 ( .A(n27534), .B(n27522), .Z(n27533) );
  XNOR U27515 ( .A(n27535), .B(n27536), .Z(n27521) );
  XOR U27516 ( .A(n27537), .B(n27538), .Z(n27536) );
  XNOR U27517 ( .A(n27539), .B(n27540), .Z(n27535) );
  XNOR U27518 ( .A(n27541), .B(n27542), .Z(n27540) );
  ANDN U27519 ( .B(n27534), .A(n27538), .Z(n27541) );
  ANDN U27520 ( .B(n27534), .A(n27531), .Z(n27532) );
  XNOR U27521 ( .A(n27537), .B(n27543), .Z(n27531) );
  XOR U27522 ( .A(n27544), .B(n27542), .Z(n27543) );
  NAND U27523 ( .A(n27545), .B(n27546), .Z(n27542) );
  XNOR U27524 ( .A(n27539), .B(n27522), .Z(n27546) );
  IV U27525 ( .A(n27534), .Z(n27539) );
  XNOR U27526 ( .A(n27525), .B(n27538), .Z(n27545) );
  IV U27527 ( .A(n27530), .Z(n27538) );
  XOR U27528 ( .A(n27547), .B(n27548), .Z(n27530) );
  XNOR U27529 ( .A(n27549), .B(n27550), .Z(n27548) );
  XNOR U27530 ( .A(n27551), .B(n27552), .Z(n27547) );
  ANDN U27531 ( .B(n27512), .A(n27553), .Z(n27551) );
  AND U27532 ( .A(n27522), .B(n27525), .Z(n27544) );
  XNOR U27533 ( .A(n27522), .B(n27525), .Z(n27537) );
  XNOR U27534 ( .A(n27554), .B(n27555), .Z(n27525) );
  XNOR U27535 ( .A(n27556), .B(n27550), .Z(n27555) );
  XOR U27536 ( .A(n27557), .B(n27558), .Z(n27554) );
  XNOR U27537 ( .A(n27559), .B(n27552), .Z(n27558) );
  OR U27538 ( .A(n26732), .B(n27510), .Z(n27552) );
  XNOR U27539 ( .A(n27512), .B(n27560), .Z(n27510) );
  XNOR U27540 ( .A(n27553), .B(n26593), .Z(n26732) );
  ANDN U27541 ( .B(n27561), .A(n26728), .Z(n27559) );
  XNOR U27542 ( .A(n27562), .B(n27563), .Z(n27522) );
  XNOR U27543 ( .A(n27550), .B(n27564), .Z(n27563) );
  XOR U27544 ( .A(n26723), .B(n27557), .Z(n27564) );
  XNOR U27545 ( .A(n27512), .B(n27553), .Z(n27550) );
  XNOR U27546 ( .A(n27565), .B(n27566), .Z(n27562) );
  XNOR U27547 ( .A(n27567), .B(n27568), .Z(n27566) );
  ANDN U27548 ( .B(n27506), .A(n26742), .Z(n27567) );
  XNOR U27549 ( .A(n27569), .B(n27570), .Z(n27534) );
  XNOR U27550 ( .A(n27556), .B(n27571), .Z(n27570) );
  XNOR U27551 ( .A(n26742), .B(n27549), .Z(n27571) );
  XOR U27552 ( .A(n27557), .B(n27572), .Z(n27549) );
  XNOR U27553 ( .A(n27573), .B(n27574), .Z(n27572) );
  NAND U27554 ( .A(n27516), .B(n26739), .Z(n27574) );
  XNOR U27555 ( .A(n27575), .B(n27573), .Z(n27557) );
  NANDN U27556 ( .A(n27518), .B(n26748), .Z(n27573) );
  XOR U27557 ( .A(n26749), .B(n26739), .Z(n26748) );
  XNOR U27558 ( .A(n27576), .B(n26593), .Z(n26739) );
  XOR U27559 ( .A(n27526), .B(n27516), .Z(n27518) );
  XOR U27560 ( .A(n27506), .B(n27560), .Z(n27516) );
  ANDN U27561 ( .B(n26749), .A(n27526), .Z(n27575) );
  XNOR U27562 ( .A(n27565), .B(n27512), .Z(n27526) );
  XNOR U27563 ( .A(n27577), .B(n27578), .Z(n27512) );
  XNOR U27564 ( .A(n27579), .B(n27580), .Z(n27578) );
  XOR U27565 ( .A(n27581), .B(n26733), .Z(n26749) );
  XOR U27566 ( .A(n27560), .B(n27561), .Z(n27556) );
  IV U27567 ( .A(n26593), .Z(n27561) );
  XOR U27568 ( .A(n27582), .B(n27583), .Z(n26593) );
  XNOR U27569 ( .A(n27584), .B(n27580), .Z(n27583) );
  IV U27570 ( .A(n26728), .Z(n27560) );
  XOR U27571 ( .A(n27580), .B(n27585), .Z(n26728) );
  XNOR U27572 ( .A(n27506), .B(n27586), .Z(n27569) );
  XNOR U27573 ( .A(n27587), .B(n27568), .Z(n27586) );
  OR U27574 ( .A(n26745), .B(n27505), .Z(n27568) );
  XNOR U27575 ( .A(n27565), .B(n27506), .Z(n27505) );
  XOR U27576 ( .A(n26723), .B(n27576), .Z(n26745) );
  IV U27577 ( .A(n26742), .Z(n27576) );
  XOR U27578 ( .A(n26733), .B(n27588), .Z(n26742) );
  XNOR U27579 ( .A(n27584), .B(n27577), .Z(n27588) );
  XOR U27580 ( .A(n27589), .B(n27590), .Z(n27577) );
  XOR U27581 ( .A(n25246), .B(n25243), .Z(n27590) );
  XOR U27582 ( .A(n24227), .B(n27591), .Z(n27589) );
  XNOR U27583 ( .A(key[218]), .B(n26046), .Z(n27591) );
  XOR U27584 ( .A(n27592), .B(n27593), .Z(n26046) );
  XNOR U27585 ( .A(n27594), .B(n27595), .Z(n27592) );
  XNOR U27586 ( .A(n24189), .B(n25202), .Z(n24227) );
  IV U27587 ( .A(n27553), .Z(n26733) );
  XOR U27588 ( .A(n27582), .B(n27596), .Z(n27553) );
  XOR U27589 ( .A(n27580), .B(n27597), .Z(n27596) );
  ANDN U27590 ( .B(n27581), .A(n26626), .Z(n27587) );
  IV U27591 ( .A(n26723), .Z(n27581) );
  XOR U27592 ( .A(n27582), .B(n27598), .Z(n26723) );
  XOR U27593 ( .A(n27580), .B(n27599), .Z(n27598) );
  XOR U27594 ( .A(n27600), .B(n27601), .Z(n27580) );
  XNOR U27595 ( .A(n26053), .B(n26626), .Z(n27601) );
  IV U27596 ( .A(n27565), .Z(n26626) );
  XNOR U27597 ( .A(n24203), .B(n26065), .Z(n26053) );
  XNOR U27598 ( .A(n24236), .B(n25231), .Z(n26065) );
  XNOR U27599 ( .A(n27602), .B(n27603), .Z(n25231) );
  XOR U27600 ( .A(n27604), .B(n27605), .Z(n27603) );
  XOR U27601 ( .A(n27606), .B(n27607), .Z(n27602) );
  XOR U27602 ( .A(n25222), .B(n25212), .Z(n24203) );
  IV U27603 ( .A(n24196), .Z(n25222) );
  XOR U27604 ( .A(n27608), .B(n27609), .Z(n24196) );
  XOR U27605 ( .A(n24197), .B(n27610), .Z(n27600) );
  XOR U27606 ( .A(key[222]), .B(n25224), .Z(n27610) );
  XOR U27607 ( .A(n27611), .B(n27612), .Z(n25224) );
  XNOR U27608 ( .A(n27613), .B(n27614), .Z(n27612) );
  XOR U27609 ( .A(n27615), .B(n25229), .Z(n24197) );
  IV U27610 ( .A(n27585), .Z(n27582) );
  XOR U27611 ( .A(n27616), .B(n27617), .Z(n27585) );
  XOR U27612 ( .A(n25212), .B(n26060), .Z(n27617) );
  XOR U27613 ( .A(n24204), .B(n25219), .Z(n26060) );
  XOR U27614 ( .A(n27618), .B(n27619), .Z(n24204) );
  XNOR U27615 ( .A(n27620), .B(n27621), .Z(n27619) );
  XNOR U27616 ( .A(n27622), .B(n27623), .Z(n27618) );
  XNOR U27617 ( .A(n27624), .B(n27625), .Z(n27623) );
  ANDN U27618 ( .B(n27626), .A(n27627), .Z(n27625) );
  XOR U27619 ( .A(n25220), .B(n27630), .Z(n27616) );
  XNOR U27620 ( .A(key[221]), .B(n26055), .Z(n27630) );
  XNOR U27621 ( .A(n27595), .B(n27631), .Z(n26055) );
  XNOR U27622 ( .A(n27632), .B(n27633), .Z(n27595) );
  XOR U27623 ( .A(n27634), .B(n27635), .Z(n27633) );
  NOR U27624 ( .A(n27636), .B(n27637), .Z(n27634) );
  XNOR U27625 ( .A(n27638), .B(n27639), .Z(n25220) );
  XNOR U27626 ( .A(n27640), .B(n27641), .Z(n27639) );
  XNOR U27627 ( .A(n27642), .B(n27643), .Z(n27638) );
  XNOR U27628 ( .A(n27644), .B(n27645), .Z(n27643) );
  ANDN U27629 ( .B(n27646), .A(n27647), .Z(n27644) );
  XOR U27630 ( .A(n27648), .B(n27649), .Z(n27506) );
  XNOR U27631 ( .A(n27599), .B(n27597), .Z(n27649) );
  XNOR U27632 ( .A(n27650), .B(n27651), .Z(n27597) );
  XOR U27633 ( .A(n25254), .B(n26066), .Z(n27651) );
  XOR U27634 ( .A(n25216), .B(n25229), .Z(n26066) );
  XNOR U27635 ( .A(n27652), .B(n27653), .Z(n25229) );
  XOR U27636 ( .A(n27629), .B(n27654), .Z(n27653) );
  XOR U27637 ( .A(n27655), .B(n27656), .Z(n27652) );
  XOR U27638 ( .A(n27657), .B(n27658), .Z(n25216) );
  XNOR U27639 ( .A(n27609), .B(n27621), .Z(n27658) );
  XNOR U27640 ( .A(n27659), .B(n27660), .Z(n27621) );
  XNOR U27641 ( .A(n27661), .B(n27662), .Z(n27660) );
  NANDN U27642 ( .A(n27663), .B(n27664), .Z(n27662) );
  XOR U27643 ( .A(n27665), .B(n27666), .Z(n27657) );
  XOR U27644 ( .A(n27667), .B(n27615), .Z(n25254) );
  XNOR U27645 ( .A(key[223]), .B(n26057), .Z(n27650) );
  XOR U27646 ( .A(n27668), .B(n27669), .Z(n26057) );
  XNOR U27647 ( .A(n27670), .B(n27641), .Z(n27669) );
  XNOR U27648 ( .A(n27671), .B(n27672), .Z(n27641) );
  XNOR U27649 ( .A(n27673), .B(n27674), .Z(n27672) );
  NANDN U27650 ( .A(n27675), .B(n27676), .Z(n27674) );
  XOR U27651 ( .A(n27677), .B(n27678), .Z(n27668) );
  XNOR U27652 ( .A(n27679), .B(n26068), .Z(n27599) );
  XNOR U27653 ( .A(n27680), .B(n27681), .Z(n26068) );
  XOR U27654 ( .A(n24218), .B(n25238), .Z(n27681) );
  XOR U27655 ( .A(n27620), .B(n24189), .Z(n24218) );
  XNOR U27656 ( .A(n27665), .B(n27682), .Z(n24189) );
  XNOR U27657 ( .A(n24236), .B(n25221), .Z(n27680) );
  XOR U27658 ( .A(n27683), .B(n27684), .Z(n25221) );
  XNOR U27659 ( .A(n27685), .B(n27605), .Z(n27684) );
  XNOR U27660 ( .A(n27686), .B(n27687), .Z(n27605) );
  XNOR U27661 ( .A(n27688), .B(n27689), .Z(n27687) );
  OR U27662 ( .A(n27690), .B(n27691), .Z(n27689) );
  XNOR U27663 ( .A(n27692), .B(n27693), .Z(n27683) );
  XNOR U27664 ( .A(n27635), .B(n27694), .Z(n27693) );
  ANDN U27665 ( .B(n27695), .A(n27696), .Z(n27694) );
  NANDN U27666 ( .A(n27697), .B(n27698), .Z(n27635) );
  IV U27667 ( .A(n27667), .Z(n24236) );
  XOR U27668 ( .A(n24215), .B(n27699), .Z(n27679) );
  XNOR U27669 ( .A(key[220]), .B(n25236), .Z(n27699) );
  XNOR U27670 ( .A(n27642), .B(n25246), .Z(n25236) );
  XOR U27671 ( .A(n27613), .B(n27677), .Z(n25246) );
  XOR U27672 ( .A(n27615), .B(n25219), .Z(n24215) );
  XNOR U27673 ( .A(n27700), .B(n27701), .Z(n25219) );
  XOR U27674 ( .A(n27702), .B(n27654), .Z(n27701) );
  XNOR U27675 ( .A(n27703), .B(n27704), .Z(n27654) );
  XNOR U27676 ( .A(n27705), .B(n27706), .Z(n27704) );
  NANDN U27677 ( .A(n27707), .B(n27708), .Z(n27706) );
  XOR U27678 ( .A(n27709), .B(n27710), .Z(n27700) );
  XOR U27679 ( .A(n27711), .B(n27712), .Z(n27710) );
  ANDN U27680 ( .B(n27713), .A(n27714), .Z(n27712) );
  XOR U27681 ( .A(n27565), .B(n27579), .Z(n27648) );
  XOR U27682 ( .A(n27715), .B(n27716), .Z(n27579) );
  XNOR U27683 ( .A(n27584), .B(n27717), .Z(n27716) );
  XOR U27684 ( .A(n24188), .B(n26072), .Z(n27717) );
  XOR U27685 ( .A(n27667), .B(n25235), .Z(n26072) );
  XOR U27686 ( .A(n27692), .B(n27718), .Z(n25235) );
  XOR U27687 ( .A(n27692), .B(n27719), .Z(n27667) );
  XNOR U27688 ( .A(n27686), .B(n27720), .Z(n27692) );
  XNOR U27689 ( .A(n27721), .B(n27722), .Z(n27720) );
  NOR U27690 ( .A(n27723), .B(n27637), .Z(n27721) );
  XNOR U27691 ( .A(n27724), .B(n27725), .Z(n27686) );
  XNOR U27692 ( .A(n27726), .B(n27727), .Z(n27725) );
  NANDN U27693 ( .A(n27728), .B(n27729), .Z(n27727) );
  IV U27694 ( .A(n26077), .Z(n24188) );
  XOR U27695 ( .A(n24229), .B(n25243), .Z(n26077) );
  XNOR U27696 ( .A(n27730), .B(n27731), .Z(n25243) );
  XOR U27697 ( .A(n27732), .B(n27628), .Z(n27731) );
  XNOR U27698 ( .A(n27733), .B(n27734), .Z(n27628) );
  XNOR U27699 ( .A(n27735), .B(n27711), .Z(n27734) );
  NOR U27700 ( .A(n27736), .B(n27737), .Z(n27711) );
  ANDN U27701 ( .B(n27738), .A(n27739), .Z(n27735) );
  XNOR U27702 ( .A(n27740), .B(n27656), .Z(n27730) );
  XNOR U27703 ( .A(n27741), .B(n27742), .Z(n24229) );
  XOR U27704 ( .A(n27743), .B(n27608), .Z(n27742) );
  XNOR U27705 ( .A(n27744), .B(n27745), .Z(n27608) );
  XOR U27706 ( .A(n27746), .B(n27624), .Z(n27745) );
  NANDN U27707 ( .A(n27747), .B(n27748), .Z(n27624) );
  ANDN U27708 ( .B(n27749), .A(n27750), .Z(n27746) );
  XNOR U27709 ( .A(n27751), .B(n27666), .Z(n27741) );
  XOR U27710 ( .A(n27752), .B(n27753), .Z(n27584) );
  XNOR U27711 ( .A(n25202), .B(n27718), .Z(n27753) );
  IV U27712 ( .A(n26045), .Z(n27718) );
  XNOR U27713 ( .A(n27719), .B(n27606), .Z(n26045) );
  XOR U27714 ( .A(n25253), .B(n27754), .Z(n27752) );
  XOR U27715 ( .A(key[217]), .B(n24235), .Z(n27754) );
  XOR U27716 ( .A(n27755), .B(n24228), .Z(n24235) );
  XOR U27717 ( .A(n27609), .B(n27756), .Z(n24228) );
  XOR U27718 ( .A(n27751), .B(n27666), .Z(n27756) );
  XOR U27719 ( .A(n27744), .B(n27757), .Z(n27666) );
  XOR U27720 ( .A(n27758), .B(n27759), .Z(n27757) );
  ANDN U27721 ( .B(n27760), .A(n27663), .Z(n27758) );
  XNOR U27722 ( .A(n27622), .B(n27761), .Z(n27744) );
  XNOR U27723 ( .A(n27762), .B(n27763), .Z(n27761) );
  NAND U27724 ( .A(n27764), .B(n27765), .Z(n27763) );
  IV U27725 ( .A(n27665), .Z(n27751) );
  XOR U27726 ( .A(n27766), .B(n27767), .Z(n27665) );
  XNOR U27727 ( .A(n27768), .B(n27769), .Z(n27767) );
  NANDN U27728 ( .A(n27770), .B(n27626), .Z(n27769) );
  XOR U27729 ( .A(n27682), .B(n27743), .Z(n27609) );
  XOR U27730 ( .A(n27622), .B(n27771), .Z(n27743) );
  XNOR U27731 ( .A(n27759), .B(n27772), .Z(n27771) );
  NANDN U27732 ( .A(n27773), .B(n27774), .Z(n27772) );
  OR U27733 ( .A(n27775), .B(n27776), .Z(n27759) );
  XOR U27734 ( .A(n27777), .B(n27762), .Z(n27622) );
  NANDN U27735 ( .A(n27778), .B(n27779), .Z(n27762) );
  ANDN U27736 ( .B(n27780), .A(n27781), .Z(n27777) );
  XOR U27737 ( .A(n27670), .B(n27782), .Z(n25253) );
  XNOR U27738 ( .A(n24221), .B(n27783), .Z(n27715) );
  XNOR U27739 ( .A(key[219]), .B(n25204), .Z(n27783) );
  XOR U27740 ( .A(n27784), .B(n27782), .Z(n25204) );
  XNOR U27741 ( .A(n27677), .B(n27678), .Z(n27782) );
  XOR U27742 ( .A(n27785), .B(n27786), .Z(n27678) );
  XNOR U27743 ( .A(n27787), .B(n27788), .Z(n27786) );
  NANDN U27744 ( .A(n27675), .B(n27789), .Z(n27788) );
  XOR U27745 ( .A(n27790), .B(n27791), .Z(n27677) );
  XOR U27746 ( .A(n27792), .B(n27793), .Z(n27791) );
  XOR U27747 ( .A(n27614), .B(n27611), .Z(n27784) );
  XNOR U27748 ( .A(n27640), .B(n27795), .Z(n27611) );
  XOR U27749 ( .A(n27796), .B(n27787), .Z(n27795) );
  OR U27750 ( .A(n27797), .B(n27798), .Z(n27787) );
  ANDN U27751 ( .B(n27799), .A(n27800), .Z(n27796) );
  XNOR U27752 ( .A(n27785), .B(n27801), .Z(n27614) );
  XNOR U27753 ( .A(n27645), .B(n27802), .Z(n27801) );
  NANDN U27754 ( .A(n27803), .B(n27804), .Z(n27802) );
  NANDN U27755 ( .A(n27805), .B(n27806), .Z(n27645) );
  XNOR U27756 ( .A(n27640), .B(n27807), .Z(n27785) );
  XNOR U27757 ( .A(n27808), .B(n27809), .Z(n27807) );
  NANDN U27758 ( .A(n27810), .B(n27811), .Z(n27809) );
  XOR U27759 ( .A(n27812), .B(n27808), .Z(n27640) );
  NANDN U27760 ( .A(n27813), .B(n27814), .Z(n27808) );
  ANDN U27761 ( .B(n27815), .A(n27816), .Z(n27812) );
  XNOR U27762 ( .A(n27615), .B(n25238), .Z(n24221) );
  XNOR U27763 ( .A(n25202), .B(n27702), .Z(n25238) );
  XOR U27764 ( .A(n27740), .B(n27817), .Z(n25202) );
  XOR U27765 ( .A(n27818), .B(n27819), .Z(n27565) );
  XNOR U27766 ( .A(n26081), .B(n24211), .Z(n27819) );
  IV U27767 ( .A(n27615), .Z(n24211) );
  XOR U27768 ( .A(n27817), .B(n27702), .Z(n27615) );
  XOR U27769 ( .A(n27703), .B(n27820), .Z(n27702) );
  XNOR U27770 ( .A(n27821), .B(n27822), .Z(n27820) );
  NOR U27771 ( .A(n27823), .B(n27739), .Z(n27821) );
  XNOR U27772 ( .A(n27824), .B(n27825), .Z(n27703) );
  XNOR U27773 ( .A(n27826), .B(n27827), .Z(n27825) );
  NANDN U27774 ( .A(n27828), .B(n27829), .Z(n27827) );
  XOR U27775 ( .A(n27604), .B(n27593), .Z(n26081) );
  XNOR U27776 ( .A(n27606), .B(n27607), .Z(n27593) );
  XOR U27777 ( .A(n27632), .B(n27830), .Z(n27607) );
  XNOR U27778 ( .A(n27831), .B(n27832), .Z(n27830) );
  OR U27779 ( .A(n27690), .B(n27833), .Z(n27832) );
  XNOR U27780 ( .A(n27685), .B(n27834), .Z(n27632) );
  XNOR U27781 ( .A(n27835), .B(n27836), .Z(n27834) );
  OR U27782 ( .A(n27728), .B(n27837), .Z(n27836) );
  XOR U27783 ( .A(n27724), .B(n27838), .Z(n27606) );
  XOR U27784 ( .A(n27722), .B(n27839), .Z(n27838) );
  OR U27785 ( .A(n27840), .B(n27696), .Z(n27839) );
  ANDN U27786 ( .B(n27698), .A(n27841), .Z(n27722) );
  XOR U27787 ( .A(n27637), .B(n27696), .Z(n27698) );
  IV U27788 ( .A(n27631), .Z(n27604) );
  XOR U27789 ( .A(n27719), .B(n27594), .Z(n27631) );
  XOR U27790 ( .A(n27685), .B(n27842), .Z(n27594) );
  XNOR U27791 ( .A(n27831), .B(n27843), .Z(n27842) );
  NANDN U27792 ( .A(n27844), .B(n27845), .Z(n27843) );
  OR U27793 ( .A(n27846), .B(n27847), .Z(n27831) );
  XOR U27794 ( .A(n27848), .B(n27835), .Z(n27685) );
  NANDN U27795 ( .A(n27849), .B(n27850), .Z(n27835) );
  AND U27796 ( .A(n27851), .B(n27852), .Z(n27848) );
  XNOR U27797 ( .A(n27724), .B(n27853), .Z(n27719) );
  XOR U27798 ( .A(n27854), .B(n27688), .Z(n27853) );
  OR U27799 ( .A(n27855), .B(n27846), .Z(n27688) );
  XOR U27800 ( .A(n27690), .B(n27856), .Z(n27846) );
  ANDN U27801 ( .B(n27857), .A(n27844), .Z(n27854) );
  XOR U27802 ( .A(n27858), .B(n27726), .Z(n27724) );
  OR U27803 ( .A(n27849), .B(n27859), .Z(n27726) );
  XOR U27804 ( .A(n27851), .B(n27728), .Z(n27849) );
  XOR U27805 ( .A(n27856), .B(n27696), .Z(n27728) );
  XNOR U27806 ( .A(n27860), .B(n27861), .Z(n27696) );
  NANDN U27807 ( .A(n27862), .B(n27863), .Z(n27861) );
  IV U27808 ( .A(n27844), .Z(n27856) );
  XNOR U27809 ( .A(n27864), .B(n27865), .Z(n27844) );
  NANDN U27810 ( .A(n27862), .B(n27866), .Z(n27865) );
  ANDN U27811 ( .B(n27851), .A(n27867), .Z(n27858) );
  XOR U27812 ( .A(n27637), .B(n27690), .Z(n27851) );
  XOR U27813 ( .A(n27868), .B(n27864), .Z(n27690) );
  NANDN U27814 ( .A(n27869), .B(n27870), .Z(n27864) );
  NANDN U27815 ( .A(n27869), .B(n27874), .Z(n27860) );
  XOR U27816 ( .A(n27875), .B(n27876), .Z(n27862) );
  XOR U27817 ( .A(n27877), .B(n27872), .Z(n27876) );
  XNOR U27818 ( .A(n27878), .B(n27879), .Z(n27875) );
  XNOR U27819 ( .A(n27880), .B(n27881), .Z(n27879) );
  ANDN U27820 ( .B(n27877), .A(n27872), .Z(n27880) );
  ANDN U27821 ( .B(n27877), .A(n27871), .Z(n27873) );
  XNOR U27822 ( .A(n27878), .B(n27882), .Z(n27871) );
  XOR U27823 ( .A(n27883), .B(n27881), .Z(n27882) );
  NAND U27824 ( .A(n27870), .B(n27874), .Z(n27881) );
  XNOR U27825 ( .A(n27866), .B(n27872), .Z(n27870) );
  XOR U27826 ( .A(n27884), .B(n27885), .Z(n27872) );
  XOR U27827 ( .A(n27886), .B(n27887), .Z(n27885) );
  XNOR U27828 ( .A(n27888), .B(n27889), .Z(n27884) );
  ANDN U27829 ( .B(n27890), .A(n27636), .Z(n27888) );
  AND U27830 ( .A(n27863), .B(n27866), .Z(n27883) );
  XNOR U27831 ( .A(n27863), .B(n27866), .Z(n27878) );
  XNOR U27832 ( .A(n27891), .B(n27892), .Z(n27866) );
  XNOR U27833 ( .A(n27893), .B(n27894), .Z(n27892) );
  XOR U27834 ( .A(n27886), .B(n27895), .Z(n27891) );
  XNOR U27835 ( .A(n27896), .B(n27889), .Z(n27895) );
  OR U27836 ( .A(n27697), .B(n27841), .Z(n27889) );
  XNOR U27837 ( .A(n27723), .B(n27840), .Z(n27841) );
  XNOR U27838 ( .A(n27636), .B(n27897), .Z(n27697) );
  NOR U27839 ( .A(n27897), .B(n27840), .Z(n27896) );
  XNOR U27840 ( .A(n27898), .B(n27899), .Z(n27863) );
  XNOR U27841 ( .A(n27900), .B(n27901), .Z(n27899) );
  XOR U27842 ( .A(n27833), .B(n27886), .Z(n27901) );
  XOR U27843 ( .A(n27890), .B(n27902), .Z(n27886) );
  XNOR U27844 ( .A(n27691), .B(n27903), .Z(n27898) );
  XNOR U27845 ( .A(n27904), .B(n27905), .Z(n27903) );
  ANDN U27846 ( .B(n27845), .A(n27906), .Z(n27904) );
  XNOR U27847 ( .A(n27907), .B(n27908), .Z(n27877) );
  XNOR U27848 ( .A(n27887), .B(n27909), .Z(n27908) );
  XNOR U27849 ( .A(n27845), .B(n27894), .Z(n27909) );
  XOR U27850 ( .A(n27840), .B(n27897), .Z(n27894) );
  XNOR U27851 ( .A(n27900), .B(n27910), .Z(n27887) );
  XNOR U27852 ( .A(n27911), .B(n27912), .Z(n27910) );
  NANDN U27853 ( .A(n27837), .B(n27729), .Z(n27912) );
  IV U27854 ( .A(n27893), .Z(n27900) );
  XNOR U27855 ( .A(n27913), .B(n27911), .Z(n27893) );
  NANDN U27856 ( .A(n27859), .B(n27850), .Z(n27911) );
  XOR U27857 ( .A(n27845), .B(n27897), .Z(n27837) );
  IV U27858 ( .A(n27695), .Z(n27897) );
  XOR U27859 ( .A(n27914), .B(n27915), .Z(n27695) );
  XNOR U27860 ( .A(n27916), .B(n27917), .Z(n27915) );
  XOR U27861 ( .A(n27867), .B(n27729), .Z(n27859) );
  XNOR U27862 ( .A(n27857), .B(n27840), .Z(n27729) );
  XNOR U27863 ( .A(n27917), .B(n27914), .Z(n27840) );
  ANDN U27864 ( .B(n27852), .A(n27867), .Z(n27913) );
  XNOR U27865 ( .A(n27918), .B(n27890), .Z(n27867) );
  IV U27866 ( .A(n27723), .Z(n27890) );
  XNOR U27867 ( .A(n27919), .B(n27920), .Z(n27723) );
  XNOR U27868 ( .A(n27921), .B(n27917), .Z(n27920) );
  XOR U27869 ( .A(n27922), .B(n27902), .Z(n27852) );
  XNOR U27870 ( .A(n27906), .B(n27923), .Z(n27907) );
  XNOR U27871 ( .A(n27924), .B(n27905), .Z(n27923) );
  OR U27872 ( .A(n27847), .B(n27855), .Z(n27905) );
  XOR U27873 ( .A(n27691), .B(n27857), .Z(n27855) );
  IV U27874 ( .A(n27906), .Z(n27857) );
  XOR U27875 ( .A(n27833), .B(n27845), .Z(n27847) );
  XNOR U27876 ( .A(n27902), .B(n27925), .Z(n27845) );
  XNOR U27877 ( .A(n27916), .B(n27919), .Z(n27925) );
  XNOR U27878 ( .A(msg[90]), .B(key[90]), .Z(n27919) );
  IV U27879 ( .A(n27636), .Z(n27902) );
  XOR U27880 ( .A(n27926), .B(n27927), .Z(n27636) );
  XOR U27881 ( .A(n27917), .B(n27928), .Z(n27927) );
  IV U27882 ( .A(n27922), .Z(n27833) );
  ANDN U27883 ( .B(n27922), .A(n27691), .Z(n27924) );
  XOR U27884 ( .A(n27914), .B(n27929), .Z(n27922) );
  XNOR U27885 ( .A(n27917), .B(n27930), .Z(n27929) );
  XOR U27886 ( .A(n27918), .B(n27931), .Z(n27917) );
  XNOR U27887 ( .A(msg[94]), .B(key[94]), .Z(n27931) );
  IV U27888 ( .A(n27926), .Z(n27914) );
  XOR U27889 ( .A(msg[93]), .B(key[93]), .Z(n27926) );
  XOR U27890 ( .A(n27932), .B(n27933), .Z(n27906) );
  XOR U27891 ( .A(n27930), .B(n27928), .Z(n27933) );
  XOR U27892 ( .A(msg[95]), .B(key[95]), .Z(n27928) );
  XNOR U27893 ( .A(msg[92]), .B(key[92]), .Z(n27930) );
  XOR U27894 ( .A(n27691), .B(n27921), .Z(n27932) );
  XNOR U27895 ( .A(n27916), .B(n27934), .Z(n27921) );
  XNOR U27896 ( .A(msg[91]), .B(key[91]), .Z(n27934) );
  XNOR U27897 ( .A(msg[89]), .B(key[89]), .Z(n27916) );
  IV U27898 ( .A(n27918), .Z(n27691) );
  XOR U27899 ( .A(msg[88]), .B(key[88]), .Z(n27918) );
  XOR U27900 ( .A(n24234), .B(n27935), .Z(n27818) );
  XOR U27901 ( .A(key[216]), .B(n27755), .Z(n27935) );
  IV U27902 ( .A(n25248), .Z(n27755) );
  XOR U27903 ( .A(n27629), .B(n27936), .Z(n25248) );
  XOR U27904 ( .A(n27740), .B(n27656), .Z(n27936) );
  XNOR U27905 ( .A(n27938), .B(n27939), .Z(n27937) );
  NANDN U27906 ( .A(n27707), .B(n27940), .Z(n27939) );
  XOR U27907 ( .A(n27709), .B(n27941), .Z(n27733) );
  XNOR U27908 ( .A(n27942), .B(n27943), .Z(n27941) );
  NANDN U27909 ( .A(n27828), .B(n27944), .Z(n27943) );
  IV U27910 ( .A(n27655), .Z(n27740) );
  XOR U27911 ( .A(n27824), .B(n27945), .Z(n27655) );
  XOR U27912 ( .A(n27822), .B(n27946), .Z(n27945) );
  NANDN U27913 ( .A(n27947), .B(n27948), .Z(n27946) );
  NOR U27914 ( .A(n27736), .B(n27949), .Z(n27822) );
  XOR U27915 ( .A(n27739), .B(n27948), .Z(n27736) );
  XOR U27916 ( .A(n27817), .B(n27732), .Z(n27629) );
  XNOR U27917 ( .A(n27709), .B(n27950), .Z(n27732) );
  XNOR U27918 ( .A(n27938), .B(n27951), .Z(n27950) );
  OR U27919 ( .A(n27952), .B(n27953), .Z(n27951) );
  OR U27920 ( .A(n27954), .B(n27955), .Z(n27938) );
  XNOR U27921 ( .A(n27956), .B(n27942), .Z(n27709) );
  NANDN U27922 ( .A(n27957), .B(n27958), .Z(n27942) );
  AND U27923 ( .A(n27959), .B(n27960), .Z(n27956) );
  XOR U27924 ( .A(n27824), .B(n27961), .Z(n27817) );
  XOR U27925 ( .A(n27962), .B(n27705), .Z(n27961) );
  OR U27926 ( .A(n27963), .B(n27954), .Z(n27705) );
  XNOR U27927 ( .A(n27707), .B(n27952), .Z(n27954) );
  NOR U27928 ( .A(n27964), .B(n27952), .Z(n27962) );
  XOR U27929 ( .A(n27965), .B(n27826), .Z(n27824) );
  OR U27930 ( .A(n27957), .B(n27966), .Z(n27826) );
  XOR U27931 ( .A(n27952), .B(n27948), .Z(n27828) );
  IV U27932 ( .A(n27714), .Z(n27948) );
  XNOR U27933 ( .A(n27967), .B(n27968), .Z(n27714) );
  NANDN U27934 ( .A(n27969), .B(n27970), .Z(n27968) );
  XNOR U27935 ( .A(n27971), .B(n27972), .Z(n27952) );
  NANDN U27936 ( .A(n27969), .B(n27973), .Z(n27972) );
  ANDN U27937 ( .B(n27959), .A(n27974), .Z(n27965) );
  XOR U27938 ( .A(n27707), .B(n27739), .Z(n27959) );
  XOR U27939 ( .A(n27975), .B(n27967), .Z(n27739) );
  NANDN U27940 ( .A(n27976), .B(n27977), .Z(n27967) );
  XOR U27941 ( .A(n27970), .B(n27978), .Z(n27977) );
  ANDN U27942 ( .B(n27978), .A(n27979), .Z(n27975) );
  NANDN U27943 ( .A(n27976), .B(n27981), .Z(n27971) );
  XOR U27944 ( .A(n27982), .B(n27983), .Z(n27969) );
  XOR U27945 ( .A(n27984), .B(n27985), .Z(n27983) );
  XNOR U27946 ( .A(n27986), .B(n27987), .Z(n27982) );
  XNOR U27947 ( .A(n27988), .B(n27989), .Z(n27987) );
  ANDN U27948 ( .B(n27985), .A(n27984), .Z(n27988) );
  ANDN U27949 ( .B(n27985), .A(n27979), .Z(n27980) );
  XNOR U27950 ( .A(n27986), .B(n27990), .Z(n27979) );
  XOR U27951 ( .A(n27991), .B(n27989), .Z(n27990) );
  NAND U27952 ( .A(n27981), .B(n27992), .Z(n27989) );
  XNOR U27953 ( .A(n27970), .B(n27984), .Z(n27992) );
  IV U27954 ( .A(n27978), .Z(n27984) );
  XNOR U27955 ( .A(n27993), .B(n27994), .Z(n27978) );
  XNOR U27956 ( .A(n27995), .B(n27996), .Z(n27994) );
  XOR U27957 ( .A(n27953), .B(n27997), .Z(n27996) );
  XNOR U27958 ( .A(n27964), .B(n27998), .Z(n27993) );
  XNOR U27959 ( .A(n27999), .B(n28000), .Z(n27998) );
  AND U27960 ( .A(n27940), .B(n27708), .Z(n27999) );
  XOR U27961 ( .A(n27973), .B(n27985), .Z(n27981) );
  AND U27962 ( .A(n27970), .B(n27973), .Z(n27991) );
  XNOR U27963 ( .A(n27970), .B(n27973), .Z(n27986) );
  XNOR U27964 ( .A(n28001), .B(n28002), .Z(n27973) );
  XNOR U27965 ( .A(n28003), .B(n27997), .Z(n28002) );
  XOR U27966 ( .A(n28004), .B(n28005), .Z(n28001) );
  XNOR U27967 ( .A(n28006), .B(n28007), .Z(n28005) );
  ANDN U27968 ( .B(n27713), .A(n27947), .Z(n28006) );
  XNOR U27969 ( .A(n28008), .B(n28009), .Z(n27970) );
  XNOR U27970 ( .A(n27940), .B(n28004), .Z(n28010) );
  XOR U27971 ( .A(n27708), .B(n28011), .Z(n28008) );
  XNOR U27972 ( .A(n28012), .B(n28000), .Z(n28011) );
  OR U27973 ( .A(n27955), .B(n27963), .Z(n28000) );
  XOR U27974 ( .A(n27708), .B(n27964), .Z(n27963) );
  XNOR U27975 ( .A(n27940), .B(n28013), .Z(n27955) );
  ANDN U27976 ( .B(n28014), .A(n27953), .Z(n28012) );
  XNOR U27977 ( .A(n28015), .B(n28016), .Z(n27985) );
  XOR U27978 ( .A(n28003), .B(n27995), .Z(n28016) );
  XOR U27979 ( .A(n28004), .B(n28017), .Z(n27995) );
  XNOR U27980 ( .A(n28018), .B(n28019), .Z(n28017) );
  NAND U27981 ( .A(n27829), .B(n27944), .Z(n28019) );
  XNOR U27982 ( .A(n28020), .B(n28018), .Z(n28004) );
  NANDN U27983 ( .A(n27966), .B(n27958), .Z(n28018) );
  XOR U27984 ( .A(n27960), .B(n27944), .Z(n27958) );
  XOR U27985 ( .A(n28013), .B(n27713), .Z(n27944) );
  IV U27986 ( .A(n27953), .Z(n28013) );
  XOR U27987 ( .A(n27738), .B(n28021), .Z(n27953) );
  XNOR U27988 ( .A(n28022), .B(n28023), .Z(n28021) );
  XOR U27989 ( .A(n27974), .B(n27829), .Z(n27966) );
  XNOR U27990 ( .A(n28014), .B(n27947), .Z(n27829) );
  IV U27991 ( .A(n27964), .Z(n28014) );
  XOR U27992 ( .A(n28024), .B(n28025), .Z(n27964) );
  XOR U27993 ( .A(n28026), .B(n28027), .Z(n28025) );
  XNOR U27994 ( .A(n27708), .B(n28028), .Z(n28024) );
  ANDN U27995 ( .B(n27960), .A(n27974), .Z(n28020) );
  XNOR U27996 ( .A(n27708), .B(n28029), .Z(n27974) );
  XOR U27997 ( .A(n27940), .B(n27738), .Z(n27960) );
  XOR U27998 ( .A(n28030), .B(n28031), .Z(n27940) );
  XOR U27999 ( .A(n28032), .B(n28027), .Z(n28031) );
  XOR U28000 ( .A(msg[52]), .B(key[52]), .Z(n28027) );
  XOR U28001 ( .A(n28029), .B(n27738), .Z(n28003) );
  IV U28002 ( .A(n27823), .Z(n28029) );
  XNOR U28003 ( .A(n28033), .B(n28007), .Z(n28015) );
  OR U28004 ( .A(n27737), .B(n27949), .Z(n28007) );
  XNOR U28005 ( .A(n27823), .B(n27947), .Z(n27949) );
  XOR U28006 ( .A(n28034), .B(n28030), .Z(n27947) );
  XNOR U28007 ( .A(n27738), .B(n27713), .Z(n27737) );
  XOR U28008 ( .A(n28030), .B(n28035), .Z(n27713) );
  XOR U28009 ( .A(n28022), .B(n28034), .Z(n28035) );
  ANDN U28010 ( .B(n27738), .A(n27823), .Z(n28033) );
  XNOR U28011 ( .A(n28023), .B(n28036), .Z(n27823) );
  XOR U28012 ( .A(n28028), .B(n28034), .Z(n28036) );
  IV U28013 ( .A(n28032), .Z(n28034) );
  XNOR U28014 ( .A(n28022), .B(n28037), .Z(n28028) );
  XNOR U28015 ( .A(msg[51]), .B(key[51]), .Z(n28037) );
  XNOR U28016 ( .A(msg[49]), .B(key[49]), .Z(n28022) );
  XNOR U28017 ( .A(msg[50]), .B(key[50]), .Z(n28023) );
  XOR U28018 ( .A(n28030), .B(n28038), .Z(n27738) );
  XNOR U28019 ( .A(n28032), .B(n28026), .Z(n28038) );
  XNOR U28020 ( .A(msg[55]), .B(key[55]), .Z(n28026) );
  XOR U28021 ( .A(n27708), .B(n28039), .Z(n28032) );
  XNOR U28022 ( .A(msg[54]), .B(key[54]), .Z(n28039) );
  XOR U28023 ( .A(msg[48]), .B(key[48]), .Z(n27708) );
  XNOR U28024 ( .A(msg[53]), .B(key[53]), .Z(n28030) );
  XOR U28025 ( .A(n26056), .B(n25215), .Z(n24234) );
  IV U28026 ( .A(n26082), .Z(n25215) );
  XNOR U28027 ( .A(n27659), .B(n28040), .Z(n27620) );
  XNOR U28028 ( .A(n27768), .B(n28041), .Z(n28040) );
  NANDN U28029 ( .A(n28042), .B(n27749), .Z(n28041) );
  NANDN U28030 ( .A(n28043), .B(n27748), .Z(n27768) );
  XOR U28031 ( .A(n27749), .B(n27626), .Z(n27748) );
  XNOR U28032 ( .A(n27766), .B(n28044), .Z(n27659) );
  XNOR U28033 ( .A(n28045), .B(n28046), .Z(n28044) );
  NAND U28034 ( .A(n27765), .B(n28047), .Z(n28046) );
  XNOR U28035 ( .A(n27766), .B(n28048), .Z(n27682) );
  XOR U28036 ( .A(n28049), .B(n27661), .Z(n28048) );
  OR U28037 ( .A(n28050), .B(n27775), .Z(n27661) );
  XNOR U28038 ( .A(n27663), .B(n27773), .Z(n27775) );
  NOR U28039 ( .A(n28051), .B(n27773), .Z(n28049) );
  XOR U28040 ( .A(n28052), .B(n28045), .Z(n27766) );
  OR U28041 ( .A(n27778), .B(n28053), .Z(n28045) );
  XNOR U28042 ( .A(n28054), .B(n27765), .Z(n27778) );
  XNOR U28043 ( .A(n27773), .B(n27626), .Z(n27765) );
  XOR U28044 ( .A(n28055), .B(n28056), .Z(n27626) );
  NAND U28045 ( .A(n28057), .B(n28058), .Z(n28056) );
  XNOR U28046 ( .A(n28059), .B(n28060), .Z(n27773) );
  NANDN U28047 ( .A(n28061), .B(n28057), .Z(n28060) );
  ANDN U28048 ( .B(n28054), .A(n28062), .Z(n28052) );
  IV U28049 ( .A(n27781), .Z(n28054) );
  XOR U28050 ( .A(n27663), .B(n27749), .Z(n27781) );
  XOR U28051 ( .A(n28055), .B(n28063), .Z(n27749) );
  NANDN U28052 ( .A(n28064), .B(n28065), .Z(n28063) );
  NAND U28053 ( .A(n28066), .B(n28067), .Z(n28055) );
  NANDN U28054 ( .A(n28069), .B(n28067), .Z(n28059) );
  XNOR U28055 ( .A(n28064), .B(n28057), .Z(n28067) );
  XNOR U28056 ( .A(n28070), .B(n28071), .Z(n28057) );
  XOR U28057 ( .A(n28072), .B(n28065), .Z(n28071) );
  IV U28058 ( .A(n28073), .Z(n28065) );
  XNOR U28059 ( .A(n28074), .B(n28075), .Z(n28070) );
  XNOR U28060 ( .A(n28076), .B(n28077), .Z(n28075) );
  NOR U28061 ( .A(n28073), .B(n28074), .Z(n28076) );
  NOR U28062 ( .A(n28064), .B(n28074), .Z(n28068) );
  XNOR U28063 ( .A(n28072), .B(n28078), .Z(n28064) );
  XNOR U28064 ( .A(n28077), .B(n28079), .Z(n28078) );
  NANDN U28065 ( .A(n28061), .B(n28058), .Z(n28079) );
  NANDN U28066 ( .A(n28069), .B(n28066), .Z(n28077) );
  XNOR U28067 ( .A(n28058), .B(n28073), .Z(n28066) );
  XOR U28068 ( .A(n28080), .B(n28081), .Z(n28073) );
  XOR U28069 ( .A(n28082), .B(n28083), .Z(n28081) );
  XOR U28070 ( .A(n27774), .B(n28084), .Z(n28083) );
  XNOR U28071 ( .A(n28051), .B(n28085), .Z(n28080) );
  XNOR U28072 ( .A(n28086), .B(n28087), .Z(n28085) );
  AND U28073 ( .A(n27664), .B(n27760), .Z(n28086) );
  XOR U28074 ( .A(n28088), .B(n28089), .Z(n28074) );
  XNOR U28075 ( .A(n28090), .B(n28084), .Z(n28089) );
  XNOR U28076 ( .A(n28091), .B(n28092), .Z(n28084) );
  XNOR U28077 ( .A(n28093), .B(n28094), .Z(n28092) );
  NAND U28078 ( .A(n28047), .B(n27764), .Z(n28094) );
  XNOR U28079 ( .A(n28095), .B(n28096), .Z(n28088) );
  ANDN U28080 ( .B(n28097), .A(n27750), .Z(n28095) );
  XOR U28081 ( .A(n28061), .B(n28058), .Z(n28072) );
  XNOR U28082 ( .A(n28098), .B(n28099), .Z(n28058) );
  XOR U28083 ( .A(n28100), .B(n28101), .Z(n28099) );
  XOR U28084 ( .A(n28090), .B(n27760), .Z(n28101) );
  XOR U28085 ( .A(n27664), .B(n28102), .Z(n28098) );
  XNOR U28086 ( .A(n28103), .B(n28087), .Z(n28102) );
  OR U28087 ( .A(n27776), .B(n28050), .Z(n28087) );
  XNOR U28088 ( .A(n27664), .B(n28104), .Z(n28050) );
  XNOR U28089 ( .A(n27760), .B(n27774), .Z(n27776) );
  ANDN U28090 ( .B(n27774), .A(n28051), .Z(n28103) );
  XOR U28091 ( .A(n28105), .B(n28106), .Z(n28061) );
  XOR U28092 ( .A(n28091), .B(n28082), .Z(n28106) );
  XOR U28093 ( .A(n28107), .B(n28108), .Z(n28082) );
  IV U28094 ( .A(n28100), .Z(n28091) );
  XNOR U28095 ( .A(n28109), .B(n28093), .Z(n28100) );
  NANDN U28096 ( .A(n28053), .B(n27779), .Z(n28093) );
  XOR U28097 ( .A(n27780), .B(n27764), .Z(n27779) );
  XOR U28098 ( .A(n28108), .B(n27774), .Z(n27764) );
  XNOR U28099 ( .A(n28110), .B(n28111), .Z(n27774) );
  XNOR U28100 ( .A(n28112), .B(n28113), .Z(n28111) );
  IV U28101 ( .A(n27627), .Z(n28108) );
  XOR U28102 ( .A(n28062), .B(n28047), .Z(n28053) );
  XNOR U28103 ( .A(n28104), .B(n27770), .Z(n28047) );
  IV U28104 ( .A(n28051), .Z(n28104) );
  XOR U28105 ( .A(n28114), .B(n28115), .Z(n28051) );
  XOR U28106 ( .A(n28116), .B(n28117), .Z(n28115) );
  XNOR U28107 ( .A(n27664), .B(n28118), .Z(n28114) );
  ANDN U28108 ( .B(n27780), .A(n28062), .Z(n28109) );
  XNOR U28109 ( .A(n27664), .B(n28097), .Z(n28062) );
  XOR U28110 ( .A(n28110), .B(n27760), .Z(n27780) );
  XNOR U28111 ( .A(n28119), .B(n28120), .Z(n27760) );
  XOR U28112 ( .A(n28121), .B(n28117), .Z(n28120) );
  XOR U28113 ( .A(msg[12]), .B(key[12]), .Z(n28117) );
  IV U28114 ( .A(n27750), .Z(n28110) );
  XNOR U28115 ( .A(n28090), .B(n28122), .Z(n28105) );
  XNOR U28116 ( .A(n28123), .B(n28096), .Z(n28122) );
  OR U28117 ( .A(n27747), .B(n28043), .Z(n28096) );
  XNOR U28118 ( .A(n28042), .B(n27770), .Z(n28043) );
  IV U28119 ( .A(n28107), .Z(n27770) );
  XNOR U28120 ( .A(n27750), .B(n27627), .Z(n27747) );
  ANDN U28121 ( .B(n28107), .A(n27627), .Z(n28123) );
  XOR U28122 ( .A(n28119), .B(n28124), .Z(n27627) );
  XOR U28123 ( .A(n28113), .B(n28125), .Z(n28124) );
  XOR U28124 ( .A(n28097), .B(n27750), .Z(n28090) );
  XOR U28125 ( .A(n28119), .B(n28126), .Z(n27750) );
  XNOR U28126 ( .A(n28121), .B(n28116), .Z(n28126) );
  XNOR U28127 ( .A(msg[15]), .B(key[15]), .Z(n28116) );
  XOR U28128 ( .A(msg[13]), .B(key[13]), .Z(n28119) );
  IV U28129 ( .A(n28042), .Z(n28097) );
  XOR U28130 ( .A(n28125), .B(n28127), .Z(n28042) );
  XNOR U28131 ( .A(n28112), .B(n28118), .Z(n28127) );
  XNOR U28132 ( .A(n28113), .B(n28128), .Z(n28118) );
  XNOR U28133 ( .A(msg[11]), .B(key[11]), .Z(n28128) );
  XNOR U28134 ( .A(msg[9]), .B(key[9]), .Z(n28113) );
  XNOR U28135 ( .A(msg[10]), .B(key[10]), .Z(n28112) );
  IV U28136 ( .A(n28121), .Z(n28125) );
  XOR U28137 ( .A(n27664), .B(n28129), .Z(n28121) );
  XNOR U28138 ( .A(msg[14]), .B(key[14]), .Z(n28129) );
  XOR U28139 ( .A(msg[8]), .B(key[8]), .Z(n27664) );
  XOR U28140 ( .A(n27613), .B(n27642), .Z(n26056) );
  XNOR U28141 ( .A(n27671), .B(n28130), .Z(n27642) );
  XNOR U28142 ( .A(n28131), .B(n27792), .Z(n28130) );
  ANDN U28143 ( .B(n27806), .A(n28132), .Z(n27792) );
  XOR U28144 ( .A(n27803), .B(n27647), .Z(n27806) );
  NOR U28145 ( .A(n28133), .B(n27803), .Z(n28131) );
  XNOR U28146 ( .A(n27790), .B(n28134), .Z(n27671) );
  XNOR U28147 ( .A(n28135), .B(n28136), .Z(n28134) );
  NANDN U28148 ( .A(n27810), .B(n28137), .Z(n28136) );
  XNOR U28149 ( .A(n27790), .B(n28138), .Z(n27613) );
  XOR U28150 ( .A(n28139), .B(n27673), .Z(n28138) );
  OR U28151 ( .A(n28140), .B(n27797), .Z(n27673) );
  XOR U28152 ( .A(n27675), .B(n28141), .Z(n27797) );
  ANDN U28153 ( .B(n28142), .A(n27800), .Z(n28139) );
  IV U28154 ( .A(n28141), .Z(n27800) );
  XOR U28155 ( .A(n28143), .B(n28135), .Z(n27790) );
  OR U28156 ( .A(n27813), .B(n28144), .Z(n28135) );
  XOR U28157 ( .A(n28145), .B(n27810), .Z(n27813) );
  XOR U28158 ( .A(n28141), .B(n27647), .Z(n27810) );
  XNOR U28159 ( .A(n28146), .B(n28147), .Z(n27647) );
  NANDN U28160 ( .A(n28148), .B(n28149), .Z(n28147) );
  XOR U28161 ( .A(n28150), .B(n28151), .Z(n28141) );
  NANDN U28162 ( .A(n28148), .B(n28152), .Z(n28151) );
  ANDN U28163 ( .B(n28145), .A(n28153), .Z(n28143) );
  IV U28164 ( .A(n27816), .Z(n28145) );
  XNOR U28165 ( .A(n27675), .B(n27803), .Z(n27816) );
  XOR U28166 ( .A(n28154), .B(n28146), .Z(n27803) );
  NANDN U28167 ( .A(n28155), .B(n28156), .Z(n28146) );
  XOR U28168 ( .A(n28149), .B(n28157), .Z(n28156) );
  ANDN U28169 ( .B(n28157), .A(n28158), .Z(n28154) );
  NANDN U28170 ( .A(n28155), .B(n28160), .Z(n28150) );
  XOR U28171 ( .A(n28161), .B(n28162), .Z(n28148) );
  XOR U28172 ( .A(n28163), .B(n28164), .Z(n28162) );
  XNOR U28173 ( .A(n28165), .B(n28166), .Z(n28161) );
  XNOR U28174 ( .A(n28167), .B(n28168), .Z(n28166) );
  ANDN U28175 ( .B(n28164), .A(n28163), .Z(n28167) );
  ANDN U28176 ( .B(n28164), .A(n28158), .Z(n28159) );
  XNOR U28177 ( .A(n28165), .B(n28169), .Z(n28158) );
  XOR U28178 ( .A(n28170), .B(n28168), .Z(n28169) );
  NAND U28179 ( .A(n28160), .B(n28171), .Z(n28168) );
  XNOR U28180 ( .A(n28149), .B(n28163), .Z(n28171) );
  IV U28181 ( .A(n28157), .Z(n28163) );
  XNOR U28182 ( .A(n28172), .B(n28173), .Z(n28157) );
  XNOR U28183 ( .A(n28174), .B(n28175), .Z(n28173) );
  XOR U28184 ( .A(n28176), .B(n28177), .Z(n28175) );
  XNOR U28185 ( .A(n28178), .B(n28179), .Z(n28172) );
  XNOR U28186 ( .A(n28180), .B(n28181), .Z(n28179) );
  AND U28187 ( .A(n27789), .B(n27676), .Z(n28180) );
  XOR U28188 ( .A(n28152), .B(n28164), .Z(n28160) );
  AND U28189 ( .A(n28149), .B(n28152), .Z(n28170) );
  XNOR U28190 ( .A(n28149), .B(n28152), .Z(n28165) );
  XNOR U28191 ( .A(n28182), .B(n28183), .Z(n28152) );
  XNOR U28192 ( .A(n28184), .B(n28177), .Z(n28183) );
  XOR U28193 ( .A(n28185), .B(n28186), .Z(n28182) );
  XNOR U28194 ( .A(n28187), .B(n28188), .Z(n28186) );
  ANDN U28195 ( .B(n27646), .A(n27794), .Z(n28187) );
  XNOR U28196 ( .A(n28189), .B(n28190), .Z(n28149) );
  XNOR U28197 ( .A(n27789), .B(n28185), .Z(n28191) );
  XOR U28198 ( .A(n27676), .B(n28192), .Z(n28189) );
  XNOR U28199 ( .A(n28193), .B(n28181), .Z(n28192) );
  OR U28200 ( .A(n27798), .B(n28140), .Z(n28181) );
  XOR U28201 ( .A(n27676), .B(n28178), .Z(n28140) );
  XNOR U28202 ( .A(n27789), .B(n27799), .Z(n27798) );
  ANDN U28203 ( .B(n28142), .A(n28176), .Z(n28193) );
  XNOR U28204 ( .A(n28194), .B(n28195), .Z(n28164) );
  XOR U28205 ( .A(n28184), .B(n28174), .Z(n28195) );
  XOR U28206 ( .A(n28185), .B(n28196), .Z(n28174) );
  XNOR U28207 ( .A(n28197), .B(n28198), .Z(n28196) );
  NAND U28208 ( .A(n28137), .B(n27811), .Z(n28198) );
  XNOR U28209 ( .A(n28199), .B(n28197), .Z(n28185) );
  NANDN U28210 ( .A(n28144), .B(n27814), .Z(n28197) );
  XOR U28211 ( .A(n27815), .B(n27811), .Z(n27814) );
  XOR U28212 ( .A(n27799), .B(n27646), .Z(n27811) );
  IV U28213 ( .A(n28176), .Z(n27799) );
  XOR U28214 ( .A(n27804), .B(n28200), .Z(n28176) );
  XNOR U28215 ( .A(n28201), .B(n28202), .Z(n28200) );
  XOR U28216 ( .A(n28153), .B(n28137), .Z(n28144) );
  XNOR U28217 ( .A(n28142), .B(n27794), .Z(n28137) );
  IV U28218 ( .A(n28178), .Z(n28142) );
  XOR U28219 ( .A(n28203), .B(n28204), .Z(n28178) );
  XOR U28220 ( .A(n28205), .B(n28206), .Z(n28204) );
  XOR U28221 ( .A(n27676), .B(n28207), .Z(n28203) );
  ANDN U28222 ( .B(n27815), .A(n28153), .Z(n28199) );
  XOR U28223 ( .A(n27676), .B(n28133), .Z(n28153) );
  XOR U28224 ( .A(n27789), .B(n27804), .Z(n27815) );
  XOR U28225 ( .A(n28208), .B(n28209), .Z(n27789) );
  XOR U28226 ( .A(n28210), .B(n28206), .Z(n28209) );
  XOR U28227 ( .A(msg[100]), .B(key[100]), .Z(n28206) );
  XNOR U28228 ( .A(n28133), .B(n27804), .Z(n28184) );
  XNOR U28229 ( .A(n28211), .B(n28188), .Z(n28194) );
  OR U28230 ( .A(n27805), .B(n28132), .Z(n28188) );
  XNOR U28231 ( .A(n28133), .B(n27794), .Z(n28132) );
  XOR U28232 ( .A(n28212), .B(n28208), .Z(n27794) );
  XNOR U28233 ( .A(n27804), .B(n27646), .Z(n27805) );
  XOR U28234 ( .A(n28208), .B(n28213), .Z(n27646) );
  XOR U28235 ( .A(n28202), .B(n28212), .Z(n28213) );
  ANDN U28236 ( .B(n27804), .A(n28133), .Z(n28211) );
  XOR U28237 ( .A(n28212), .B(n28214), .Z(n28133) );
  XOR U28238 ( .A(n28201), .B(n28207), .Z(n28214) );
  XOR U28239 ( .A(n28202), .B(n28215), .Z(n28207) );
  XNOR U28240 ( .A(msg[99]), .B(key[99]), .Z(n28215) );
  XNOR U28241 ( .A(msg[97]), .B(key[97]), .Z(n28202) );
  XNOR U28242 ( .A(msg[98]), .B(key[98]), .Z(n28201) );
  IV U28243 ( .A(n28210), .Z(n28212) );
  XOR U28244 ( .A(n28208), .B(n28216), .Z(n27804) );
  XNOR U28245 ( .A(n28210), .B(n28205), .Z(n28216) );
  XNOR U28246 ( .A(msg[103]), .B(key[103]), .Z(n28205) );
  XOR U28247 ( .A(n27676), .B(n28217), .Z(n28210) );
  XNOR U28248 ( .A(msg[102]), .B(key[102]), .Z(n28217) );
  XOR U28249 ( .A(msg[96]), .B(key[96]), .Z(n27676) );
  XNOR U28250 ( .A(msg[101]), .B(key[101]), .Z(n28208) );
  XNOR U28251 ( .A(n26709), .B(n28218), .Z(n23036) );
  XOR U28252 ( .A(n26634), .B(n26635), .Z(n28218) );
  XOR U28253 ( .A(n28219), .B(n28220), .Z(n26635) );
  XOR U28254 ( .A(n28221), .B(n28222), .Z(n28220) );
  NAND U28255 ( .A(n28223), .B(n26662), .Z(n28222) );
  XNOR U28256 ( .A(n26607), .B(n26608), .Z(n26634) );
  XNOR U28257 ( .A(n26651), .B(n28224), .Z(n26608) );
  XOR U28258 ( .A(n28225), .B(n28226), .Z(n28224) );
  AND U28259 ( .A(n28227), .B(n28228), .Z(n28225) );
  IV U28260 ( .A(n26632), .Z(n26709) );
  XOR U28261 ( .A(n26710), .B(n28229), .Z(n26632) );
  XNOR U28262 ( .A(n28226), .B(n28230), .Z(n28229) );
  NANDN U28263 ( .A(n26656), .B(n28231), .Z(n28230) );
  OR U28264 ( .A(n28232), .B(n28233), .Z(n28226) );
  XNOR U28265 ( .A(n26651), .B(n28234), .Z(n26710) );
  XNOR U28266 ( .A(n28235), .B(n28236), .Z(n28234) );
  NAND U28267 ( .A(n28237), .B(n28238), .Z(n28236) );
  XOR U28268 ( .A(n28239), .B(n28235), .Z(n26651) );
  NANDN U28269 ( .A(n28240), .B(n28241), .Z(n28235) );
  ANDN U28270 ( .B(n28242), .A(n28243), .Z(n28239) );
  XNOR U28271 ( .A(n22239), .B(n28244), .Z(n26785) );
  XOR U28272 ( .A(key[328]), .B(n26646), .Z(n28244) );
  XOR U28273 ( .A(n26607), .B(n26658), .Z(n26646) );
  XNOR U28274 ( .A(n26652), .B(n28245), .Z(n26658) );
  XNOR U28275 ( .A(n28246), .B(n28221), .Z(n28245) );
  ANDN U28276 ( .B(n26716), .A(n28247), .Z(n28221) );
  XNOR U28277 ( .A(n26713), .B(n26662), .Z(n26716) );
  NOR U28278 ( .A(n28248), .B(n26713), .Z(n28246) );
  XNOR U28279 ( .A(n28219), .B(n28249), .Z(n26652) );
  XNOR U28280 ( .A(n28250), .B(n28251), .Z(n28249) );
  NAND U28281 ( .A(n28238), .B(n28252), .Z(n28251) );
  XNOR U28282 ( .A(n28219), .B(n28253), .Z(n26607) );
  XOR U28283 ( .A(n28254), .B(n26654), .Z(n28253) );
  OR U28284 ( .A(n28255), .B(n28232), .Z(n26654) );
  XOR U28285 ( .A(n26656), .B(n28228), .Z(n28232) );
  ANDN U28286 ( .B(n28228), .A(n28256), .Z(n28254) );
  XOR U28287 ( .A(n28257), .B(n28250), .Z(n28219) );
  OR U28288 ( .A(n28258), .B(n28240), .Z(n28250) );
  XOR U28289 ( .A(n28243), .B(n28238), .Z(n28240) );
  XOR U28290 ( .A(n28228), .B(n26662), .Z(n28238) );
  XOR U28291 ( .A(n28259), .B(n28260), .Z(n26662) );
  NANDN U28292 ( .A(n28261), .B(n28262), .Z(n28260) );
  XOR U28293 ( .A(n28263), .B(n28264), .Z(n28228) );
  OR U28294 ( .A(n28261), .B(n28265), .Z(n28264) );
  IV U28295 ( .A(n28266), .Z(n28243) );
  ANDN U28296 ( .B(n28266), .A(n28267), .Z(n28257) );
  XOR U28297 ( .A(n26656), .B(n26713), .Z(n28266) );
  XOR U28298 ( .A(n28268), .B(n28259), .Z(n26713) );
  NANDN U28299 ( .A(n28269), .B(n28270), .Z(n28259) );
  ANDN U28300 ( .B(n28271), .A(n28272), .Z(n28268) );
  NANDN U28301 ( .A(n28269), .B(n28274), .Z(n28263) );
  XOR U28302 ( .A(n28275), .B(n28261), .Z(n28269) );
  XNOR U28303 ( .A(n28276), .B(n28277), .Z(n28261) );
  XOR U28304 ( .A(n28278), .B(n28271), .Z(n28277) );
  XNOR U28305 ( .A(n28279), .B(n28280), .Z(n28276) );
  XNOR U28306 ( .A(n28281), .B(n28282), .Z(n28280) );
  ANDN U28307 ( .B(n28271), .A(n28283), .Z(n28281) );
  IV U28308 ( .A(n28284), .Z(n28271) );
  ANDN U28309 ( .B(n28275), .A(n28283), .Z(n28273) );
  IV U28310 ( .A(n28279), .Z(n28283) );
  IV U28311 ( .A(n28272), .Z(n28275) );
  XNOR U28312 ( .A(n28278), .B(n28285), .Z(n28272) );
  XOR U28313 ( .A(n28286), .B(n28282), .Z(n28285) );
  NAND U28314 ( .A(n28274), .B(n28270), .Z(n28282) );
  XNOR U28315 ( .A(n28262), .B(n28284), .Z(n28270) );
  XOR U28316 ( .A(n28287), .B(n28288), .Z(n28284) );
  XOR U28317 ( .A(n28289), .B(n28290), .Z(n28288) );
  XNOR U28318 ( .A(n28227), .B(n28291), .Z(n28290) );
  XNOR U28319 ( .A(n28292), .B(n28293), .Z(n28287) );
  XNOR U28320 ( .A(n28294), .B(n28295), .Z(n28293) );
  ANDN U28321 ( .B(n28231), .A(n26657), .Z(n28294) );
  XNOR U28322 ( .A(n28279), .B(n28265), .Z(n28274) );
  XOR U28323 ( .A(n28296), .B(n28297), .Z(n28279) );
  XNOR U28324 ( .A(n28298), .B(n28291), .Z(n28297) );
  XOR U28325 ( .A(n28299), .B(n28300), .Z(n28291) );
  XNOR U28326 ( .A(n28301), .B(n28302), .Z(n28300) );
  NAND U28327 ( .A(n28252), .B(n28237), .Z(n28302) );
  XNOR U28328 ( .A(n28303), .B(n28304), .Z(n28296) );
  ANDN U28329 ( .B(n28305), .A(n28248), .Z(n28303) );
  ANDN U28330 ( .B(n28262), .A(n28265), .Z(n28286) );
  XOR U28331 ( .A(n28265), .B(n28262), .Z(n28278) );
  XNOR U28332 ( .A(n28306), .B(n28307), .Z(n28262) );
  XNOR U28333 ( .A(n28299), .B(n28308), .Z(n28307) );
  XNOR U28334 ( .A(n28298), .B(n28231), .Z(n28308) );
  XNOR U28335 ( .A(n28309), .B(n28310), .Z(n28306) );
  XNOR U28336 ( .A(n28311), .B(n28295), .Z(n28310) );
  OR U28337 ( .A(n28233), .B(n28255), .Z(n28295) );
  XNOR U28338 ( .A(n28309), .B(n28292), .Z(n28255) );
  XNOR U28339 ( .A(n28231), .B(n28227), .Z(n28233) );
  ANDN U28340 ( .B(n28227), .A(n28256), .Z(n28311) );
  XOR U28341 ( .A(n28312), .B(n28313), .Z(n28265) );
  XOR U28342 ( .A(n28299), .B(n28289), .Z(n28313) );
  XOR U28343 ( .A(n28223), .B(n26663), .Z(n28289) );
  XOR U28344 ( .A(n28314), .B(n28301), .Z(n28299) );
  NANDN U28345 ( .A(n28258), .B(n28241), .Z(n28301) );
  XOR U28346 ( .A(n28242), .B(n28237), .Z(n28241) );
  XNOR U28347 ( .A(n28305), .B(n28315), .Z(n28227) );
  XOR U28348 ( .A(n28316), .B(n28317), .Z(n28315) );
  XOR U28349 ( .A(n28267), .B(n28252), .Z(n28258) );
  XNOR U28350 ( .A(n28256), .B(n28223), .Z(n28252) );
  IV U28351 ( .A(n28292), .Z(n28256) );
  XOR U28352 ( .A(n28318), .B(n28319), .Z(n28292) );
  XOR U28353 ( .A(n28320), .B(n28321), .Z(n28319) );
  XOR U28354 ( .A(n28309), .B(n28322), .Z(n28318) );
  ANDN U28355 ( .B(n28242), .A(n28267), .Z(n28314) );
  XNOR U28356 ( .A(n28309), .B(n28323), .Z(n28267) );
  XOR U28357 ( .A(n28305), .B(n28231), .Z(n28242) );
  XNOR U28358 ( .A(n28324), .B(n28325), .Z(n28231) );
  XOR U28359 ( .A(n28326), .B(n28321), .Z(n28325) );
  XNOR U28360 ( .A(n28327), .B(n28328), .Z(n28321) );
  XNOR U28361 ( .A(n24320), .B(n26166), .Z(n28328) );
  XNOR U28362 ( .A(n26180), .B(n24339), .Z(n26166) );
  XNOR U28363 ( .A(n28329), .B(n28330), .Z(n24339) );
  XNOR U28364 ( .A(n28331), .B(n28332), .Z(n28330) );
  XNOR U28365 ( .A(n28333), .B(n28334), .Z(n28329) );
  XNOR U28366 ( .A(n28335), .B(n28336), .Z(n28334) );
  ANDN U28367 ( .B(n28337), .A(n28338), .Z(n28336) );
  XNOR U28368 ( .A(n25413), .B(n25399), .Z(n24320) );
  XOR U28369 ( .A(n28339), .B(n25370), .Z(n25399) );
  XNOR U28370 ( .A(n28340), .B(n24365), .Z(n25413) );
  IV U28371 ( .A(n26210), .Z(n24365) );
  XNOR U28372 ( .A(n24321), .B(n28341), .Z(n28327) );
  XNOR U28373 ( .A(key[228]), .B(n26167), .Z(n28341) );
  XOR U28374 ( .A(n25416), .B(n26184), .Z(n24321) );
  IV U28375 ( .A(n26714), .Z(n28305) );
  XOR U28376 ( .A(n28298), .B(n28342), .Z(n28312) );
  XNOR U28377 ( .A(n28343), .B(n28304), .Z(n28342) );
  OR U28378 ( .A(n26715), .B(n28247), .Z(n28304) );
  XNOR U28379 ( .A(n28323), .B(n28223), .Z(n28247) );
  XNOR U28380 ( .A(n26714), .B(n26663), .Z(n26715) );
  ANDN U28381 ( .B(n28223), .A(n26663), .Z(n28343) );
  XOR U28382 ( .A(n28324), .B(n28344), .Z(n26663) );
  XNOR U28383 ( .A(n28317), .B(n28345), .Z(n28344) );
  XOR U28384 ( .A(n28326), .B(n28324), .Z(n28223) );
  XNOR U28385 ( .A(n28248), .B(n26714), .Z(n28298) );
  XOR U28386 ( .A(n28324), .B(n28346), .Z(n26714) );
  XNOR U28387 ( .A(n28326), .B(n28320), .Z(n28346) );
  XOR U28388 ( .A(n28347), .B(n28348), .Z(n28320) );
  XNOR U28389 ( .A(n28349), .B(n24334), .Z(n28348) );
  XOR U28390 ( .A(n25382), .B(n26197), .Z(n24334) );
  XNOR U28391 ( .A(n28350), .B(n28351), .Z(n26197) );
  XNOR U28392 ( .A(n28352), .B(n28353), .Z(n28351) );
  XOR U28393 ( .A(n28354), .B(n28355), .Z(n28350) );
  XOR U28394 ( .A(n28356), .B(n28357), .Z(n25382) );
  XNOR U28395 ( .A(n28358), .B(n28359), .Z(n28357) );
  XNOR U28396 ( .A(key[231]), .B(n26180), .Z(n28347) );
  XNOR U28397 ( .A(n28360), .B(n28361), .Z(n28324) );
  XNOR U28398 ( .A(n24337), .B(n26196), .Z(n28361) );
  XNOR U28399 ( .A(n24347), .B(n24338), .Z(n26196) );
  XNOR U28400 ( .A(n28362), .B(n28363), .Z(n24347) );
  XNOR U28401 ( .A(n25401), .B(n25385), .Z(n24337) );
  XOR U28402 ( .A(n28364), .B(n28365), .Z(n25385) );
  XNOR U28403 ( .A(n28366), .B(n28353), .Z(n28365) );
  XNOR U28404 ( .A(n28367), .B(n28368), .Z(n28353) );
  XNOR U28405 ( .A(n28369), .B(n28370), .Z(n28368) );
  OR U28406 ( .A(n28371), .B(n28372), .Z(n28370) );
  XNOR U28407 ( .A(n28339), .B(n28373), .Z(n28364) );
  XNOR U28408 ( .A(n28374), .B(n28375), .Z(n28373) );
  ANDN U28409 ( .B(n28376), .A(n28377), .Z(n28375) );
  IV U28410 ( .A(n26183), .Z(n25401) );
  XNOR U28411 ( .A(n28378), .B(n28379), .Z(n26183) );
  XNOR U28412 ( .A(n28380), .B(n28359), .Z(n28379) );
  XNOR U28413 ( .A(n28381), .B(n28382), .Z(n28359) );
  XNOR U28414 ( .A(n28383), .B(n28384), .Z(n28382) );
  OR U28415 ( .A(n28385), .B(n28386), .Z(n28384) );
  XNOR U28416 ( .A(n28340), .B(n28387), .Z(n28378) );
  XNOR U28417 ( .A(n28388), .B(n28389), .Z(n28387) );
  ANDN U28418 ( .B(n28390), .A(n28391), .Z(n28389) );
  XOR U28419 ( .A(key[229]), .B(n26184), .Z(n28360) );
  XNOR U28420 ( .A(n28392), .B(n28393), .Z(n26184) );
  XNOR U28421 ( .A(n28394), .B(n28395), .Z(n28393) );
  XNOR U28422 ( .A(n28396), .B(n28397), .Z(n28392) );
  XOR U28423 ( .A(n28398), .B(n28399), .Z(n28397) );
  ANDN U28424 ( .B(n28400), .A(n28401), .Z(n28399) );
  IV U28425 ( .A(n28323), .Z(n28248) );
  XOR U28426 ( .A(n28345), .B(n28402), .Z(n28323) );
  XNOR U28427 ( .A(n28316), .B(n28322), .Z(n28402) );
  XOR U28428 ( .A(n28403), .B(n28404), .Z(n28322) );
  XOR U28429 ( .A(n28317), .B(n28405), .Z(n28404) );
  XNOR U28430 ( .A(n28406), .B(n26200), .Z(n28405) );
  XNOR U28431 ( .A(n26180), .B(n24319), .Z(n26200) );
  XNOR U28432 ( .A(n28333), .B(n24374), .Z(n24319) );
  XNOR U28433 ( .A(n28407), .B(n28408), .Z(n28317) );
  XNOR U28434 ( .A(n24363), .B(n25371), .Z(n28408) );
  XOR U28435 ( .A(n24367), .B(n24374), .Z(n25371) );
  XOR U28436 ( .A(n28409), .B(n28410), .Z(n24374) );
  XNOR U28437 ( .A(n26205), .B(n26193), .Z(n24363) );
  IV U28438 ( .A(n25410), .Z(n26193) );
  XOR U28439 ( .A(n28411), .B(n28412), .Z(n25410) );
  XNOR U28440 ( .A(n28354), .B(n28355), .Z(n28412) );
  IV U28441 ( .A(n24351), .Z(n26205) );
  XNOR U28442 ( .A(n28358), .B(n28413), .Z(n24351) );
  XNOR U28443 ( .A(n28414), .B(n28415), .Z(n28413) );
  XOR U28444 ( .A(key[225]), .B(n24352), .Z(n28407) );
  XOR U28445 ( .A(n24358), .B(n28416), .Z(n28403) );
  XNOR U28446 ( .A(key[227]), .B(n24370), .Z(n28416) );
  XNOR U28447 ( .A(n25416), .B(n26167), .Z(n24370) );
  XOR U28448 ( .A(n28394), .B(n28417), .Z(n26167) );
  IV U28449 ( .A(n25372), .Z(n24358) );
  XOR U28450 ( .A(n24377), .B(n25411), .Z(n25372) );
  XNOR U28451 ( .A(n28418), .B(n28419), .Z(n25411) );
  XNOR U28452 ( .A(n28352), .B(n28420), .Z(n28419) );
  XNOR U28453 ( .A(n28354), .B(n28421), .Z(n28418) );
  XNOR U28454 ( .A(n28423), .B(n28424), .Z(n28422) );
  OR U28455 ( .A(n28371), .B(n28425), .Z(n28424) );
  XOR U28456 ( .A(n28356), .B(n28427), .Z(n24377) );
  XOR U28457 ( .A(n28428), .B(n28429), .Z(n28427) );
  XOR U28458 ( .A(n28414), .B(n28415), .Z(n28356) );
  XOR U28459 ( .A(n28430), .B(n28431), .Z(n28415) );
  XNOR U28460 ( .A(n28432), .B(n28433), .Z(n28431) );
  OR U28461 ( .A(n28385), .B(n28434), .Z(n28433) );
  XOR U28462 ( .A(n28435), .B(n28436), .Z(n28316) );
  XOR U28463 ( .A(n24375), .B(n25404), .Z(n28436) );
  XOR U28464 ( .A(n24360), .B(n24373), .Z(n25404) );
  IV U28465 ( .A(n28406), .Z(n24373) );
  XNOR U28466 ( .A(n28437), .B(n28438), .Z(n28406) );
  XOR U28467 ( .A(n28439), .B(n28440), .Z(n28438) );
  XNOR U28468 ( .A(n28441), .B(n28442), .Z(n28437) );
  XNOR U28469 ( .A(n28443), .B(n28444), .Z(n24360) );
  XOR U28470 ( .A(n28410), .B(n28363), .Z(n28444) );
  XNOR U28471 ( .A(n28445), .B(n28446), .Z(n28363) );
  XOR U28472 ( .A(n28447), .B(n28335), .Z(n28446) );
  NANDN U28473 ( .A(n28448), .B(n28449), .Z(n28335) );
  ANDN U28474 ( .B(n28450), .A(n28451), .Z(n28447) );
  XOR U28475 ( .A(n28452), .B(n28453), .Z(n28443) );
  XNOR U28476 ( .A(n26210), .B(n25370), .Z(n24375) );
  XNOR U28477 ( .A(n28454), .B(n28352), .Z(n25370) );
  IV U28478 ( .A(n28411), .Z(n28352) );
  XOR U28479 ( .A(n28455), .B(n28456), .Z(n28411) );
  XOR U28480 ( .A(n28457), .B(n28458), .Z(n28456) );
  NANDN U28481 ( .A(n28459), .B(n28376), .Z(n28458) );
  XOR U28482 ( .A(n28460), .B(n28414), .Z(n26210) );
  XOR U28483 ( .A(n28461), .B(n28462), .Z(n28414) );
  XNOR U28484 ( .A(n28463), .B(n28464), .Z(n28462) );
  NANDN U28485 ( .A(n28465), .B(n28390), .Z(n28464) );
  XOR U28486 ( .A(key[226]), .B(n28417), .Z(n28435) );
  IV U28487 ( .A(n24367), .Z(n28417) );
  XNOR U28488 ( .A(n28441), .B(n28466), .Z(n24367) );
  IV U28489 ( .A(n28326), .Z(n28345) );
  XOR U28490 ( .A(n28467), .B(n28468), .Z(n28326) );
  XOR U28491 ( .A(n26189), .B(n26657), .Z(n28468) );
  IV U28492 ( .A(n28309), .Z(n26657) );
  XOR U28493 ( .A(n28469), .B(n28470), .Z(n28309) );
  XNOR U28494 ( .A(n24332), .B(n25409), .Z(n28470) );
  XNOR U28495 ( .A(n24352), .B(n24364), .Z(n25409) );
  XNOR U28496 ( .A(n28410), .B(n28471), .Z(n24364) );
  XNOR U28497 ( .A(n28452), .B(n28362), .Z(n28471) );
  XNOR U28498 ( .A(n28472), .B(n28473), .Z(n24352) );
  XOR U28499 ( .A(n28441), .B(n28442), .Z(n28473) );
  IV U28500 ( .A(n28474), .Z(n28441) );
  IV U28501 ( .A(n26192), .Z(n24332) );
  XOR U28502 ( .A(n25394), .B(n25416), .Z(n26192) );
  IV U28503 ( .A(n24355), .Z(n25394) );
  XOR U28504 ( .A(n28340), .B(n28475), .Z(n24355) );
  XNOR U28505 ( .A(n28381), .B(n28476), .Z(n28340) );
  XOR U28506 ( .A(n28477), .B(n28463), .Z(n28476) );
  NANDN U28507 ( .A(n28478), .B(n28479), .Z(n28463) );
  NOR U28508 ( .A(n28480), .B(n28481), .Z(n28477) );
  XNOR U28509 ( .A(n28461), .B(n28482), .Z(n28381) );
  XNOR U28510 ( .A(n28483), .B(n28484), .Z(n28482) );
  NANDN U28511 ( .A(n28485), .B(n28486), .Z(n28484) );
  XOR U28512 ( .A(key[224]), .B(n26179), .Z(n28469) );
  IV U28513 ( .A(n26169), .Z(n26179) );
  XOR U28514 ( .A(n28339), .B(n28487), .Z(n26169) );
  XNOR U28515 ( .A(n28367), .B(n28488), .Z(n28339) );
  XNOR U28516 ( .A(n28489), .B(n28457), .Z(n28488) );
  ANDN U28517 ( .B(n28490), .A(n28491), .Z(n28457) );
  ANDN U28518 ( .B(n28492), .A(n28493), .Z(n28489) );
  XOR U28519 ( .A(n28494), .B(n28495), .Z(n28367) );
  XNOR U28520 ( .A(n28496), .B(n28497), .Z(n28495) );
  NAND U28521 ( .A(n28498), .B(n28499), .Z(n28497) );
  XOR U28522 ( .A(n26180), .B(n24333), .Z(n26189) );
  IV U28523 ( .A(n26178), .Z(n24333) );
  XOR U28524 ( .A(n28500), .B(n28501), .Z(n26178) );
  XOR U28525 ( .A(n28410), .B(n28332), .Z(n28501) );
  XNOR U28526 ( .A(n28502), .B(n28503), .Z(n28332) );
  XNOR U28527 ( .A(n28504), .B(n28505), .Z(n28503) );
  OR U28528 ( .A(n28506), .B(n28507), .Z(n28505) );
  XNOR U28529 ( .A(n28508), .B(n28509), .Z(n28410) );
  XOR U28530 ( .A(n28510), .B(n28511), .Z(n28509) );
  NANDN U28531 ( .A(n28512), .B(n28337), .Z(n28511) );
  XOR U28532 ( .A(n28452), .B(n28362), .Z(n28500) );
  XOR U28533 ( .A(n28409), .B(n28453), .Z(n28362) );
  XOR U28534 ( .A(n28331), .B(n28513), .Z(n28453) );
  XNOR U28535 ( .A(n28514), .B(n28515), .Z(n28513) );
  NANDN U28536 ( .A(n28516), .B(n28517), .Z(n28515) );
  XNOR U28537 ( .A(n28514), .B(n28519), .Z(n28518) );
  OR U28538 ( .A(n28506), .B(n28520), .Z(n28519) );
  OR U28539 ( .A(n28521), .B(n28522), .Z(n28514) );
  XNOR U28540 ( .A(n28331), .B(n28523), .Z(n28445) );
  XNOR U28541 ( .A(n28524), .B(n28525), .Z(n28523) );
  NANDN U28542 ( .A(n28526), .B(n28527), .Z(n28525) );
  XOR U28543 ( .A(n28528), .B(n28524), .Z(n28331) );
  NANDN U28544 ( .A(n28529), .B(n28530), .Z(n28524) );
  ANDN U28545 ( .B(n28531), .A(n28532), .Z(n28528) );
  XOR U28546 ( .A(n28333), .B(n28409), .Z(n26180) );
  XOR U28547 ( .A(n28534), .B(n28504), .Z(n28533) );
  OR U28548 ( .A(n28535), .B(n28521), .Z(n28504) );
  ANDN U28549 ( .B(n28536), .A(n28516), .Z(n28534) );
  XNOR U28550 ( .A(n28502), .B(n28537), .Z(n28333) );
  XNOR U28551 ( .A(n28538), .B(n28510), .Z(n28537) );
  ANDN U28552 ( .B(n28449), .A(n28539), .Z(n28510) );
  XOR U28553 ( .A(n28450), .B(n28337), .Z(n28449) );
  ANDN U28554 ( .B(n28450), .A(n28540), .Z(n28538) );
  XOR U28555 ( .A(n28508), .B(n28541), .Z(n28502) );
  XNOR U28556 ( .A(n28542), .B(n28543), .Z(n28541) );
  NAND U28557 ( .A(n28527), .B(n28544), .Z(n28543) );
  XNOR U28558 ( .A(n28545), .B(n28542), .Z(n28508) );
  OR U28559 ( .A(n28529), .B(n28546), .Z(n28542) );
  XNOR U28560 ( .A(n28547), .B(n28527), .Z(n28529) );
  XNOR U28561 ( .A(n28516), .B(n28337), .Z(n28527) );
  XOR U28562 ( .A(n28548), .B(n28549), .Z(n28337) );
  NANDN U28563 ( .A(n28550), .B(n28551), .Z(n28549) );
  XNOR U28564 ( .A(n28552), .B(n28553), .Z(n28516) );
  NANDN U28565 ( .A(n28550), .B(n28554), .Z(n28553) );
  ANDN U28566 ( .B(n28547), .A(n28555), .Z(n28545) );
  IV U28567 ( .A(n28532), .Z(n28547) );
  XOR U28568 ( .A(n28450), .B(n28506), .Z(n28532) );
  XOR U28569 ( .A(n28556), .B(n28552), .Z(n28506) );
  NANDN U28570 ( .A(n28557), .B(n28558), .Z(n28552) );
  NANDN U28571 ( .A(n28557), .B(n28562), .Z(n28548) );
  XOR U28572 ( .A(n28563), .B(n28564), .Z(n28550) );
  XOR U28573 ( .A(n28565), .B(n28560), .Z(n28564) );
  XNOR U28574 ( .A(n28566), .B(n28567), .Z(n28563) );
  XNOR U28575 ( .A(n28568), .B(n28569), .Z(n28567) );
  ANDN U28576 ( .B(n28565), .A(n28560), .Z(n28568) );
  ANDN U28577 ( .B(n28565), .A(n28559), .Z(n28561) );
  XNOR U28578 ( .A(n28566), .B(n28570), .Z(n28559) );
  XOR U28579 ( .A(n28571), .B(n28569), .Z(n28570) );
  NAND U28580 ( .A(n28558), .B(n28562), .Z(n28569) );
  XNOR U28581 ( .A(n28554), .B(n28560), .Z(n28558) );
  XOR U28582 ( .A(n28572), .B(n28573), .Z(n28560) );
  XOR U28583 ( .A(n28574), .B(n28575), .Z(n28573) );
  XNOR U28584 ( .A(n28576), .B(n28577), .Z(n28572) );
  ANDN U28585 ( .B(n28578), .A(n28451), .Z(n28576) );
  AND U28586 ( .A(n28551), .B(n28554), .Z(n28571) );
  XNOR U28587 ( .A(n28551), .B(n28554), .Z(n28566) );
  XNOR U28588 ( .A(n28579), .B(n28580), .Z(n28554) );
  XNOR U28589 ( .A(n28581), .B(n28582), .Z(n28580) );
  XOR U28590 ( .A(n28574), .B(n28583), .Z(n28579) );
  XNOR U28591 ( .A(n28584), .B(n28577), .Z(n28583) );
  OR U28592 ( .A(n28448), .B(n28539), .Z(n28577) );
  XNOR U28593 ( .A(n28540), .B(n28512), .Z(n28539) );
  XNOR U28594 ( .A(n28451), .B(n28338), .Z(n28448) );
  NOR U28595 ( .A(n28338), .B(n28512), .Z(n28584) );
  XNOR U28596 ( .A(n28585), .B(n28586), .Z(n28551) );
  XNOR U28597 ( .A(n28587), .B(n28588), .Z(n28586) );
  XOR U28598 ( .A(n28520), .B(n28574), .Z(n28588) );
  XOR U28599 ( .A(n28578), .B(n28589), .Z(n28574) );
  XNOR U28600 ( .A(n28507), .B(n28590), .Z(n28585) );
  XNOR U28601 ( .A(n28591), .B(n28592), .Z(n28590) );
  ANDN U28602 ( .B(n28517), .A(n28593), .Z(n28591) );
  XNOR U28603 ( .A(n28594), .B(n28595), .Z(n28565) );
  XNOR U28604 ( .A(n28575), .B(n28596), .Z(n28595) );
  XNOR U28605 ( .A(n28517), .B(n28582), .Z(n28596) );
  XOR U28606 ( .A(n28512), .B(n28338), .Z(n28582) );
  XNOR U28607 ( .A(n28587), .B(n28597), .Z(n28575) );
  XNOR U28608 ( .A(n28598), .B(n28599), .Z(n28597) );
  NANDN U28609 ( .A(n28526), .B(n28544), .Z(n28599) );
  IV U28610 ( .A(n28581), .Z(n28587) );
  XNOR U28611 ( .A(n28600), .B(n28598), .Z(n28581) );
  NANDN U28612 ( .A(n28546), .B(n28530), .Z(n28598) );
  XOR U28613 ( .A(n28517), .B(n28338), .Z(n28526) );
  XOR U28614 ( .A(n28601), .B(n28602), .Z(n28338) );
  XNOR U28615 ( .A(n28603), .B(n28604), .Z(n28602) );
  XOR U28616 ( .A(n28555), .B(n28544), .Z(n28546) );
  XNOR U28617 ( .A(n28536), .B(n28512), .Z(n28544) );
  XNOR U28618 ( .A(n28604), .B(n28605), .Z(n28512) );
  ANDN U28619 ( .B(n28531), .A(n28555), .Z(n28600) );
  XNOR U28620 ( .A(n28606), .B(n28578), .Z(n28555) );
  IV U28621 ( .A(n28540), .Z(n28578) );
  XNOR U28622 ( .A(n28607), .B(n28608), .Z(n28540) );
  XNOR U28623 ( .A(n28609), .B(n28604), .Z(n28608) );
  XOR U28624 ( .A(n28610), .B(n28589), .Z(n28531) );
  XNOR U28625 ( .A(n28593), .B(n28611), .Z(n28594) );
  XNOR U28626 ( .A(n28612), .B(n28592), .Z(n28611) );
  OR U28627 ( .A(n28522), .B(n28535), .Z(n28592) );
  XOR U28628 ( .A(n28507), .B(n28536), .Z(n28535) );
  IV U28629 ( .A(n28593), .Z(n28536) );
  XOR U28630 ( .A(n28520), .B(n28517), .Z(n28522) );
  XNOR U28631 ( .A(n28589), .B(n28613), .Z(n28517) );
  XNOR U28632 ( .A(n28603), .B(n28607), .Z(n28613) );
  XNOR U28633 ( .A(msg[2]), .B(key[2]), .Z(n28607) );
  IV U28634 ( .A(n28451), .Z(n28589) );
  XOR U28635 ( .A(n28601), .B(n28614), .Z(n28451) );
  XOR U28636 ( .A(n28604), .B(n28615), .Z(n28614) );
  IV U28637 ( .A(n28610), .Z(n28520) );
  ANDN U28638 ( .B(n28610), .A(n28507), .Z(n28612) );
  XOR U28639 ( .A(n28605), .B(n28616), .Z(n28610) );
  XNOR U28640 ( .A(n28604), .B(n28617), .Z(n28616) );
  XOR U28641 ( .A(n28606), .B(n28618), .Z(n28604) );
  XNOR U28642 ( .A(msg[6]), .B(key[6]), .Z(n28618) );
  IV U28643 ( .A(n28601), .Z(n28605) );
  XOR U28644 ( .A(msg[5]), .B(key[5]), .Z(n28601) );
  XOR U28645 ( .A(n28619), .B(n28620), .Z(n28593) );
  XOR U28646 ( .A(n28617), .B(n28615), .Z(n28620) );
  XOR U28647 ( .A(msg[7]), .B(key[7]), .Z(n28615) );
  XNOR U28648 ( .A(msg[4]), .B(key[4]), .Z(n28617) );
  XOR U28649 ( .A(n28507), .B(n28609), .Z(n28619) );
  XNOR U28650 ( .A(n28603), .B(n28621), .Z(n28609) );
  XNOR U28651 ( .A(msg[3]), .B(key[3]), .Z(n28621) );
  XNOR U28652 ( .A(msg[1]), .B(key[1]), .Z(n28603) );
  IV U28653 ( .A(n28606), .Z(n28507) );
  XOR U28654 ( .A(msg[0]), .B(key[0]), .Z(n28606) );
  XOR U28655 ( .A(n24338), .B(n28622), .Z(n28467) );
  XOR U28656 ( .A(key[230]), .B(n24346), .Z(n28622) );
  XNOR U28657 ( .A(n25387), .B(n28349), .Z(n24346) );
  XOR U28658 ( .A(n25416), .B(n26177), .Z(n28349) );
  XNOR U28659 ( .A(n28623), .B(n28624), .Z(n26177) );
  XOR U28660 ( .A(n28472), .B(n28395), .Z(n28624) );
  XNOR U28661 ( .A(n28625), .B(n28626), .Z(n28395) );
  XNOR U28662 ( .A(n28627), .B(n28628), .Z(n28626) );
  NANDN U28663 ( .A(n28629), .B(n28630), .Z(n28628) );
  XOR U28664 ( .A(n28474), .B(n28442), .Z(n28623) );
  XNOR U28665 ( .A(n28632), .B(n28633), .Z(n28631) );
  NANDN U28666 ( .A(n28629), .B(n28634), .Z(n28633) );
  XOR U28667 ( .A(n28637), .B(n28638), .Z(n28636) );
  NANDN U28668 ( .A(n28639), .B(n28640), .Z(n28638) );
  XOR U28669 ( .A(n28642), .B(n28394), .Z(n25416) );
  XNOR U28670 ( .A(n28625), .B(n28643), .Z(n28394) );
  XNOR U28671 ( .A(n28644), .B(n28637), .Z(n28643) );
  NOR U28672 ( .A(n28645), .B(n28646), .Z(n28637) );
  ANDN U28673 ( .B(n28647), .A(n28648), .Z(n28644) );
  XOR U28674 ( .A(n28641), .B(n28649), .Z(n28625) );
  XNOR U28675 ( .A(n28650), .B(n28651), .Z(n28649) );
  NANDN U28676 ( .A(n28652), .B(n28653), .Z(n28651) );
  XOR U28677 ( .A(n24341), .B(n25380), .Z(n25387) );
  XOR U28678 ( .A(n28355), .B(n28420), .Z(n25380) );
  XNOR U28679 ( .A(n28426), .B(n28654), .Z(n28420) );
  XOR U28680 ( .A(n28655), .B(n28374), .Z(n28654) );
  NANDN U28681 ( .A(n28656), .B(n28490), .Z(n28374) );
  XOR U28682 ( .A(n28492), .B(n28376), .Z(n28490) );
  ANDN U28683 ( .B(n28492), .A(n28657), .Z(n28655) );
  XNOR U28684 ( .A(n28366), .B(n28658), .Z(n28426) );
  XNOR U28685 ( .A(n28659), .B(n28660), .Z(n28658) );
  NANDN U28686 ( .A(n28661), .B(n28498), .Z(n28660) );
  XOR U28687 ( .A(n28454), .B(n28421), .Z(n28355) );
  XNOR U28688 ( .A(n28366), .B(n28662), .Z(n28421) );
  XNOR U28689 ( .A(n28423), .B(n28663), .Z(n28662) );
  NANDN U28690 ( .A(n28664), .B(n28665), .Z(n28663) );
  OR U28691 ( .A(n28666), .B(n28667), .Z(n28423) );
  XOR U28692 ( .A(n28668), .B(n28659), .Z(n28366) );
  NANDN U28693 ( .A(n28669), .B(n28670), .Z(n28659) );
  ANDN U28694 ( .B(n28671), .A(n28672), .Z(n28668) );
  IV U28695 ( .A(n28487), .Z(n28454) );
  XOR U28696 ( .A(n28455), .B(n28673), .Z(n28487) );
  XOR U28697 ( .A(n28674), .B(n28369), .Z(n28673) );
  OR U28698 ( .A(n28675), .B(n28666), .Z(n28369) );
  ANDN U28699 ( .B(n28676), .A(n28664), .Z(n28674) );
  IV U28700 ( .A(n28494), .Z(n28455) );
  XNOR U28701 ( .A(n28677), .B(n28496), .Z(n28494) );
  OR U28702 ( .A(n28669), .B(n28678), .Z(n28496) );
  XNOR U28703 ( .A(n28679), .B(n28498), .Z(n28669) );
  XNOR U28704 ( .A(n28664), .B(n28376), .Z(n28498) );
  XOR U28705 ( .A(n28680), .B(n28681), .Z(n28376) );
  NANDN U28706 ( .A(n28682), .B(n28683), .Z(n28681) );
  XNOR U28707 ( .A(n28684), .B(n28685), .Z(n28664) );
  NANDN U28708 ( .A(n28682), .B(n28686), .Z(n28685) );
  ANDN U28709 ( .B(n28679), .A(n28687), .Z(n28677) );
  IV U28710 ( .A(n28672), .Z(n28679) );
  XOR U28711 ( .A(n28492), .B(n28371), .Z(n28672) );
  XOR U28712 ( .A(n28688), .B(n28684), .Z(n28371) );
  NANDN U28713 ( .A(n28689), .B(n28690), .Z(n28684) );
  NANDN U28714 ( .A(n28689), .B(n28694), .Z(n28680) );
  XOR U28715 ( .A(n28695), .B(n28696), .Z(n28682) );
  XOR U28716 ( .A(n28697), .B(n28692), .Z(n28696) );
  XNOR U28717 ( .A(n28698), .B(n28699), .Z(n28695) );
  XNOR U28718 ( .A(n28700), .B(n28701), .Z(n28699) );
  ANDN U28719 ( .B(n28697), .A(n28692), .Z(n28700) );
  ANDN U28720 ( .B(n28697), .A(n28691), .Z(n28693) );
  XNOR U28721 ( .A(n28698), .B(n28702), .Z(n28691) );
  XOR U28722 ( .A(n28703), .B(n28701), .Z(n28702) );
  NAND U28723 ( .A(n28690), .B(n28694), .Z(n28701) );
  XNOR U28724 ( .A(n28686), .B(n28692), .Z(n28690) );
  XOR U28725 ( .A(n28704), .B(n28705), .Z(n28692) );
  XOR U28726 ( .A(n28706), .B(n28707), .Z(n28705) );
  XNOR U28727 ( .A(n28708), .B(n28709), .Z(n28704) );
  ANDN U28728 ( .B(n28710), .A(n28657), .Z(n28708) );
  AND U28729 ( .A(n28683), .B(n28686), .Z(n28703) );
  XNOR U28730 ( .A(n28683), .B(n28686), .Z(n28698) );
  XNOR U28731 ( .A(n28711), .B(n28712), .Z(n28686) );
  XNOR U28732 ( .A(n28713), .B(n28714), .Z(n28712) );
  XOR U28733 ( .A(n28706), .B(n28715), .Z(n28711) );
  XNOR U28734 ( .A(n28716), .B(n28709), .Z(n28715) );
  OR U28735 ( .A(n28656), .B(n28491), .Z(n28709) );
  XNOR U28736 ( .A(n28493), .B(n28459), .Z(n28491) );
  XNOR U28737 ( .A(n28657), .B(n28377), .Z(n28656) );
  NOR U28738 ( .A(n28377), .B(n28459), .Z(n28716) );
  XNOR U28739 ( .A(n28717), .B(n28718), .Z(n28683) );
  XNOR U28740 ( .A(n28719), .B(n28720), .Z(n28718) );
  XOR U28741 ( .A(n28425), .B(n28706), .Z(n28720) );
  XOR U28742 ( .A(n28710), .B(n28721), .Z(n28706) );
  XNOR U28743 ( .A(n28372), .B(n28722), .Z(n28717) );
  XNOR U28744 ( .A(n28723), .B(n28724), .Z(n28722) );
  ANDN U28745 ( .B(n28665), .A(n28725), .Z(n28723) );
  XNOR U28746 ( .A(n28726), .B(n28727), .Z(n28697) );
  XNOR U28747 ( .A(n28707), .B(n28728), .Z(n28727) );
  XNOR U28748 ( .A(n28665), .B(n28714), .Z(n28728) );
  XOR U28749 ( .A(n28459), .B(n28377), .Z(n28714) );
  XNOR U28750 ( .A(n28719), .B(n28729), .Z(n28707) );
  XNOR U28751 ( .A(n28730), .B(n28731), .Z(n28729) );
  NANDN U28752 ( .A(n28661), .B(n28499), .Z(n28731) );
  IV U28753 ( .A(n28713), .Z(n28719) );
  XNOR U28754 ( .A(n28732), .B(n28730), .Z(n28713) );
  NANDN U28755 ( .A(n28678), .B(n28670), .Z(n28730) );
  XOR U28756 ( .A(n28665), .B(n28377), .Z(n28661) );
  XOR U28757 ( .A(n28733), .B(n28734), .Z(n28377) );
  XNOR U28758 ( .A(n28735), .B(n28736), .Z(n28734) );
  XOR U28759 ( .A(n28687), .B(n28499), .Z(n28678) );
  XNOR U28760 ( .A(n28676), .B(n28459), .Z(n28499) );
  XNOR U28761 ( .A(n28736), .B(n28737), .Z(n28459) );
  ANDN U28762 ( .B(n28671), .A(n28687), .Z(n28732) );
  XNOR U28763 ( .A(n28738), .B(n28710), .Z(n28687) );
  IV U28764 ( .A(n28493), .Z(n28710) );
  XNOR U28765 ( .A(n28739), .B(n28740), .Z(n28493) );
  XNOR U28766 ( .A(n28741), .B(n28736), .Z(n28740) );
  XOR U28767 ( .A(n28742), .B(n28721), .Z(n28671) );
  XNOR U28768 ( .A(n28725), .B(n28743), .Z(n28726) );
  XNOR U28769 ( .A(n28744), .B(n28724), .Z(n28743) );
  OR U28770 ( .A(n28667), .B(n28675), .Z(n28724) );
  XOR U28771 ( .A(n28372), .B(n28676), .Z(n28675) );
  IV U28772 ( .A(n28725), .Z(n28676) );
  XOR U28773 ( .A(n28425), .B(n28665), .Z(n28667) );
  XNOR U28774 ( .A(n28721), .B(n28745), .Z(n28665) );
  XNOR U28775 ( .A(n28735), .B(n28739), .Z(n28745) );
  XNOR U28776 ( .A(msg[42]), .B(key[42]), .Z(n28739) );
  IV U28777 ( .A(n28657), .Z(n28721) );
  XOR U28778 ( .A(n28733), .B(n28746), .Z(n28657) );
  XOR U28779 ( .A(n28736), .B(n28747), .Z(n28746) );
  IV U28780 ( .A(n28742), .Z(n28425) );
  ANDN U28781 ( .B(n28742), .A(n28372), .Z(n28744) );
  XOR U28782 ( .A(n28737), .B(n28748), .Z(n28742) );
  XNOR U28783 ( .A(n28736), .B(n28749), .Z(n28748) );
  XOR U28784 ( .A(n28738), .B(n28750), .Z(n28736) );
  XNOR U28785 ( .A(msg[46]), .B(key[46]), .Z(n28750) );
  IV U28786 ( .A(n28733), .Z(n28737) );
  XOR U28787 ( .A(msg[45]), .B(key[45]), .Z(n28733) );
  XOR U28788 ( .A(n28751), .B(n28752), .Z(n28725) );
  XOR U28789 ( .A(n28749), .B(n28747), .Z(n28752) );
  XOR U28790 ( .A(msg[47]), .B(key[47]), .Z(n28747) );
  XNOR U28791 ( .A(msg[44]), .B(key[44]), .Z(n28749) );
  XOR U28792 ( .A(n28372), .B(n28741), .Z(n28751) );
  XNOR U28793 ( .A(n28735), .B(n28753), .Z(n28741) );
  XNOR U28794 ( .A(msg[43]), .B(key[43]), .Z(n28753) );
  XNOR U28795 ( .A(msg[41]), .B(key[41]), .Z(n28735) );
  IV U28796 ( .A(n28738), .Z(n28372) );
  XOR U28797 ( .A(msg[40]), .B(key[40]), .Z(n28738) );
  XNOR U28798 ( .A(n28358), .B(n28429), .Z(n24341) );
  XNOR U28799 ( .A(n28430), .B(n28754), .Z(n28429) );
  XOR U28800 ( .A(n28755), .B(n28388), .Z(n28754) );
  NANDN U28801 ( .A(n28756), .B(n28479), .Z(n28388) );
  XNOR U28802 ( .A(n28481), .B(n28390), .Z(n28479) );
  NOR U28803 ( .A(n28757), .B(n28481), .Z(n28755) );
  XNOR U28804 ( .A(n28380), .B(n28758), .Z(n28430) );
  XNOR U28805 ( .A(n28759), .B(n28760), .Z(n28758) );
  OR U28806 ( .A(n28485), .B(n28761), .Z(n28760) );
  XNOR U28807 ( .A(n28460), .B(n28428), .Z(n28358) );
  XOR U28808 ( .A(n28380), .B(n28762), .Z(n28428) );
  XNOR U28809 ( .A(n28432), .B(n28763), .Z(n28762) );
  NANDN U28810 ( .A(n28764), .B(n28765), .Z(n28763) );
  OR U28811 ( .A(n28766), .B(n28767), .Z(n28432) );
  XOR U28812 ( .A(n28768), .B(n28759), .Z(n28380) );
  NANDN U28813 ( .A(n28769), .B(n28770), .Z(n28759) );
  AND U28814 ( .A(n28771), .B(n28772), .Z(n28768) );
  IV U28815 ( .A(n28475), .Z(n28460) );
  XNOR U28816 ( .A(n28461), .B(n28773), .Z(n28475) );
  XOR U28817 ( .A(n28774), .B(n28383), .Z(n28773) );
  OR U28818 ( .A(n28775), .B(n28766), .Z(n28383) );
  XOR U28819 ( .A(n28385), .B(n28776), .Z(n28766) );
  ANDN U28820 ( .B(n28777), .A(n28764), .Z(n28774) );
  XOR U28821 ( .A(n28778), .B(n28483), .Z(n28461) );
  OR U28822 ( .A(n28769), .B(n28779), .Z(n28483) );
  XOR U28823 ( .A(n28771), .B(n28485), .Z(n28769) );
  XNOR U28824 ( .A(n28776), .B(n28390), .Z(n28485) );
  XOR U28825 ( .A(n28780), .B(n28781), .Z(n28390) );
  NANDN U28826 ( .A(n28782), .B(n28783), .Z(n28781) );
  IV U28827 ( .A(n28764), .Z(n28776) );
  XNOR U28828 ( .A(n28784), .B(n28785), .Z(n28764) );
  NANDN U28829 ( .A(n28782), .B(n28786), .Z(n28785) );
  ANDN U28830 ( .B(n28771), .A(n28787), .Z(n28778) );
  XOR U28831 ( .A(n28481), .B(n28385), .Z(n28771) );
  XOR U28832 ( .A(n28788), .B(n28784), .Z(n28385) );
  NANDN U28833 ( .A(n28789), .B(n28790), .Z(n28784) );
  NANDN U28834 ( .A(n28789), .B(n28794), .Z(n28780) );
  XOR U28835 ( .A(n28795), .B(n28796), .Z(n28782) );
  XOR U28836 ( .A(n28797), .B(n28792), .Z(n28796) );
  XNOR U28837 ( .A(n28798), .B(n28799), .Z(n28795) );
  XNOR U28838 ( .A(n28800), .B(n28801), .Z(n28799) );
  ANDN U28839 ( .B(n28797), .A(n28792), .Z(n28800) );
  ANDN U28840 ( .B(n28797), .A(n28791), .Z(n28793) );
  XNOR U28841 ( .A(n28798), .B(n28802), .Z(n28791) );
  XOR U28842 ( .A(n28803), .B(n28801), .Z(n28802) );
  NAND U28843 ( .A(n28790), .B(n28794), .Z(n28801) );
  XNOR U28844 ( .A(n28786), .B(n28792), .Z(n28790) );
  XOR U28845 ( .A(n28804), .B(n28805), .Z(n28792) );
  XOR U28846 ( .A(n28806), .B(n28807), .Z(n28805) );
  XNOR U28847 ( .A(n28808), .B(n28809), .Z(n28804) );
  ANDN U28848 ( .B(n28810), .A(n28757), .Z(n28808) );
  AND U28849 ( .A(n28783), .B(n28786), .Z(n28803) );
  XNOR U28850 ( .A(n28783), .B(n28786), .Z(n28798) );
  XNOR U28851 ( .A(n28811), .B(n28812), .Z(n28786) );
  XNOR U28852 ( .A(n28813), .B(n28814), .Z(n28812) );
  XOR U28853 ( .A(n28806), .B(n28815), .Z(n28811) );
  XNOR U28854 ( .A(n28816), .B(n28809), .Z(n28815) );
  OR U28855 ( .A(n28756), .B(n28478), .Z(n28809) );
  XNOR U28856 ( .A(n28480), .B(n28465), .Z(n28478) );
  XNOR U28857 ( .A(n28757), .B(n28391), .Z(n28756) );
  NOR U28858 ( .A(n28391), .B(n28465), .Z(n28816) );
  XNOR U28859 ( .A(n28817), .B(n28818), .Z(n28783) );
  XNOR U28860 ( .A(n28819), .B(n28820), .Z(n28818) );
  XOR U28861 ( .A(n28434), .B(n28806), .Z(n28820) );
  XOR U28862 ( .A(n28810), .B(n28821), .Z(n28806) );
  XNOR U28863 ( .A(n28386), .B(n28822), .Z(n28817) );
  XNOR U28864 ( .A(n28823), .B(n28824), .Z(n28822) );
  ANDN U28865 ( .B(n28765), .A(n28825), .Z(n28823) );
  XNOR U28866 ( .A(n28826), .B(n28827), .Z(n28797) );
  XNOR U28867 ( .A(n28807), .B(n28828), .Z(n28827) );
  XNOR U28868 ( .A(n28765), .B(n28814), .Z(n28828) );
  XOR U28869 ( .A(n28465), .B(n28391), .Z(n28814) );
  XNOR U28870 ( .A(n28819), .B(n28829), .Z(n28807) );
  XNOR U28871 ( .A(n28830), .B(n28831), .Z(n28829) );
  NANDN U28872 ( .A(n28761), .B(n28486), .Z(n28831) );
  IV U28873 ( .A(n28813), .Z(n28819) );
  XNOR U28874 ( .A(n28832), .B(n28830), .Z(n28813) );
  NANDN U28875 ( .A(n28779), .B(n28770), .Z(n28830) );
  XOR U28876 ( .A(n28765), .B(n28391), .Z(n28761) );
  XOR U28877 ( .A(n28833), .B(n28834), .Z(n28391) );
  XNOR U28878 ( .A(n28835), .B(n28836), .Z(n28834) );
  XOR U28879 ( .A(n28787), .B(n28486), .Z(n28779) );
  XNOR U28880 ( .A(n28777), .B(n28465), .Z(n28486) );
  XNOR U28881 ( .A(n28836), .B(n28837), .Z(n28465) );
  ANDN U28882 ( .B(n28772), .A(n28787), .Z(n28832) );
  XNOR U28883 ( .A(n28838), .B(n28810), .Z(n28787) );
  IV U28884 ( .A(n28480), .Z(n28810) );
  XNOR U28885 ( .A(n28839), .B(n28840), .Z(n28480) );
  XNOR U28886 ( .A(n28841), .B(n28836), .Z(n28840) );
  XOR U28887 ( .A(n28842), .B(n28821), .Z(n28772) );
  XNOR U28888 ( .A(n28825), .B(n28843), .Z(n28826) );
  XNOR U28889 ( .A(n28844), .B(n28824), .Z(n28843) );
  OR U28890 ( .A(n28767), .B(n28775), .Z(n28824) );
  XOR U28891 ( .A(n28386), .B(n28777), .Z(n28775) );
  IV U28892 ( .A(n28825), .Z(n28777) );
  XOR U28893 ( .A(n28434), .B(n28765), .Z(n28767) );
  XNOR U28894 ( .A(n28821), .B(n28845), .Z(n28765) );
  XNOR U28895 ( .A(n28835), .B(n28839), .Z(n28845) );
  XNOR U28896 ( .A(msg[82]), .B(key[82]), .Z(n28839) );
  IV U28897 ( .A(n28757), .Z(n28821) );
  XOR U28898 ( .A(n28833), .B(n28846), .Z(n28757) );
  XOR U28899 ( .A(n28836), .B(n28847), .Z(n28846) );
  IV U28900 ( .A(n28842), .Z(n28434) );
  ANDN U28901 ( .B(n28842), .A(n28386), .Z(n28844) );
  XOR U28902 ( .A(n28837), .B(n28848), .Z(n28842) );
  XNOR U28903 ( .A(n28836), .B(n28849), .Z(n28848) );
  XOR U28904 ( .A(n28838), .B(n28850), .Z(n28836) );
  XNOR U28905 ( .A(msg[86]), .B(key[86]), .Z(n28850) );
  IV U28906 ( .A(n28833), .Z(n28837) );
  XOR U28907 ( .A(msg[85]), .B(key[85]), .Z(n28833) );
  XOR U28908 ( .A(n28851), .B(n28852), .Z(n28825) );
  XOR U28909 ( .A(n28849), .B(n28847), .Z(n28852) );
  XOR U28910 ( .A(msg[87]), .B(key[87]), .Z(n28847) );
  XNOR U28911 ( .A(msg[84]), .B(key[84]), .Z(n28849) );
  XOR U28912 ( .A(n28386), .B(n28841), .Z(n28851) );
  XNOR U28913 ( .A(n28835), .B(n28853), .Z(n28841) );
  XNOR U28914 ( .A(msg[83]), .B(key[83]), .Z(n28853) );
  XNOR U28915 ( .A(msg[81]), .B(key[81]), .Z(n28835) );
  IV U28916 ( .A(n28838), .Z(n28386) );
  XOR U28917 ( .A(msg[80]), .B(key[80]), .Z(n28838) );
  XNOR U28918 ( .A(n28472), .B(n28440), .Z(n24338) );
  XNOR U28919 ( .A(n28635), .B(n28854), .Z(n28440) );
  XNOR U28920 ( .A(n28855), .B(n28398), .Z(n28854) );
  NOR U28921 ( .A(n28645), .B(n28856), .Z(n28398) );
  XNOR U28922 ( .A(n28647), .B(n28640), .Z(n28645) );
  AND U28923 ( .A(n28647), .B(n28857), .Z(n28855) );
  XNOR U28924 ( .A(n28396), .B(n28858), .Z(n28635) );
  XNOR U28925 ( .A(n28859), .B(n28860), .Z(n28858) );
  NANDN U28926 ( .A(n28652), .B(n28861), .Z(n28860) );
  XOR U28927 ( .A(n28642), .B(n28439), .Z(n28472) );
  XOR U28928 ( .A(n28396), .B(n28862), .Z(n28439) );
  XNOR U28929 ( .A(n28632), .B(n28863), .Z(n28862) );
  NANDN U28930 ( .A(n28864), .B(n28865), .Z(n28863) );
  OR U28931 ( .A(n28866), .B(n28867), .Z(n28632) );
  XOR U28932 ( .A(n28868), .B(n28859), .Z(n28396) );
  NANDN U28933 ( .A(n28869), .B(n28870), .Z(n28859) );
  ANDN U28934 ( .B(n28871), .A(n28872), .Z(n28868) );
  IV U28935 ( .A(n28466), .Z(n28642) );
  XOR U28936 ( .A(n28641), .B(n28873), .Z(n28466) );
  XOR U28937 ( .A(n28874), .B(n28627), .Z(n28873) );
  OR U28938 ( .A(n28875), .B(n28866), .Z(n28627) );
  XOR U28939 ( .A(n28629), .B(n28865), .Z(n28866) );
  ANDN U28940 ( .B(n28865), .A(n28876), .Z(n28874) );
  XNOR U28941 ( .A(n28877), .B(n28650), .Z(n28641) );
  OR U28942 ( .A(n28869), .B(n28878), .Z(n28650) );
  XNOR U28943 ( .A(n28872), .B(n28652), .Z(n28869) );
  XNOR U28944 ( .A(n28865), .B(n28640), .Z(n28652) );
  IV U28945 ( .A(n28401), .Z(n28640) );
  XNOR U28946 ( .A(n28879), .B(n28880), .Z(n28401) );
  NANDN U28947 ( .A(n28881), .B(n28882), .Z(n28880) );
  XOR U28948 ( .A(n28883), .B(n28884), .Z(n28865) );
  NANDN U28949 ( .A(n28881), .B(n28885), .Z(n28884) );
  XOR U28950 ( .A(n28629), .B(n28647), .Z(n28872) );
  XNOR U28951 ( .A(n28887), .B(n28879), .Z(n28647) );
  NANDN U28952 ( .A(n28888), .B(n28889), .Z(n28879) );
  XOR U28953 ( .A(n28882), .B(n28890), .Z(n28889) );
  ANDN U28954 ( .B(n28890), .A(n28891), .Z(n28887) );
  NANDN U28955 ( .A(n28888), .B(n28893), .Z(n28883) );
  XOR U28956 ( .A(n28894), .B(n28895), .Z(n28881) );
  XOR U28957 ( .A(n28896), .B(n28897), .Z(n28895) );
  XNOR U28958 ( .A(n28898), .B(n28899), .Z(n28894) );
  XNOR U28959 ( .A(n28900), .B(n28901), .Z(n28899) );
  ANDN U28960 ( .B(n28897), .A(n28896), .Z(n28900) );
  ANDN U28961 ( .B(n28897), .A(n28891), .Z(n28892) );
  XNOR U28962 ( .A(n28898), .B(n28902), .Z(n28891) );
  XOR U28963 ( .A(n28903), .B(n28901), .Z(n28902) );
  NAND U28964 ( .A(n28893), .B(n28904), .Z(n28901) );
  XNOR U28965 ( .A(n28882), .B(n28896), .Z(n28904) );
  IV U28966 ( .A(n28890), .Z(n28896) );
  XNOR U28967 ( .A(n28905), .B(n28906), .Z(n28890) );
  XNOR U28968 ( .A(n28907), .B(n28908), .Z(n28906) );
  XOR U28969 ( .A(n28864), .B(n28909), .Z(n28908) );
  XNOR U28970 ( .A(n28876), .B(n28910), .Z(n28905) );
  XNOR U28971 ( .A(n28911), .B(n28912), .Z(n28910) );
  AND U28972 ( .A(n28634), .B(n28630), .Z(n28911) );
  XOR U28973 ( .A(n28885), .B(n28897), .Z(n28893) );
  AND U28974 ( .A(n28882), .B(n28885), .Z(n28903) );
  XNOR U28975 ( .A(n28882), .B(n28885), .Z(n28898) );
  XNOR U28976 ( .A(n28913), .B(n28914), .Z(n28885) );
  XNOR U28977 ( .A(n28915), .B(n28909), .Z(n28914) );
  XOR U28978 ( .A(n28916), .B(n28917), .Z(n28913) );
  XNOR U28979 ( .A(n28918), .B(n28919), .Z(n28917) );
  ANDN U28980 ( .B(n28400), .A(n28639), .Z(n28918) );
  XNOR U28981 ( .A(n28920), .B(n28921), .Z(n28882) );
  XNOR U28982 ( .A(n28634), .B(n28916), .Z(n28922) );
  XOR U28983 ( .A(n28630), .B(n28923), .Z(n28920) );
  XNOR U28984 ( .A(n28924), .B(n28912), .Z(n28923) );
  OR U28985 ( .A(n28867), .B(n28875), .Z(n28912) );
  XOR U28986 ( .A(n28630), .B(n28876), .Z(n28875) );
  XNOR U28987 ( .A(n28634), .B(n28925), .Z(n28867) );
  ANDN U28988 ( .B(n28926), .A(n28864), .Z(n28924) );
  XNOR U28989 ( .A(n28927), .B(n28928), .Z(n28897) );
  XOR U28990 ( .A(n28915), .B(n28907), .Z(n28928) );
  XOR U28991 ( .A(n28916), .B(n28929), .Z(n28907) );
  XNOR U28992 ( .A(n28930), .B(n28931), .Z(n28929) );
  NAND U28993 ( .A(n28653), .B(n28861), .Z(n28931) );
  XNOR U28994 ( .A(n28932), .B(n28930), .Z(n28916) );
  NANDN U28995 ( .A(n28878), .B(n28870), .Z(n28930) );
  XOR U28996 ( .A(n28871), .B(n28861), .Z(n28870) );
  XOR U28997 ( .A(n28925), .B(n28400), .Z(n28861) );
  IV U28998 ( .A(n28864), .Z(n28925) );
  XOR U28999 ( .A(n28857), .B(n28933), .Z(n28864) );
  XNOR U29000 ( .A(n28934), .B(n28935), .Z(n28933) );
  XOR U29001 ( .A(n28886), .B(n28653), .Z(n28878) );
  XNOR U29002 ( .A(n28926), .B(n28639), .Z(n28653) );
  IV U29003 ( .A(n28876), .Z(n28926) );
  XOR U29004 ( .A(n28936), .B(n28937), .Z(n28876) );
  XOR U29005 ( .A(n28938), .B(n28939), .Z(n28937) );
  XNOR U29006 ( .A(n28630), .B(n28940), .Z(n28936) );
  ANDN U29007 ( .B(n28871), .A(n28886), .Z(n28932) );
  XNOR U29008 ( .A(n28630), .B(n28941), .Z(n28886) );
  XOR U29009 ( .A(n28634), .B(n28857), .Z(n28871) );
  XOR U29010 ( .A(n28942), .B(n28943), .Z(n28634) );
  XOR U29011 ( .A(n28944), .B(n28939), .Z(n28943) );
  XOR U29012 ( .A(msg[124]), .B(key[124]), .Z(n28939) );
  XOR U29013 ( .A(n28941), .B(n28857), .Z(n28915) );
  IV U29014 ( .A(n28648), .Z(n28941) );
  XNOR U29015 ( .A(n28945), .B(n28919), .Z(n28927) );
  OR U29016 ( .A(n28856), .B(n28646), .Z(n28919) );
  XNOR U29017 ( .A(n28648), .B(n28639), .Z(n28646) );
  XOR U29018 ( .A(n28946), .B(n28942), .Z(n28639) );
  XNOR U29019 ( .A(n28857), .B(n28400), .Z(n28856) );
  XOR U29020 ( .A(n28942), .B(n28947), .Z(n28400) );
  XOR U29021 ( .A(n28934), .B(n28946), .Z(n28947) );
  ANDN U29022 ( .B(n28857), .A(n28648), .Z(n28945) );
  XNOR U29023 ( .A(n28935), .B(n28948), .Z(n28648) );
  XOR U29024 ( .A(n28940), .B(n28946), .Z(n28948) );
  IV U29025 ( .A(n28944), .Z(n28946) );
  XNOR U29026 ( .A(n28934), .B(n28949), .Z(n28940) );
  XNOR U29027 ( .A(msg[123]), .B(key[123]), .Z(n28949) );
  XNOR U29028 ( .A(msg[121]), .B(key[121]), .Z(n28934) );
  XNOR U29029 ( .A(msg[122]), .B(key[122]), .Z(n28935) );
  XOR U29030 ( .A(n28942), .B(n28950), .Z(n28857) );
  XNOR U29031 ( .A(n28944), .B(n28938), .Z(n28950) );
  XNOR U29032 ( .A(msg[127]), .B(key[127]), .Z(n28938) );
  XOR U29033 ( .A(n28630), .B(n28951), .Z(n28944) );
  XNOR U29034 ( .A(msg[126]), .B(key[126]), .Z(n28951) );
  XOR U29035 ( .A(msg[120]), .B(key[120]), .Z(n28630) );
  XNOR U29036 ( .A(msg[125]), .B(key[125]), .Z(n28942) );
  XNOR U29037 ( .A(n26573), .B(n28952), .Z(n22239) );
  XOR U29038 ( .A(n26575), .B(n26576), .Z(n28952) );
  XOR U29039 ( .A(n26609), .B(n28953), .Z(n26576) );
  XOR U29040 ( .A(n28954), .B(n28955), .Z(n28953) );
  ANDN U29041 ( .B(n28956), .A(n26673), .Z(n28954) );
  XNOR U29042 ( .A(n26675), .B(n28957), .Z(n26609) );
  XNOR U29043 ( .A(n28958), .B(n28959), .Z(n28957) );
  NAND U29044 ( .A(n28960), .B(n26695), .Z(n28959) );
  XNOR U29045 ( .A(n26691), .B(n28961), .Z(n26575) );
  XNOR U29046 ( .A(n26688), .B(n28962), .Z(n28961) );
  NANDN U29047 ( .A(n26679), .B(n28963), .Z(n28962) );
  OR U29048 ( .A(n28964), .B(n26680), .Z(n26688) );
  XOR U29049 ( .A(n26614), .B(n28965), .Z(n26680) );
  XNOR U29050 ( .A(n26702), .B(n26564), .Z(n26573) );
  XNOR U29051 ( .A(n26675), .B(n28966), .Z(n26564) );
  XNOR U29052 ( .A(n28955), .B(n28967), .Z(n28966) );
  NANDN U29053 ( .A(n28968), .B(n28969), .Z(n28967) );
  OR U29054 ( .A(n28970), .B(n28971), .Z(n28955) );
  XOR U29055 ( .A(n28972), .B(n28958), .Z(n26675) );
  NANDN U29056 ( .A(n28973), .B(n28974), .Z(n28958) );
  AND U29057 ( .A(n28975), .B(n28976), .Z(n28972) );
  XNOR U29058 ( .A(n26691), .B(n28977), .Z(n26702) );
  XOR U29059 ( .A(n28978), .B(n26671), .Z(n28977) );
  OR U29060 ( .A(n28979), .B(n28970), .Z(n26671) );
  XNOR U29061 ( .A(n26673), .B(n28968), .Z(n28970) );
  NOR U29062 ( .A(n28980), .B(n28968), .Z(n28978) );
  XOR U29063 ( .A(n28981), .B(n26693), .Z(n26691) );
  OR U29064 ( .A(n28973), .B(n28982), .Z(n26693) );
  XNOR U29065 ( .A(n28975), .B(n26695), .Z(n28973) );
  XOR U29066 ( .A(n28968), .B(n26679), .Z(n26695) );
  IV U29067 ( .A(n28965), .Z(n26679) );
  XOR U29068 ( .A(n28983), .B(n28984), .Z(n28965) );
  NANDN U29069 ( .A(n28985), .B(n28986), .Z(n28984) );
  XNOR U29070 ( .A(n28987), .B(n28988), .Z(n28968) );
  OR U29071 ( .A(n28985), .B(n28989), .Z(n28988) );
  ANDN U29072 ( .B(n28975), .A(n28990), .Z(n28981) );
  XOR U29073 ( .A(n26673), .B(n26614), .Z(n28975) );
  XNOR U29074 ( .A(n28983), .B(n28991), .Z(n26614) );
  NANDN U29075 ( .A(n28992), .B(n28993), .Z(n28991) );
  NANDN U29076 ( .A(n28994), .B(n28995), .Z(n28983) );
  OR U29077 ( .A(n28997), .B(n28994), .Z(n28987) );
  XOR U29078 ( .A(n28998), .B(n28985), .Z(n28994) );
  XNOR U29079 ( .A(n28999), .B(n29000), .Z(n28985) );
  XOR U29080 ( .A(n29001), .B(n28993), .Z(n29000) );
  XNOR U29081 ( .A(n29002), .B(n29003), .Z(n28999) );
  XNOR U29082 ( .A(n29004), .B(n29005), .Z(n29003) );
  ANDN U29083 ( .B(n28993), .A(n29006), .Z(n29004) );
  IV U29084 ( .A(n29007), .Z(n28993) );
  ANDN U29085 ( .B(n28998), .A(n29006), .Z(n28996) );
  IV U29086 ( .A(n28992), .Z(n28998) );
  XNOR U29087 ( .A(n29001), .B(n29008), .Z(n28992) );
  XNOR U29088 ( .A(n29005), .B(n29009), .Z(n29008) );
  NANDN U29089 ( .A(n28989), .B(n28986), .Z(n29009) );
  NANDN U29090 ( .A(n28997), .B(n28995), .Z(n29005) );
  XNOR U29091 ( .A(n28986), .B(n29007), .Z(n28995) );
  XOR U29092 ( .A(n29010), .B(n29011), .Z(n29007) );
  XOR U29093 ( .A(n29012), .B(n29013), .Z(n29011) );
  XNOR U29094 ( .A(n28969), .B(n29014), .Z(n29013) );
  XNOR U29095 ( .A(n29015), .B(n29016), .Z(n29010) );
  XNOR U29096 ( .A(n29017), .B(n29018), .Z(n29016) );
  ANDN U29097 ( .B(n28956), .A(n26674), .Z(n29017) );
  XNOR U29098 ( .A(n29006), .B(n28989), .Z(n28997) );
  IV U29099 ( .A(n29002), .Z(n29006) );
  XOR U29100 ( .A(n29019), .B(n29020), .Z(n29002) );
  XNOR U29101 ( .A(n29021), .B(n29014), .Z(n29020) );
  XOR U29102 ( .A(n29022), .B(n29023), .Z(n29014) );
  XNOR U29103 ( .A(n29024), .B(n29025), .Z(n29023) );
  NAND U29104 ( .A(n26696), .B(n28960), .Z(n29025) );
  XNOR U29105 ( .A(n29026), .B(n29027), .Z(n29019) );
  ANDN U29106 ( .B(n29028), .A(n26690), .Z(n29026) );
  XOR U29107 ( .A(n28989), .B(n28986), .Z(n29001) );
  XNOR U29108 ( .A(n29029), .B(n29030), .Z(n28986) );
  XNOR U29109 ( .A(n29022), .B(n29031), .Z(n29030) );
  XNOR U29110 ( .A(n29021), .B(n28956), .Z(n29031) );
  XNOR U29111 ( .A(n29032), .B(n29033), .Z(n29029) );
  XNOR U29112 ( .A(n29034), .B(n29018), .Z(n29033) );
  OR U29113 ( .A(n28971), .B(n28979), .Z(n29018) );
  XNOR U29114 ( .A(n29032), .B(n29015), .Z(n28979) );
  XNOR U29115 ( .A(n28956), .B(n28969), .Z(n28971) );
  ANDN U29116 ( .B(n28969), .A(n28980), .Z(n29034) );
  XOR U29117 ( .A(n29035), .B(n29036), .Z(n28989) );
  XOR U29118 ( .A(n29022), .B(n29012), .Z(n29036) );
  XNOR U29119 ( .A(n28963), .B(n26678), .Z(n29012) );
  XOR U29120 ( .A(n29037), .B(n29024), .Z(n29022) );
  NANDN U29121 ( .A(n28982), .B(n28974), .Z(n29024) );
  XOR U29122 ( .A(n28976), .B(n28960), .Z(n28974) );
  XOR U29123 ( .A(n26678), .B(n28969), .Z(n28960) );
  XNOR U29124 ( .A(n29028), .B(n29038), .Z(n28969) );
  XOR U29125 ( .A(n29039), .B(n29040), .Z(n29038) );
  XOR U29126 ( .A(n28990), .B(n26696), .Z(n28982) );
  XNOR U29127 ( .A(n28980), .B(n28963), .Z(n26696) );
  IV U29128 ( .A(n29015), .Z(n28980) );
  XOR U29129 ( .A(n29041), .B(n29042), .Z(n29015) );
  XOR U29130 ( .A(n29043), .B(n29044), .Z(n29042) );
  XOR U29131 ( .A(n29032), .B(n29045), .Z(n29041) );
  ANDN U29132 ( .B(n28976), .A(n28990), .Z(n29037) );
  XNOR U29133 ( .A(n29032), .B(n29046), .Z(n28990) );
  XOR U29134 ( .A(n29028), .B(n28956), .Z(n28976) );
  XNOR U29135 ( .A(n29047), .B(n29048), .Z(n28956) );
  XOR U29136 ( .A(n29049), .B(n29044), .Z(n29048) );
  XNOR U29137 ( .A(n29050), .B(n29051), .Z(n29044) );
  XOR U29138 ( .A(n25517), .B(n26449), .Z(n29051) );
  XNOR U29139 ( .A(n29052), .B(n29053), .Z(n26449) );
  XOR U29140 ( .A(n24495), .B(n25535), .Z(n29053) );
  IV U29141 ( .A(n26439), .Z(n25535) );
  XOR U29142 ( .A(n29054), .B(n29055), .Z(n26439) );
  XNOR U29143 ( .A(n29056), .B(n29057), .Z(n29055) );
  XNOR U29144 ( .A(n29058), .B(n29059), .Z(n29054) );
  XOR U29145 ( .A(n29060), .B(n29061), .Z(n29059) );
  ANDN U29146 ( .B(n29062), .A(n29063), .Z(n29061) );
  XOR U29147 ( .A(n29064), .B(n24466), .Z(n24495) );
  XOR U29148 ( .A(n29065), .B(n25519), .Z(n29052) );
  XNOR U29149 ( .A(n29066), .B(n25562), .Z(n25517) );
  XNOR U29150 ( .A(key[140]), .B(n24493), .Z(n29050) );
  XOR U29151 ( .A(n24488), .B(n25534), .Z(n24493) );
  XOR U29152 ( .A(n29021), .B(n29067), .Z(n29035) );
  XNOR U29153 ( .A(n29068), .B(n29027), .Z(n29067) );
  OR U29154 ( .A(n26681), .B(n28964), .Z(n29027) );
  XNOR U29155 ( .A(n29046), .B(n28963), .Z(n28964) );
  XNOR U29156 ( .A(n29028), .B(n26678), .Z(n26681) );
  IV U29157 ( .A(n26613), .Z(n29028) );
  AND U29158 ( .A(n26678), .B(n28963), .Z(n29068) );
  XOR U29159 ( .A(n29049), .B(n29047), .Z(n28963) );
  XNOR U29160 ( .A(n29047), .B(n29069), .Z(n26678) );
  XNOR U29161 ( .A(n29040), .B(n29070), .Z(n29069) );
  XNOR U29162 ( .A(n26690), .B(n26613), .Z(n29021) );
  XOR U29163 ( .A(n29047), .B(n29071), .Z(n26613) );
  XNOR U29164 ( .A(n29049), .B(n29043), .Z(n29071) );
  XOR U29165 ( .A(n29072), .B(n29073), .Z(n29043) );
  XNOR U29166 ( .A(n25546), .B(n26446), .Z(n29073) );
  XOR U29167 ( .A(n25554), .B(n25529), .Z(n26446) );
  XOR U29168 ( .A(n29074), .B(n29075), .Z(n25554) );
  XOR U29169 ( .A(n29076), .B(n29077), .Z(n29075) );
  XOR U29170 ( .A(n29065), .B(n24488), .Z(n25546) );
  XOR U29171 ( .A(key[143]), .B(n25531), .Z(n29072) );
  XNOR U29172 ( .A(n29078), .B(n29079), .Z(n25531) );
  XNOR U29173 ( .A(n29080), .B(n29081), .Z(n29079) );
  XOR U29174 ( .A(n29082), .B(n29083), .Z(n29078) );
  XNOR U29175 ( .A(n29084), .B(n29085), .Z(n29047) );
  XNOR U29176 ( .A(n25550), .B(n26440), .Z(n29085) );
  XNOR U29177 ( .A(n25534), .B(n24481), .Z(n26440) );
  XOR U29178 ( .A(n29086), .B(n29087), .Z(n24481) );
  XNOR U29179 ( .A(n29064), .B(n29077), .Z(n29087) );
  XNOR U29180 ( .A(n29088), .B(n29089), .Z(n29077) );
  XNOR U29181 ( .A(n29090), .B(n29091), .Z(n29089) );
  NANDN U29182 ( .A(n29092), .B(n29093), .Z(n29091) );
  XOR U29183 ( .A(n29094), .B(n29095), .Z(n29086) );
  XOR U29184 ( .A(n29096), .B(n29097), .Z(n29095) );
  ANDN U29185 ( .B(n29098), .A(n29099), .Z(n29097) );
  XNOR U29186 ( .A(n29100), .B(n29101), .Z(n25534) );
  XOR U29187 ( .A(n29102), .B(n29103), .Z(n29101) );
  XOR U29188 ( .A(n29104), .B(n29105), .Z(n29100) );
  XOR U29189 ( .A(n29106), .B(n29107), .Z(n29105) );
  ANDN U29190 ( .B(n29108), .A(n29109), .Z(n29107) );
  XOR U29191 ( .A(n25536), .B(n29110), .Z(n29084) );
  XNOR U29192 ( .A(key[141]), .B(n26435), .Z(n29110) );
  XOR U29193 ( .A(n29111), .B(n29112), .Z(n26435) );
  XNOR U29194 ( .A(n29113), .B(n29114), .Z(n25536) );
  XNOR U29195 ( .A(n29115), .B(n29081), .Z(n29114) );
  XNOR U29196 ( .A(n29116), .B(n29117), .Z(n29081) );
  XNOR U29197 ( .A(n29118), .B(n29119), .Z(n29117) );
  OR U29198 ( .A(n29120), .B(n29121), .Z(n29119) );
  XNOR U29199 ( .A(n29066), .B(n29122), .Z(n29113) );
  XOR U29200 ( .A(n29123), .B(n29124), .Z(n29122) );
  ANDN U29201 ( .B(n29125), .A(n29126), .Z(n29124) );
  IV U29202 ( .A(n29046), .Z(n26690) );
  XOR U29203 ( .A(n29070), .B(n29127), .Z(n29046) );
  XNOR U29204 ( .A(n29039), .B(n29045), .Z(n29127) );
  XOR U29205 ( .A(n29128), .B(n29129), .Z(n29045) );
  XOR U29206 ( .A(n29040), .B(n29130), .Z(n29129) );
  XNOR U29207 ( .A(n24464), .B(n26452), .Z(n29130) );
  XOR U29208 ( .A(n24513), .B(n25516), .Z(n26452) );
  XNOR U29209 ( .A(n29058), .B(n26425), .Z(n25516) );
  IV U29210 ( .A(n26457), .Z(n24464) );
  XOR U29211 ( .A(n24506), .B(n25559), .Z(n26457) );
  XNOR U29212 ( .A(n29074), .B(n29131), .Z(n24506) );
  XOR U29213 ( .A(n29132), .B(n29133), .Z(n29131) );
  XOR U29214 ( .A(n29134), .B(n29135), .Z(n29074) );
  XNOR U29215 ( .A(n29136), .B(n29137), .Z(n29040) );
  XNOR U29216 ( .A(n26462), .B(n26425), .Z(n29137) );
  XNOR U29217 ( .A(n29138), .B(n29139), .Z(n26425) );
  IV U29218 ( .A(n25545), .Z(n26462) );
  XNOR U29219 ( .A(n29082), .B(n29083), .Z(n29140) );
  XNOR U29220 ( .A(n25571), .B(n29141), .Z(n29136) );
  XNOR U29221 ( .A(key[137]), .B(n24511), .Z(n29141) );
  XOR U29222 ( .A(n25549), .B(n25564), .Z(n24511) );
  IV U29223 ( .A(n24505), .Z(n25549) );
  XNOR U29224 ( .A(n29076), .B(n29142), .Z(n24505) );
  XNOR U29225 ( .A(n29134), .B(n29135), .Z(n29142) );
  XNOR U29226 ( .A(n29144), .B(n29145), .Z(n29143) );
  NANDN U29227 ( .A(n29092), .B(n29146), .Z(n29145) );
  XOR U29228 ( .A(n25569), .B(n29148), .Z(n29128) );
  XNOR U29229 ( .A(key[139]), .B(n24508), .Z(n29148) );
  XOR U29230 ( .A(n24488), .B(n25519), .Z(n24508) );
  XNOR U29231 ( .A(n29102), .B(n25571), .Z(n25519) );
  XNOR U29232 ( .A(n29149), .B(n29150), .Z(n25569) );
  XNOR U29233 ( .A(n29080), .B(n29151), .Z(n29150) );
  XOR U29234 ( .A(n29082), .B(n29152), .Z(n29149) );
  XNOR U29235 ( .A(n29154), .B(n29155), .Z(n29153) );
  OR U29236 ( .A(n29120), .B(n29156), .Z(n29155) );
  XOR U29237 ( .A(n29158), .B(n29159), .Z(n29039) );
  XOR U29238 ( .A(n25559), .B(n25562), .Z(n29159) );
  XNOR U29239 ( .A(n29160), .B(n29080), .Z(n25562) );
  XOR U29240 ( .A(n29161), .B(n29162), .Z(n29080) );
  XNOR U29241 ( .A(n29163), .B(n29164), .Z(n29162) );
  NANDN U29242 ( .A(n29165), .B(n29166), .Z(n29164) );
  XNOR U29243 ( .A(n29167), .B(n29168), .Z(n25559) );
  XOR U29244 ( .A(n29169), .B(n29170), .Z(n29168) );
  XNOR U29245 ( .A(n29171), .B(n29172), .Z(n29167) );
  XNOR U29246 ( .A(n26426), .B(n29173), .Z(n29158) );
  XOR U29247 ( .A(key[138]), .B(n24504), .Z(n29173) );
  XNOR U29248 ( .A(n29134), .B(n29174), .Z(n24466) );
  XNOR U29249 ( .A(n29175), .B(n29176), .Z(n29134) );
  XNOR U29250 ( .A(n29177), .B(n29178), .Z(n29176) );
  NANDN U29251 ( .A(n29179), .B(n29180), .Z(n29178) );
  XNOR U29252 ( .A(n29181), .B(n29182), .Z(n25571) );
  XOR U29253 ( .A(n29183), .B(n29184), .Z(n26426) );
  XNOR U29254 ( .A(n29139), .B(n29112), .Z(n29184) );
  XNOR U29255 ( .A(n29185), .B(n29186), .Z(n29112) );
  XNOR U29256 ( .A(n29187), .B(n29060), .Z(n29186) );
  NOR U29257 ( .A(n29188), .B(n29189), .Z(n29060) );
  ANDN U29258 ( .B(n29190), .A(n29191), .Z(n29187) );
  IV U29259 ( .A(n29192), .Z(n29139) );
  XOR U29260 ( .A(n29193), .B(n29194), .Z(n29183) );
  IV U29261 ( .A(n29049), .Z(n29070) );
  XOR U29262 ( .A(n29195), .B(n29196), .Z(n29049) );
  XNOR U29263 ( .A(n26433), .B(n26674), .Z(n29196) );
  IV U29264 ( .A(n29032), .Z(n26674) );
  XOR U29265 ( .A(n29197), .B(n29198), .Z(n29032) );
  XOR U29266 ( .A(n24488), .B(n26461), .Z(n29198) );
  IV U29267 ( .A(n26456), .Z(n26461) );
  XOR U29268 ( .A(n29192), .B(n29199), .Z(n26456) );
  XNOR U29269 ( .A(n29193), .B(n29111), .Z(n29199) );
  XOR U29270 ( .A(n24512), .B(n29200), .Z(n29197) );
  XOR U29271 ( .A(key[136]), .B(n25564), .Z(n29200) );
  XNOR U29272 ( .A(n29201), .B(n29202), .Z(n25564) );
  XOR U29273 ( .A(n29171), .B(n29172), .Z(n29202) );
  XOR U29274 ( .A(n26436), .B(n25553), .Z(n24512) );
  XOR U29275 ( .A(n29174), .B(n29064), .Z(n25553) );
  XNOR U29276 ( .A(n29088), .B(n29203), .Z(n29064) );
  XOR U29277 ( .A(n29204), .B(n29177), .Z(n29203) );
  OR U29278 ( .A(n29205), .B(n29206), .Z(n29177) );
  ANDN U29279 ( .B(n29207), .A(n29208), .Z(n29204) );
  XOR U29280 ( .A(n29175), .B(n29209), .Z(n29088) );
  XNOR U29281 ( .A(n29210), .B(n29211), .Z(n29209) );
  NAND U29282 ( .A(n29212), .B(n29213), .Z(n29211) );
  XOR U29283 ( .A(n29066), .B(n29160), .Z(n26436) );
  IV U29284 ( .A(n29214), .Z(n29160) );
  XNOR U29285 ( .A(n29116), .B(n29215), .Z(n29066) );
  XOR U29286 ( .A(n29216), .B(n29163), .Z(n29215) );
  OR U29287 ( .A(n29217), .B(n29218), .Z(n29163) );
  XOR U29288 ( .A(n29161), .B(n29221), .Z(n29116) );
  XNOR U29289 ( .A(n29222), .B(n29223), .Z(n29221) );
  NANDN U29290 ( .A(n29224), .B(n29225), .Z(n29223) );
  XNOR U29291 ( .A(n24480), .B(n26445), .Z(n26433) );
  XOR U29292 ( .A(n29065), .B(n25530), .Z(n26445) );
  XNOR U29293 ( .A(n29226), .B(n29227), .Z(n25530) );
  XOR U29294 ( .A(n29192), .B(n29057), .Z(n29227) );
  XNOR U29295 ( .A(n29228), .B(n29229), .Z(n29057) );
  XNOR U29296 ( .A(n29230), .B(n29231), .Z(n29229) );
  OR U29297 ( .A(n29232), .B(n29233), .Z(n29231) );
  XOR U29298 ( .A(n29234), .B(n29235), .Z(n29192) );
  XNOR U29299 ( .A(n29236), .B(n29237), .Z(n29235) );
  NANDN U29300 ( .A(n29238), .B(n29239), .Z(n29237) );
  XOR U29301 ( .A(n29193), .B(n29111), .Z(n29226) );
  XOR U29302 ( .A(n29138), .B(n29194), .Z(n29111) );
  XOR U29303 ( .A(n29056), .B(n29240), .Z(n29194) );
  XNOR U29304 ( .A(n29241), .B(n29242), .Z(n29240) );
  NANDN U29305 ( .A(n29243), .B(n29244), .Z(n29242) );
  XNOR U29306 ( .A(n29241), .B(n29246), .Z(n29245) );
  OR U29307 ( .A(n29232), .B(n29247), .Z(n29246) );
  OR U29308 ( .A(n29248), .B(n29249), .Z(n29241) );
  XNOR U29309 ( .A(n29056), .B(n29250), .Z(n29185) );
  XNOR U29310 ( .A(n29251), .B(n29252), .Z(n29250) );
  OR U29311 ( .A(n29253), .B(n29254), .Z(n29252) );
  XOR U29312 ( .A(n29255), .B(n29251), .Z(n29056) );
  NANDN U29313 ( .A(n29256), .B(n29257), .Z(n29251) );
  ANDN U29314 ( .B(n29258), .A(n29259), .Z(n29255) );
  IV U29315 ( .A(n24513), .Z(n29065) );
  XOR U29316 ( .A(n29058), .B(n29138), .Z(n24513) );
  XOR U29317 ( .A(n29234), .B(n29260), .Z(n29138) );
  XOR U29318 ( .A(n29261), .B(n29230), .Z(n29260) );
  OR U29319 ( .A(n29262), .B(n29248), .Z(n29230) );
  XOR U29320 ( .A(n29232), .B(n29263), .Z(n29248) );
  ANDN U29321 ( .B(n29264), .A(n29243), .Z(n29261) );
  XNOR U29322 ( .A(n29228), .B(n29265), .Z(n29058) );
  XOR U29323 ( .A(n29266), .B(n29236), .Z(n29265) );
  OR U29324 ( .A(n29267), .B(n29188), .Z(n29236) );
  XNOR U29325 ( .A(n29190), .B(n29239), .Z(n29188) );
  XNOR U29326 ( .A(n29234), .B(n29269), .Z(n29228) );
  XNOR U29327 ( .A(n29270), .B(n29271), .Z(n29269) );
  NANDN U29328 ( .A(n29253), .B(n29272), .Z(n29271) );
  XOR U29329 ( .A(n29273), .B(n29270), .Z(n29234) );
  OR U29330 ( .A(n29256), .B(n29274), .Z(n29270) );
  XOR U29331 ( .A(n29275), .B(n29253), .Z(n29256) );
  XOR U29332 ( .A(n29263), .B(n29063), .Z(n29253) );
  IV U29333 ( .A(n29239), .Z(n29063) );
  XOR U29334 ( .A(n29276), .B(n29277), .Z(n29239) );
  NANDN U29335 ( .A(n29278), .B(n29279), .Z(n29277) );
  IV U29336 ( .A(n29243), .Z(n29263) );
  XNOR U29337 ( .A(n29280), .B(n29281), .Z(n29243) );
  NANDN U29338 ( .A(n29278), .B(n29282), .Z(n29281) );
  ANDN U29339 ( .B(n29275), .A(n29283), .Z(n29273) );
  IV U29340 ( .A(n29259), .Z(n29275) );
  XOR U29341 ( .A(n29190), .B(n29232), .Z(n29259) );
  XOR U29342 ( .A(n29284), .B(n29280), .Z(n29232) );
  NANDN U29343 ( .A(n29285), .B(n29286), .Z(n29280) );
  NANDN U29344 ( .A(n29285), .B(n29290), .Z(n29276) );
  XOR U29345 ( .A(n29291), .B(n29292), .Z(n29278) );
  XOR U29346 ( .A(n29293), .B(n29288), .Z(n29292) );
  XNOR U29347 ( .A(n29294), .B(n29295), .Z(n29291) );
  XNOR U29348 ( .A(n29296), .B(n29297), .Z(n29295) );
  ANDN U29349 ( .B(n29293), .A(n29288), .Z(n29296) );
  ANDN U29350 ( .B(n29293), .A(n29287), .Z(n29289) );
  XNOR U29351 ( .A(n29294), .B(n29298), .Z(n29287) );
  XOR U29352 ( .A(n29299), .B(n29297), .Z(n29298) );
  NAND U29353 ( .A(n29286), .B(n29290), .Z(n29297) );
  XNOR U29354 ( .A(n29282), .B(n29288), .Z(n29286) );
  XOR U29355 ( .A(n29300), .B(n29301), .Z(n29288) );
  XOR U29356 ( .A(n29302), .B(n29303), .Z(n29301) );
  XNOR U29357 ( .A(n29304), .B(n29305), .Z(n29300) );
  ANDN U29358 ( .B(n29268), .A(n29191), .Z(n29304) );
  AND U29359 ( .A(n29279), .B(n29282), .Z(n29299) );
  XNOR U29360 ( .A(n29279), .B(n29282), .Z(n29294) );
  XNOR U29361 ( .A(n29306), .B(n29307), .Z(n29282) );
  XNOR U29362 ( .A(n29308), .B(n29309), .Z(n29307) );
  XOR U29363 ( .A(n29302), .B(n29310), .Z(n29306) );
  XNOR U29364 ( .A(n29311), .B(n29305), .Z(n29310) );
  OR U29365 ( .A(n29189), .B(n29267), .Z(n29305) );
  XNOR U29366 ( .A(n29312), .B(n29238), .Z(n29267) );
  XNOR U29367 ( .A(n29191), .B(n29313), .Z(n29189) );
  NOR U29368 ( .A(n29313), .B(n29238), .Z(n29311) );
  XNOR U29369 ( .A(n29314), .B(n29315), .Z(n29279) );
  XNOR U29370 ( .A(n29316), .B(n29317), .Z(n29315) );
  XOR U29371 ( .A(n29247), .B(n29302), .Z(n29317) );
  XOR U29372 ( .A(n29268), .B(n29318), .Z(n29302) );
  XNOR U29373 ( .A(n29233), .B(n29319), .Z(n29314) );
  XNOR U29374 ( .A(n29320), .B(n29321), .Z(n29319) );
  ANDN U29375 ( .B(n29244), .A(n29322), .Z(n29320) );
  XNOR U29376 ( .A(n29323), .B(n29324), .Z(n29293) );
  XNOR U29377 ( .A(n29303), .B(n29325), .Z(n29324) );
  XNOR U29378 ( .A(n29244), .B(n29309), .Z(n29325) );
  XOR U29379 ( .A(n29238), .B(n29313), .Z(n29309) );
  XNOR U29380 ( .A(n29316), .B(n29326), .Z(n29303) );
  XNOR U29381 ( .A(n29327), .B(n29328), .Z(n29326) );
  NANDN U29382 ( .A(n29254), .B(n29272), .Z(n29328) );
  IV U29383 ( .A(n29308), .Z(n29316) );
  XNOR U29384 ( .A(n29329), .B(n29327), .Z(n29308) );
  NANDN U29385 ( .A(n29274), .B(n29257), .Z(n29327) );
  XOR U29386 ( .A(n29244), .B(n29313), .Z(n29254) );
  IV U29387 ( .A(n29062), .Z(n29313) );
  XOR U29388 ( .A(n29330), .B(n29331), .Z(n29062) );
  XNOR U29389 ( .A(n29332), .B(n29333), .Z(n29331) );
  XOR U29390 ( .A(n29283), .B(n29272), .Z(n29274) );
  XNOR U29391 ( .A(n29264), .B(n29238), .Z(n29272) );
  XNOR U29392 ( .A(n29333), .B(n29330), .Z(n29238) );
  ANDN U29393 ( .B(n29258), .A(n29283), .Z(n29329) );
  XNOR U29394 ( .A(n29334), .B(n29268), .Z(n29283) );
  IV U29395 ( .A(n29312), .Z(n29268) );
  XNOR U29396 ( .A(n29335), .B(n29336), .Z(n29312) );
  XNOR U29397 ( .A(n29337), .B(n29333), .Z(n29336) );
  XOR U29398 ( .A(n29338), .B(n29318), .Z(n29258) );
  XNOR U29399 ( .A(n29322), .B(n29339), .Z(n29323) );
  XNOR U29400 ( .A(n29340), .B(n29321), .Z(n29339) );
  OR U29401 ( .A(n29249), .B(n29262), .Z(n29321) );
  XOR U29402 ( .A(n29233), .B(n29264), .Z(n29262) );
  IV U29403 ( .A(n29322), .Z(n29264) );
  XOR U29404 ( .A(n29247), .B(n29244), .Z(n29249) );
  XNOR U29405 ( .A(n29318), .B(n29341), .Z(n29244) );
  XNOR U29406 ( .A(n29332), .B(n29335), .Z(n29341) );
  XNOR U29407 ( .A(msg[74]), .B(key[74]), .Z(n29335) );
  IV U29408 ( .A(n29191), .Z(n29318) );
  XOR U29409 ( .A(n29342), .B(n29343), .Z(n29191) );
  XOR U29410 ( .A(n29333), .B(n29344), .Z(n29343) );
  IV U29411 ( .A(n29338), .Z(n29247) );
  ANDN U29412 ( .B(n29338), .A(n29233), .Z(n29340) );
  XOR U29413 ( .A(n29330), .B(n29345), .Z(n29338) );
  XNOR U29414 ( .A(n29333), .B(n29346), .Z(n29345) );
  XOR U29415 ( .A(n29334), .B(n29347), .Z(n29333) );
  XNOR U29416 ( .A(msg[78]), .B(key[78]), .Z(n29347) );
  IV U29417 ( .A(n29342), .Z(n29330) );
  XOR U29418 ( .A(msg[77]), .B(key[77]), .Z(n29342) );
  XOR U29419 ( .A(n29348), .B(n29349), .Z(n29322) );
  XOR U29420 ( .A(n29346), .B(n29344), .Z(n29349) );
  XOR U29421 ( .A(msg[79]), .B(key[79]), .Z(n29344) );
  XNOR U29422 ( .A(msg[76]), .B(key[76]), .Z(n29346) );
  XOR U29423 ( .A(n29233), .B(n29337), .Z(n29348) );
  XNOR U29424 ( .A(n29332), .B(n29350), .Z(n29337) );
  XNOR U29425 ( .A(msg[75]), .B(key[75]), .Z(n29350) );
  XNOR U29426 ( .A(msg[73]), .B(key[73]), .Z(n29332) );
  IV U29427 ( .A(n29334), .Z(n29233) );
  XOR U29428 ( .A(msg[72]), .B(key[72]), .Z(n29334) );
  XNOR U29429 ( .A(n24473), .B(n25550), .Z(n24480) );
  XNOR U29430 ( .A(n29351), .B(n29352), .Z(n29170) );
  XNOR U29431 ( .A(n29353), .B(n29106), .Z(n29352) );
  NOR U29432 ( .A(n29354), .B(n29355), .Z(n29106) );
  ANDN U29433 ( .B(n29356), .A(n29357), .Z(n29353) );
  XNOR U29434 ( .A(n29076), .B(n29133), .Z(n24473) );
  XNOR U29435 ( .A(n29147), .B(n29358), .Z(n29133) );
  XNOR U29436 ( .A(n29359), .B(n29096), .Z(n29358) );
  NOR U29437 ( .A(n29206), .B(n29360), .Z(n29096) );
  XNOR U29438 ( .A(n29207), .B(n29180), .Z(n29206) );
  ANDN U29439 ( .B(n29207), .A(n29361), .Z(n29359) );
  XOR U29440 ( .A(n29094), .B(n29362), .Z(n29147) );
  XNOR U29441 ( .A(n29363), .B(n29364), .Z(n29362) );
  NAND U29442 ( .A(n29212), .B(n29365), .Z(n29364) );
  XNOR U29443 ( .A(n29174), .B(n29132), .Z(n29076) );
  XNOR U29444 ( .A(n29094), .B(n29366), .Z(n29132) );
  XNOR U29445 ( .A(n29144), .B(n29367), .Z(n29366) );
  OR U29446 ( .A(n29368), .B(n29369), .Z(n29367) );
  OR U29447 ( .A(n29370), .B(n29371), .Z(n29144) );
  XNOR U29448 ( .A(n29372), .B(n29363), .Z(n29094) );
  NANDN U29449 ( .A(n29373), .B(n29374), .Z(n29363) );
  ANDN U29450 ( .B(n29375), .A(n29376), .Z(n29372) );
  XOR U29451 ( .A(n29378), .B(n29090), .Z(n29377) );
  OR U29452 ( .A(n29370), .B(n29379), .Z(n29090) );
  XNOR U29453 ( .A(n29092), .B(n29368), .Z(n29370) );
  NOR U29454 ( .A(n29380), .B(n29368), .Z(n29378) );
  XNOR U29455 ( .A(n29381), .B(n29210), .Z(n29175) );
  OR U29456 ( .A(n29373), .B(n29382), .Z(n29210) );
  XNOR U29457 ( .A(n29383), .B(n29212), .Z(n29373) );
  XNOR U29458 ( .A(n29368), .B(n29180), .Z(n29212) );
  IV U29459 ( .A(n29099), .Z(n29180) );
  XNOR U29460 ( .A(n29384), .B(n29385), .Z(n29099) );
  NANDN U29461 ( .A(n29386), .B(n29387), .Z(n29385) );
  XNOR U29462 ( .A(n29388), .B(n29389), .Z(n29368) );
  NANDN U29463 ( .A(n29386), .B(n29390), .Z(n29389) );
  ANDN U29464 ( .B(n29383), .A(n29391), .Z(n29381) );
  IV U29465 ( .A(n29376), .Z(n29383) );
  XOR U29466 ( .A(n29092), .B(n29207), .Z(n29376) );
  XNOR U29467 ( .A(n29392), .B(n29384), .Z(n29207) );
  NANDN U29468 ( .A(n29393), .B(n29394), .Z(n29384) );
  XOR U29469 ( .A(n29387), .B(n29395), .Z(n29394) );
  ANDN U29470 ( .B(n29395), .A(n29396), .Z(n29392) );
  NANDN U29471 ( .A(n29393), .B(n29398), .Z(n29388) );
  XOR U29472 ( .A(n29399), .B(n29400), .Z(n29386) );
  XOR U29473 ( .A(n29401), .B(n29402), .Z(n29400) );
  XNOR U29474 ( .A(n29403), .B(n29404), .Z(n29399) );
  XNOR U29475 ( .A(n29405), .B(n29406), .Z(n29404) );
  ANDN U29476 ( .B(n29402), .A(n29401), .Z(n29405) );
  ANDN U29477 ( .B(n29402), .A(n29396), .Z(n29397) );
  XNOR U29478 ( .A(n29403), .B(n29407), .Z(n29396) );
  XOR U29479 ( .A(n29408), .B(n29406), .Z(n29407) );
  NAND U29480 ( .A(n29398), .B(n29409), .Z(n29406) );
  XNOR U29481 ( .A(n29387), .B(n29401), .Z(n29409) );
  IV U29482 ( .A(n29395), .Z(n29401) );
  XNOR U29483 ( .A(n29410), .B(n29411), .Z(n29395) );
  XNOR U29484 ( .A(n29412), .B(n29413), .Z(n29411) );
  XOR U29485 ( .A(n29369), .B(n29414), .Z(n29413) );
  XNOR U29486 ( .A(n29380), .B(n29415), .Z(n29410) );
  XNOR U29487 ( .A(n29416), .B(n29417), .Z(n29415) );
  AND U29488 ( .A(n29146), .B(n29093), .Z(n29416) );
  XOR U29489 ( .A(n29390), .B(n29402), .Z(n29398) );
  AND U29490 ( .A(n29387), .B(n29390), .Z(n29408) );
  XNOR U29491 ( .A(n29387), .B(n29390), .Z(n29403) );
  XNOR U29492 ( .A(n29418), .B(n29419), .Z(n29390) );
  XNOR U29493 ( .A(n29420), .B(n29414), .Z(n29419) );
  XOR U29494 ( .A(n29421), .B(n29422), .Z(n29418) );
  XNOR U29495 ( .A(n29423), .B(n29424), .Z(n29422) );
  ANDN U29496 ( .B(n29098), .A(n29179), .Z(n29423) );
  XNOR U29497 ( .A(n29425), .B(n29426), .Z(n29387) );
  XNOR U29498 ( .A(n29146), .B(n29421), .Z(n29427) );
  XOR U29499 ( .A(n29093), .B(n29428), .Z(n29425) );
  XNOR U29500 ( .A(n29429), .B(n29417), .Z(n29428) );
  OR U29501 ( .A(n29371), .B(n29379), .Z(n29417) );
  XOR U29502 ( .A(n29093), .B(n29380), .Z(n29379) );
  XNOR U29503 ( .A(n29146), .B(n29430), .Z(n29371) );
  ANDN U29504 ( .B(n29431), .A(n29369), .Z(n29429) );
  XNOR U29505 ( .A(n29432), .B(n29433), .Z(n29402) );
  XOR U29506 ( .A(n29420), .B(n29412), .Z(n29433) );
  XOR U29507 ( .A(n29421), .B(n29434), .Z(n29412) );
  XNOR U29508 ( .A(n29435), .B(n29436), .Z(n29434) );
  NAND U29509 ( .A(n29213), .B(n29365), .Z(n29436) );
  XNOR U29510 ( .A(n29437), .B(n29435), .Z(n29421) );
  NANDN U29511 ( .A(n29382), .B(n29374), .Z(n29435) );
  XOR U29512 ( .A(n29375), .B(n29365), .Z(n29374) );
  XOR U29513 ( .A(n29430), .B(n29098), .Z(n29365) );
  IV U29514 ( .A(n29369), .Z(n29430) );
  XOR U29515 ( .A(n29438), .B(n29439), .Z(n29369) );
  XNOR U29516 ( .A(n29440), .B(n29441), .Z(n29439) );
  XOR U29517 ( .A(n29391), .B(n29213), .Z(n29382) );
  XNOR U29518 ( .A(n29431), .B(n29179), .Z(n29213) );
  IV U29519 ( .A(n29380), .Z(n29431) );
  XOR U29520 ( .A(n29442), .B(n29443), .Z(n29380) );
  XOR U29521 ( .A(n29444), .B(n29445), .Z(n29443) );
  XNOR U29522 ( .A(n29093), .B(n29446), .Z(n29442) );
  ANDN U29523 ( .B(n29375), .A(n29391), .Z(n29437) );
  XNOR U29524 ( .A(n29093), .B(n29447), .Z(n29391) );
  XOR U29525 ( .A(n29146), .B(n29438), .Z(n29375) );
  XOR U29526 ( .A(n29448), .B(n29449), .Z(n29146) );
  XOR U29527 ( .A(n29450), .B(n29445), .Z(n29449) );
  XOR U29528 ( .A(msg[28]), .B(key[28]), .Z(n29445) );
  XNOR U29529 ( .A(n29447), .B(n29361), .Z(n29420) );
  XNOR U29530 ( .A(n29451), .B(n29424), .Z(n29432) );
  OR U29531 ( .A(n29360), .B(n29205), .Z(n29424) );
  XNOR U29532 ( .A(n29208), .B(n29179), .Z(n29205) );
  XOR U29533 ( .A(n29452), .B(n29448), .Z(n29179) );
  XNOR U29534 ( .A(n29438), .B(n29098), .Z(n29360) );
  XOR U29535 ( .A(n29448), .B(n29453), .Z(n29098) );
  XOR U29536 ( .A(n29440), .B(n29452), .Z(n29453) );
  IV U29537 ( .A(n29361), .Z(n29438) );
  ANDN U29538 ( .B(n29447), .A(n29361), .Z(n29451) );
  XNOR U29539 ( .A(n29448), .B(n29454), .Z(n29361) );
  XNOR U29540 ( .A(n29450), .B(n29444), .Z(n29454) );
  XNOR U29541 ( .A(msg[31]), .B(key[31]), .Z(n29444) );
  XNOR U29542 ( .A(msg[29]), .B(key[29]), .Z(n29448) );
  IV U29543 ( .A(n29208), .Z(n29447) );
  XNOR U29544 ( .A(n29441), .B(n29455), .Z(n29208) );
  XOR U29545 ( .A(n29446), .B(n29452), .Z(n29455) );
  IV U29546 ( .A(n29450), .Z(n29452) );
  XOR U29547 ( .A(n29093), .B(n29456), .Z(n29450) );
  XNOR U29548 ( .A(msg[30]), .B(key[30]), .Z(n29456) );
  XOR U29549 ( .A(msg[24]), .B(key[24]), .Z(n29093) );
  XNOR U29550 ( .A(n29440), .B(n29457), .Z(n29446) );
  XNOR U29551 ( .A(msg[27]), .B(key[27]), .Z(n29457) );
  XNOR U29552 ( .A(msg[25]), .B(key[25]), .Z(n29440) );
  XNOR U29553 ( .A(msg[26]), .B(key[26]), .Z(n29441) );
  XOR U29554 ( .A(n24474), .B(n29458), .Z(n29195) );
  XNOR U29555 ( .A(key[142]), .B(n25538), .Z(n29458) );
  XOR U29556 ( .A(n29083), .B(n29151), .Z(n25538) );
  XNOR U29557 ( .A(n29157), .B(n29459), .Z(n29151) );
  XNOR U29558 ( .A(n29460), .B(n29123), .Z(n29459) );
  NOR U29559 ( .A(n29218), .B(n29461), .Z(n29123) );
  XNOR U29560 ( .A(n29220), .B(n29166), .Z(n29218) );
  ANDN U29561 ( .B(n29220), .A(n29462), .Z(n29460) );
  XNOR U29562 ( .A(n29115), .B(n29463), .Z(n29157) );
  XNOR U29563 ( .A(n29464), .B(n29465), .Z(n29463) );
  OR U29564 ( .A(n29224), .B(n29466), .Z(n29465) );
  XOR U29565 ( .A(n29214), .B(n29152), .Z(n29083) );
  XOR U29566 ( .A(n29115), .B(n29467), .Z(n29152) );
  XNOR U29567 ( .A(n29154), .B(n29468), .Z(n29467) );
  NANDN U29568 ( .A(n29469), .B(n29470), .Z(n29468) );
  OR U29569 ( .A(n29471), .B(n29472), .Z(n29154) );
  XOR U29570 ( .A(n29473), .B(n29464), .Z(n29115) );
  NANDN U29571 ( .A(n29474), .B(n29475), .Z(n29464) );
  ANDN U29572 ( .B(n29476), .A(n29477), .Z(n29473) );
  XOR U29573 ( .A(n29479), .B(n29118), .Z(n29478) );
  OR U29574 ( .A(n29471), .B(n29480), .Z(n29118) );
  XOR U29575 ( .A(n29120), .B(n29481), .Z(n29471) );
  ANDN U29576 ( .B(n29482), .A(n29469), .Z(n29479) );
  XNOR U29577 ( .A(n29483), .B(n29222), .Z(n29161) );
  OR U29578 ( .A(n29474), .B(n29484), .Z(n29222) );
  XOR U29579 ( .A(n29485), .B(n29224), .Z(n29474) );
  XOR U29580 ( .A(n29481), .B(n29126), .Z(n29224) );
  IV U29581 ( .A(n29166), .Z(n29126) );
  XOR U29582 ( .A(n29486), .B(n29487), .Z(n29166) );
  NANDN U29583 ( .A(n29488), .B(n29489), .Z(n29487) );
  IV U29584 ( .A(n29469), .Z(n29481) );
  XNOR U29585 ( .A(n29490), .B(n29491), .Z(n29469) );
  NANDN U29586 ( .A(n29488), .B(n29492), .Z(n29491) );
  ANDN U29587 ( .B(n29485), .A(n29493), .Z(n29483) );
  IV U29588 ( .A(n29477), .Z(n29485) );
  XOR U29589 ( .A(n29220), .B(n29120), .Z(n29477) );
  XOR U29590 ( .A(n29494), .B(n29490), .Z(n29120) );
  NANDN U29591 ( .A(n29495), .B(n29496), .Z(n29490) );
  NANDN U29592 ( .A(n29495), .B(n29500), .Z(n29486) );
  XOR U29593 ( .A(n29501), .B(n29502), .Z(n29488) );
  XOR U29594 ( .A(n29503), .B(n29498), .Z(n29502) );
  XNOR U29595 ( .A(n29504), .B(n29505), .Z(n29501) );
  XNOR U29596 ( .A(n29506), .B(n29507), .Z(n29505) );
  ANDN U29597 ( .B(n29503), .A(n29498), .Z(n29506) );
  ANDN U29598 ( .B(n29503), .A(n29497), .Z(n29499) );
  XNOR U29599 ( .A(n29504), .B(n29508), .Z(n29497) );
  XOR U29600 ( .A(n29509), .B(n29507), .Z(n29508) );
  NAND U29601 ( .A(n29496), .B(n29500), .Z(n29507) );
  XNOR U29602 ( .A(n29492), .B(n29498), .Z(n29496) );
  XOR U29603 ( .A(n29510), .B(n29511), .Z(n29498) );
  XOR U29604 ( .A(n29512), .B(n29513), .Z(n29511) );
  XNOR U29605 ( .A(n29514), .B(n29515), .Z(n29510) );
  ANDN U29606 ( .B(n29219), .A(n29462), .Z(n29514) );
  AND U29607 ( .A(n29489), .B(n29492), .Z(n29509) );
  XNOR U29608 ( .A(n29489), .B(n29492), .Z(n29504) );
  XNOR U29609 ( .A(n29516), .B(n29517), .Z(n29492) );
  XNOR U29610 ( .A(n29518), .B(n29519), .Z(n29517) );
  XOR U29611 ( .A(n29512), .B(n29520), .Z(n29516) );
  XNOR U29612 ( .A(n29521), .B(n29515), .Z(n29520) );
  OR U29613 ( .A(n29461), .B(n29217), .Z(n29515) );
  XNOR U29614 ( .A(n29522), .B(n29165), .Z(n29217) );
  XNOR U29615 ( .A(n29462), .B(n29523), .Z(n29461) );
  NOR U29616 ( .A(n29523), .B(n29165), .Z(n29521) );
  XNOR U29617 ( .A(n29524), .B(n29525), .Z(n29489) );
  XNOR U29618 ( .A(n29526), .B(n29527), .Z(n29525) );
  XOR U29619 ( .A(n29156), .B(n29512), .Z(n29527) );
  XOR U29620 ( .A(n29219), .B(n29528), .Z(n29512) );
  XNOR U29621 ( .A(n29121), .B(n29529), .Z(n29524) );
  XNOR U29622 ( .A(n29530), .B(n29531), .Z(n29529) );
  ANDN U29623 ( .B(n29470), .A(n29532), .Z(n29530) );
  XNOR U29624 ( .A(n29533), .B(n29534), .Z(n29503) );
  XNOR U29625 ( .A(n29513), .B(n29535), .Z(n29534) );
  XNOR U29626 ( .A(n29470), .B(n29519), .Z(n29535) );
  XOR U29627 ( .A(n29165), .B(n29523), .Z(n29519) );
  XNOR U29628 ( .A(n29526), .B(n29536), .Z(n29513) );
  XNOR U29629 ( .A(n29537), .B(n29538), .Z(n29536) );
  NANDN U29630 ( .A(n29466), .B(n29225), .Z(n29538) );
  IV U29631 ( .A(n29518), .Z(n29526) );
  XNOR U29632 ( .A(n29539), .B(n29537), .Z(n29518) );
  NANDN U29633 ( .A(n29484), .B(n29475), .Z(n29537) );
  XOR U29634 ( .A(n29470), .B(n29523), .Z(n29466) );
  IV U29635 ( .A(n29125), .Z(n29523) );
  XOR U29636 ( .A(n29540), .B(n29541), .Z(n29125) );
  XNOR U29637 ( .A(n29542), .B(n29543), .Z(n29541) );
  XOR U29638 ( .A(n29493), .B(n29225), .Z(n29484) );
  XNOR U29639 ( .A(n29482), .B(n29165), .Z(n29225) );
  XNOR U29640 ( .A(n29543), .B(n29540), .Z(n29165) );
  ANDN U29641 ( .B(n29476), .A(n29493), .Z(n29539) );
  XNOR U29642 ( .A(n29544), .B(n29219), .Z(n29493) );
  IV U29643 ( .A(n29522), .Z(n29219) );
  XNOR U29644 ( .A(n29545), .B(n29546), .Z(n29522) );
  XNOR U29645 ( .A(n29547), .B(n29543), .Z(n29546) );
  XOR U29646 ( .A(n29548), .B(n29528), .Z(n29476) );
  XNOR U29647 ( .A(n29532), .B(n29549), .Z(n29533) );
  XNOR U29648 ( .A(n29550), .B(n29531), .Z(n29549) );
  OR U29649 ( .A(n29472), .B(n29480), .Z(n29531) );
  XOR U29650 ( .A(n29121), .B(n29482), .Z(n29480) );
  IV U29651 ( .A(n29532), .Z(n29482) );
  XOR U29652 ( .A(n29156), .B(n29470), .Z(n29472) );
  XNOR U29653 ( .A(n29528), .B(n29551), .Z(n29470) );
  XNOR U29654 ( .A(n29542), .B(n29545), .Z(n29551) );
  XNOR U29655 ( .A(msg[114]), .B(key[114]), .Z(n29545) );
  IV U29656 ( .A(n29462), .Z(n29528) );
  XOR U29657 ( .A(n29552), .B(n29553), .Z(n29462) );
  XOR U29658 ( .A(n29543), .B(n29554), .Z(n29553) );
  IV U29659 ( .A(n29548), .Z(n29156) );
  ANDN U29660 ( .B(n29548), .A(n29121), .Z(n29550) );
  XOR U29661 ( .A(n29540), .B(n29555), .Z(n29548) );
  XNOR U29662 ( .A(n29543), .B(n29556), .Z(n29555) );
  XOR U29663 ( .A(n29544), .B(n29557), .Z(n29543) );
  XNOR U29664 ( .A(msg[118]), .B(key[118]), .Z(n29557) );
  IV U29665 ( .A(n29552), .Z(n29540) );
  XOR U29666 ( .A(msg[117]), .B(key[117]), .Z(n29552) );
  XOR U29667 ( .A(n29558), .B(n29559), .Z(n29532) );
  XOR U29668 ( .A(n29556), .B(n29554), .Z(n29559) );
  XOR U29669 ( .A(msg[119]), .B(key[119]), .Z(n29554) );
  XNOR U29670 ( .A(msg[116]), .B(key[116]), .Z(n29556) );
  XOR U29671 ( .A(n29121), .B(n29547), .Z(n29558) );
  XNOR U29672 ( .A(n29542), .B(n29560), .Z(n29547) );
  XNOR U29673 ( .A(msg[115]), .B(key[115]), .Z(n29560) );
  XNOR U29674 ( .A(msg[113]), .B(key[113]), .Z(n29542) );
  IV U29675 ( .A(n29544), .Z(n29121) );
  XOR U29676 ( .A(msg[112]), .B(key[112]), .Z(n29544) );
  XNOR U29677 ( .A(n24488), .B(n25529), .Z(n24474) );
  XNOR U29678 ( .A(n29561), .B(n29562), .Z(n25529) );
  XOR U29679 ( .A(n29201), .B(n29103), .Z(n29562) );
  XNOR U29680 ( .A(n29563), .B(n29564), .Z(n29103) );
  XNOR U29681 ( .A(n29565), .B(n29566), .Z(n29564) );
  NANDN U29682 ( .A(n29567), .B(n29568), .Z(n29566) );
  XOR U29683 ( .A(n29182), .B(n29169), .Z(n29201) );
  XNOR U29684 ( .A(n29104), .B(n29569), .Z(n29169) );
  XNOR U29685 ( .A(n29570), .B(n29571), .Z(n29569) );
  OR U29686 ( .A(n29572), .B(n29573), .Z(n29571) );
  XOR U29687 ( .A(n29181), .B(n29172), .Z(n29561) );
  XNOR U29688 ( .A(n29570), .B(n29575), .Z(n29574) );
  NANDN U29689 ( .A(n29567), .B(n29576), .Z(n29575) );
  OR U29690 ( .A(n29577), .B(n29578), .Z(n29570) );
  XOR U29691 ( .A(n29104), .B(n29579), .Z(n29351) );
  XNOR U29692 ( .A(n29580), .B(n29581), .Z(n29579) );
  NAND U29693 ( .A(n29582), .B(n29583), .Z(n29581) );
  XNOR U29694 ( .A(n29584), .B(n29580), .Z(n29104) );
  NANDN U29695 ( .A(n29585), .B(n29586), .Z(n29580) );
  ANDN U29696 ( .B(n29587), .A(n29588), .Z(n29584) );
  IV U29697 ( .A(n29171), .Z(n29181) );
  XOR U29698 ( .A(n29589), .B(n29590), .Z(n29171) );
  XNOR U29699 ( .A(n29591), .B(n29592), .Z(n29590) );
  NANDN U29700 ( .A(n29593), .B(n29594), .Z(n29592) );
  XOR U29701 ( .A(n29563), .B(n29595), .Z(n29102) );
  XOR U29702 ( .A(n29596), .B(n29591), .Z(n29595) );
  OR U29703 ( .A(n29597), .B(n29354), .Z(n29591) );
  XNOR U29704 ( .A(n29356), .B(n29594), .Z(n29354) );
  ANDN U29705 ( .B(n29356), .A(n29598), .Z(n29596) );
  XOR U29706 ( .A(n29589), .B(n29599), .Z(n29563) );
  XNOR U29707 ( .A(n29600), .B(n29601), .Z(n29599) );
  NAND U29708 ( .A(n29582), .B(n29602), .Z(n29601) );
  XOR U29709 ( .A(n29604), .B(n29565), .Z(n29603) );
  OR U29710 ( .A(n29605), .B(n29577), .Z(n29565) );
  XNOR U29711 ( .A(n29567), .B(n29572), .Z(n29577) );
  NOR U29712 ( .A(n29606), .B(n29572), .Z(n29604) );
  XNOR U29713 ( .A(n29607), .B(n29600), .Z(n29589) );
  OR U29714 ( .A(n29585), .B(n29608), .Z(n29600) );
  XNOR U29715 ( .A(n29609), .B(n29582), .Z(n29585) );
  XNOR U29716 ( .A(n29572), .B(n29594), .Z(n29582) );
  IV U29717 ( .A(n29109), .Z(n29594) );
  XNOR U29718 ( .A(n29610), .B(n29611), .Z(n29109) );
  NANDN U29719 ( .A(n29612), .B(n29613), .Z(n29611) );
  XNOR U29720 ( .A(n29614), .B(n29615), .Z(n29572) );
  NANDN U29721 ( .A(n29612), .B(n29616), .Z(n29615) );
  ANDN U29722 ( .B(n29609), .A(n29617), .Z(n29607) );
  IV U29723 ( .A(n29588), .Z(n29609) );
  XOR U29724 ( .A(n29567), .B(n29356), .Z(n29588) );
  XNOR U29725 ( .A(n29618), .B(n29610), .Z(n29356) );
  NANDN U29726 ( .A(n29619), .B(n29620), .Z(n29610) );
  XOR U29727 ( .A(n29613), .B(n29621), .Z(n29620) );
  ANDN U29728 ( .B(n29621), .A(n29622), .Z(n29618) );
  NANDN U29729 ( .A(n29619), .B(n29624), .Z(n29614) );
  XOR U29730 ( .A(n29625), .B(n29626), .Z(n29612) );
  XOR U29731 ( .A(n29627), .B(n29628), .Z(n29626) );
  XNOR U29732 ( .A(n29629), .B(n29630), .Z(n29625) );
  XNOR U29733 ( .A(n29631), .B(n29632), .Z(n29630) );
  ANDN U29734 ( .B(n29628), .A(n29627), .Z(n29631) );
  ANDN U29735 ( .B(n29628), .A(n29622), .Z(n29623) );
  XNOR U29736 ( .A(n29629), .B(n29633), .Z(n29622) );
  XOR U29737 ( .A(n29634), .B(n29632), .Z(n29633) );
  NAND U29738 ( .A(n29624), .B(n29635), .Z(n29632) );
  XNOR U29739 ( .A(n29613), .B(n29627), .Z(n29635) );
  IV U29740 ( .A(n29621), .Z(n29627) );
  XNOR U29741 ( .A(n29636), .B(n29637), .Z(n29621) );
  XNOR U29742 ( .A(n29638), .B(n29639), .Z(n29637) );
  XOR U29743 ( .A(n29573), .B(n29640), .Z(n29639) );
  XNOR U29744 ( .A(n29606), .B(n29641), .Z(n29636) );
  XNOR U29745 ( .A(n29642), .B(n29643), .Z(n29641) );
  AND U29746 ( .A(n29576), .B(n29568), .Z(n29642) );
  XOR U29747 ( .A(n29616), .B(n29628), .Z(n29624) );
  AND U29748 ( .A(n29613), .B(n29616), .Z(n29634) );
  XNOR U29749 ( .A(n29613), .B(n29616), .Z(n29629) );
  XNOR U29750 ( .A(n29644), .B(n29645), .Z(n29616) );
  XNOR U29751 ( .A(n29646), .B(n29640), .Z(n29645) );
  XOR U29752 ( .A(n29647), .B(n29648), .Z(n29644) );
  XNOR U29753 ( .A(n29649), .B(n29650), .Z(n29648) );
  ANDN U29754 ( .B(n29108), .A(n29593), .Z(n29649) );
  XNOR U29755 ( .A(n29651), .B(n29652), .Z(n29613) );
  XNOR U29756 ( .A(n29576), .B(n29647), .Z(n29653) );
  XOR U29757 ( .A(n29568), .B(n29654), .Z(n29651) );
  XNOR U29758 ( .A(n29655), .B(n29643), .Z(n29654) );
  OR U29759 ( .A(n29578), .B(n29605), .Z(n29643) );
  XOR U29760 ( .A(n29568), .B(n29606), .Z(n29605) );
  XNOR U29761 ( .A(n29576), .B(n29656), .Z(n29578) );
  ANDN U29762 ( .B(n29657), .A(n29573), .Z(n29655) );
  XNOR U29763 ( .A(n29658), .B(n29659), .Z(n29628) );
  XOR U29764 ( .A(n29646), .B(n29638), .Z(n29659) );
  XOR U29765 ( .A(n29647), .B(n29660), .Z(n29638) );
  XNOR U29766 ( .A(n29661), .B(n29662), .Z(n29660) );
  NAND U29767 ( .A(n29602), .B(n29583), .Z(n29662) );
  XNOR U29768 ( .A(n29663), .B(n29661), .Z(n29647) );
  NANDN U29769 ( .A(n29608), .B(n29586), .Z(n29661) );
  XOR U29770 ( .A(n29587), .B(n29583), .Z(n29586) );
  XOR U29771 ( .A(n29656), .B(n29108), .Z(n29583) );
  IV U29772 ( .A(n29573), .Z(n29656) );
  XOR U29773 ( .A(n29664), .B(n29665), .Z(n29573) );
  XNOR U29774 ( .A(n29666), .B(n29667), .Z(n29665) );
  XOR U29775 ( .A(n29617), .B(n29602), .Z(n29608) );
  XNOR U29776 ( .A(n29657), .B(n29593), .Z(n29602) );
  IV U29777 ( .A(n29606), .Z(n29657) );
  XOR U29778 ( .A(n29668), .B(n29669), .Z(n29606) );
  XOR U29779 ( .A(n29670), .B(n29671), .Z(n29669) );
  XNOR U29780 ( .A(n29568), .B(n29672), .Z(n29668) );
  ANDN U29781 ( .B(n29587), .A(n29617), .Z(n29663) );
  XNOR U29782 ( .A(n29568), .B(n29673), .Z(n29617) );
  XOR U29783 ( .A(n29576), .B(n29664), .Z(n29587) );
  XOR U29784 ( .A(n29674), .B(n29675), .Z(n29576) );
  XOR U29785 ( .A(n29676), .B(n29671), .Z(n29675) );
  XOR U29786 ( .A(msg[36]), .B(key[36]), .Z(n29671) );
  XNOR U29787 ( .A(n29673), .B(n29357), .Z(n29646) );
  XNOR U29788 ( .A(n29677), .B(n29650), .Z(n29658) );
  OR U29789 ( .A(n29355), .B(n29597), .Z(n29650) );
  XNOR U29790 ( .A(n29598), .B(n29593), .Z(n29597) );
  XOR U29791 ( .A(n29678), .B(n29674), .Z(n29593) );
  XNOR U29792 ( .A(n29664), .B(n29108), .Z(n29355) );
  XOR U29793 ( .A(n29674), .B(n29679), .Z(n29108) );
  XOR U29794 ( .A(n29666), .B(n29678), .Z(n29679) );
  IV U29795 ( .A(n29357), .Z(n29664) );
  ANDN U29796 ( .B(n29673), .A(n29357), .Z(n29677) );
  XNOR U29797 ( .A(n29674), .B(n29680), .Z(n29357) );
  XNOR U29798 ( .A(n29676), .B(n29670), .Z(n29680) );
  XNOR U29799 ( .A(msg[39]), .B(key[39]), .Z(n29670) );
  XNOR U29800 ( .A(msg[37]), .B(key[37]), .Z(n29674) );
  IV U29801 ( .A(n29598), .Z(n29673) );
  XNOR U29802 ( .A(n29667), .B(n29681), .Z(n29598) );
  XOR U29803 ( .A(n29672), .B(n29678), .Z(n29681) );
  IV U29804 ( .A(n29676), .Z(n29678) );
  XOR U29805 ( .A(n29568), .B(n29682), .Z(n29676) );
  XNOR U29806 ( .A(msg[38]), .B(key[38]), .Z(n29682) );
  XOR U29807 ( .A(msg[32]), .B(key[32]), .Z(n29568) );
  XNOR U29808 ( .A(n29666), .B(n29683), .Z(n29672) );
  XNOR U29809 ( .A(msg[35]), .B(key[35]), .Z(n29683) );
  XNOR U29810 ( .A(msg[33]), .B(key[33]), .Z(n29666) );
  XNOR U29811 ( .A(msg[34]), .B(key[34]), .Z(n29667) );
endmodule

