
module matrixMult_N_M_1_N16_M32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_3 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_8 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_4 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_10 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_5 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_12 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_6 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_14 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_7 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_16 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_8 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_18 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_9 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_20 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_10 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_22 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_11 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_24 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_12 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_26 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_13 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_28 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_14 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32_DW01_add_30 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[31]) );
  XNOR U16 ( .A(B[31]), .B(A[31]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n15) );
  NAND U18 ( .A(n19), .B(B[30]), .Z(n18) );
  NANDN U19 ( .A(A[30]), .B(n20), .Z(n19) );
  NANDN U20 ( .A(n20), .B(A[30]), .Z(n17) );
  XOR U21 ( .A(n20), .B(n21), .Z(SUM[30]) );
  XNOR U22 ( .A(B[30]), .B(A[30]), .Z(n21) );
  AND U23 ( .A(n22), .B(n23), .Z(n20) );
  NAND U24 ( .A(n24), .B(B[29]), .Z(n23) );
  NANDN U25 ( .A(A[29]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(n25), .B(A[29]), .Z(n22) );
  XOR U27 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n27) );
  XOR U29 ( .A(n25), .B(n28), .Z(SUM[29]) );
  XNOR U30 ( .A(B[29]), .B(A[29]), .Z(n28) );
  AND U31 ( .A(n29), .B(n30), .Z(n25) );
  NAND U32 ( .A(n31), .B(B[28]), .Z(n30) );
  NANDN U33 ( .A(A[28]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(n32), .B(A[28]), .Z(n29) );
  XOR U35 ( .A(n32), .B(n33), .Z(SUM[28]) );
  XNOR U36 ( .A(B[28]), .B(A[28]), .Z(n33) );
  AND U37 ( .A(n34), .B(n35), .Z(n32) );
  NAND U38 ( .A(n36), .B(B[27]), .Z(n35) );
  NANDN U39 ( .A(A[27]), .B(n37), .Z(n36) );
  NANDN U40 ( .A(n37), .B(A[27]), .Z(n34) );
  XOR U41 ( .A(n37), .B(n38), .Z(SUM[27]) );
  XNOR U42 ( .A(B[27]), .B(A[27]), .Z(n38) );
  AND U43 ( .A(n39), .B(n40), .Z(n37) );
  NAND U44 ( .A(n41), .B(B[26]), .Z(n40) );
  NANDN U45 ( .A(A[26]), .B(n42), .Z(n41) );
  NANDN U46 ( .A(n42), .B(A[26]), .Z(n39) );
  XOR U47 ( .A(n42), .B(n43), .Z(SUM[26]) );
  XNOR U48 ( .A(B[26]), .B(A[26]), .Z(n43) );
  AND U49 ( .A(n44), .B(n45), .Z(n42) );
  NAND U50 ( .A(n46), .B(B[25]), .Z(n45) );
  NANDN U51 ( .A(A[25]), .B(n47), .Z(n46) );
  NANDN U52 ( .A(n47), .B(A[25]), .Z(n44) );
  XOR U53 ( .A(n47), .B(n48), .Z(SUM[25]) );
  XNOR U54 ( .A(B[25]), .B(A[25]), .Z(n48) );
  AND U55 ( .A(n49), .B(n50), .Z(n47) );
  NAND U56 ( .A(n51), .B(B[24]), .Z(n50) );
  NANDN U57 ( .A(A[24]), .B(n52), .Z(n51) );
  NANDN U58 ( .A(n52), .B(A[24]), .Z(n49) );
  XOR U59 ( .A(n52), .B(n53), .Z(SUM[24]) );
  XNOR U60 ( .A(B[24]), .B(A[24]), .Z(n53) );
  AND U61 ( .A(n54), .B(n55), .Z(n52) );
  NAND U62 ( .A(n56), .B(B[23]), .Z(n55) );
  NANDN U63 ( .A(A[23]), .B(n57), .Z(n56) );
  NANDN U64 ( .A(n57), .B(A[23]), .Z(n54) );
  XOR U65 ( .A(n57), .B(n58), .Z(SUM[23]) );
  XNOR U66 ( .A(B[23]), .B(A[23]), .Z(n58) );
  AND U67 ( .A(n59), .B(n60), .Z(n57) );
  NAND U68 ( .A(n61), .B(B[22]), .Z(n60) );
  NANDN U69 ( .A(A[22]), .B(n62), .Z(n61) );
  NANDN U70 ( .A(n62), .B(A[22]), .Z(n59) );
  XOR U71 ( .A(n62), .B(n63), .Z(SUM[22]) );
  XNOR U72 ( .A(B[22]), .B(A[22]), .Z(n63) );
  AND U73 ( .A(n64), .B(n65), .Z(n62) );
  NAND U74 ( .A(n66), .B(B[21]), .Z(n65) );
  NANDN U75 ( .A(A[21]), .B(n67), .Z(n66) );
  NANDN U76 ( .A(n67), .B(A[21]), .Z(n64) );
  XOR U77 ( .A(n67), .B(n68), .Z(SUM[21]) );
  XNOR U78 ( .A(B[21]), .B(A[21]), .Z(n68) );
  AND U79 ( .A(n69), .B(n70), .Z(n67) );
  NAND U80 ( .A(n71), .B(B[20]), .Z(n70) );
  NANDN U81 ( .A(A[20]), .B(n72), .Z(n71) );
  NANDN U82 ( .A(n72), .B(A[20]), .Z(n69) );
  XOR U83 ( .A(n72), .B(n73), .Z(SUM[20]) );
  XNOR U84 ( .A(B[20]), .B(A[20]), .Z(n73) );
  AND U85 ( .A(n74), .B(n75), .Z(n72) );
  NAND U86 ( .A(n76), .B(B[19]), .Z(n75) );
  NANDN U87 ( .A(A[19]), .B(n77), .Z(n76) );
  NANDN U88 ( .A(n77), .B(A[19]), .Z(n74) );
  XOR U89 ( .A(n78), .B(n79), .Z(SUM[1]) );
  XOR U90 ( .A(B[1]), .B(A[1]), .Z(n79) );
  XOR U91 ( .A(n77), .B(n80), .Z(SUM[19]) );
  XNOR U92 ( .A(B[19]), .B(A[19]), .Z(n80) );
  AND U93 ( .A(n81), .B(n82), .Z(n77) );
  NAND U94 ( .A(n83), .B(B[18]), .Z(n82) );
  NANDN U95 ( .A(A[18]), .B(n84), .Z(n83) );
  NANDN U96 ( .A(n84), .B(A[18]), .Z(n81) );
  XOR U97 ( .A(n84), .B(n85), .Z(SUM[18]) );
  XNOR U98 ( .A(B[18]), .B(A[18]), .Z(n85) );
  AND U99 ( .A(n86), .B(n87), .Z(n84) );
  NAND U100 ( .A(n88), .B(B[17]), .Z(n87) );
  NANDN U101 ( .A(A[17]), .B(n89), .Z(n88) );
  NANDN U102 ( .A(n89), .B(A[17]), .Z(n86) );
  XOR U103 ( .A(n89), .B(n90), .Z(SUM[17]) );
  XNOR U104 ( .A(B[17]), .B(A[17]), .Z(n90) );
  AND U105 ( .A(n91), .B(n92), .Z(n89) );
  NAND U106 ( .A(n93), .B(B[16]), .Z(n92) );
  NANDN U107 ( .A(A[16]), .B(n94), .Z(n93) );
  NANDN U108 ( .A(n94), .B(A[16]), .Z(n91) );
  XOR U109 ( .A(n94), .B(n95), .Z(SUM[16]) );
  XNOR U110 ( .A(B[16]), .B(A[16]), .Z(n95) );
  AND U111 ( .A(n96), .B(n97), .Z(n94) );
  NAND U112 ( .A(n98), .B(B[15]), .Z(n97) );
  NANDN U113 ( .A(A[15]), .B(n99), .Z(n98) );
  NANDN U114 ( .A(n99), .B(A[15]), .Z(n96) );
  XOR U115 ( .A(n99), .B(n100), .Z(SUM[15]) );
  XNOR U116 ( .A(B[15]), .B(A[15]), .Z(n100) );
  AND U117 ( .A(n101), .B(n102), .Z(n99) );
  NAND U118 ( .A(n103), .B(B[14]), .Z(n102) );
  NANDN U119 ( .A(A[14]), .B(n104), .Z(n103) );
  NANDN U120 ( .A(n104), .B(A[14]), .Z(n101) );
  XOR U121 ( .A(n104), .B(n105), .Z(SUM[14]) );
  XNOR U122 ( .A(B[14]), .B(A[14]), .Z(n105) );
  AND U123 ( .A(n106), .B(n107), .Z(n104) );
  NAND U124 ( .A(n108), .B(B[13]), .Z(n107) );
  NANDN U125 ( .A(A[13]), .B(n109), .Z(n108) );
  NANDN U126 ( .A(n109), .B(A[13]), .Z(n106) );
  XOR U127 ( .A(n109), .B(n110), .Z(SUM[13]) );
  XNOR U128 ( .A(B[13]), .B(A[13]), .Z(n110) );
  AND U129 ( .A(n111), .B(n112), .Z(n109) );
  NAND U130 ( .A(n113), .B(B[12]), .Z(n112) );
  NANDN U131 ( .A(A[12]), .B(n114), .Z(n113) );
  NANDN U132 ( .A(n114), .B(A[12]), .Z(n111) );
  XOR U133 ( .A(n114), .B(n115), .Z(SUM[12]) );
  XNOR U134 ( .A(B[12]), .B(A[12]), .Z(n115) );
  AND U135 ( .A(n116), .B(n117), .Z(n114) );
  NAND U136 ( .A(n118), .B(B[11]), .Z(n117) );
  NANDN U137 ( .A(A[11]), .B(n119), .Z(n118) );
  NANDN U138 ( .A(n119), .B(A[11]), .Z(n116) );
  XOR U139 ( .A(n119), .B(n120), .Z(SUM[11]) );
  XNOR U140 ( .A(B[11]), .B(A[11]), .Z(n120) );
  AND U141 ( .A(n121), .B(n122), .Z(n119) );
  NAND U142 ( .A(n123), .B(B[10]), .Z(n122) );
  NANDN U143 ( .A(A[10]), .B(n124), .Z(n123) );
  NANDN U144 ( .A(n124), .B(A[10]), .Z(n121) );
  XOR U145 ( .A(n124), .B(n125), .Z(SUM[10]) );
  XNOR U146 ( .A(B[10]), .B(A[10]), .Z(n125) );
  AND U147 ( .A(n126), .B(n127), .Z(n124) );
  NAND U148 ( .A(n128), .B(B[9]), .Z(n127) );
  NANDN U149 ( .A(A[9]), .B(n1), .Z(n128) );
  NANDN U150 ( .A(n1), .B(A[9]), .Z(n126) );
  AND U151 ( .A(n129), .B(n130), .Z(n1) );
  NAND U152 ( .A(n131), .B(B[8]), .Z(n130) );
  NANDN U153 ( .A(A[8]), .B(n3), .Z(n131) );
  NANDN U154 ( .A(n3), .B(A[8]), .Z(n129) );
  AND U155 ( .A(n132), .B(n133), .Z(n3) );
  NAND U156 ( .A(n134), .B(B[7]), .Z(n133) );
  NANDN U157 ( .A(A[7]), .B(n5), .Z(n134) );
  NANDN U158 ( .A(n5), .B(A[7]), .Z(n132) );
  AND U159 ( .A(n135), .B(n136), .Z(n5) );
  NAND U160 ( .A(n137), .B(B[6]), .Z(n136) );
  NANDN U161 ( .A(A[6]), .B(n7), .Z(n137) );
  NANDN U162 ( .A(n7), .B(A[6]), .Z(n135) );
  AND U163 ( .A(n138), .B(n139), .Z(n7) );
  NAND U164 ( .A(n140), .B(B[5]), .Z(n139) );
  NANDN U165 ( .A(A[5]), .B(n9), .Z(n140) );
  NANDN U166 ( .A(n9), .B(A[5]), .Z(n138) );
  AND U167 ( .A(n141), .B(n142), .Z(n9) );
  NAND U168 ( .A(n143), .B(B[4]), .Z(n142) );
  NANDN U169 ( .A(A[4]), .B(n11), .Z(n143) );
  NANDN U170 ( .A(n11), .B(A[4]), .Z(n141) );
  AND U171 ( .A(n144), .B(n145), .Z(n11) );
  NAND U172 ( .A(n146), .B(B[3]), .Z(n145) );
  NANDN U173 ( .A(A[3]), .B(n13), .Z(n146) );
  NANDN U174 ( .A(n13), .B(A[3]), .Z(n144) );
  AND U175 ( .A(n147), .B(n148), .Z(n13) );
  NAND U176 ( .A(n149), .B(B[2]), .Z(n148) );
  NANDN U177 ( .A(A[2]), .B(n26), .Z(n149) );
  NANDN U178 ( .A(n26), .B(A[2]), .Z(n147) );
  AND U179 ( .A(n150), .B(n151), .Z(n26) );
  NAND U180 ( .A(n152), .B(B[1]), .Z(n151) );
  OR U181 ( .A(n78), .B(A[1]), .Z(n152) );
  NAND U182 ( .A(n78), .B(A[1]), .Z(n150) );
  AND U183 ( .A(B[0]), .B(A[0]), .Z(n78) );
  XOR U184 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module matrixMult_N_M_1_N16_M32_DW02_mult_15 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298;

  IV U2 ( .A(A[31]), .Z(n3) );
  IV U3 ( .A(n2908), .Z(n4) );
  IV U4 ( .A(n2909), .Z(n5) );
  IV U5 ( .A(n2923), .Z(n6) );
  IV U6 ( .A(n2924), .Z(n7) );
  IV U7 ( .A(n2938), .Z(n8) );
  IV U8 ( .A(n2939), .Z(n9) );
  IV U9 ( .A(n2953), .Z(n10) );
  IV U10 ( .A(n2954), .Z(n11) );
  IV U11 ( .A(n365), .Z(n12) );
  IV U12 ( .A(n565), .Z(n13) );
  IV U13 ( .A(n758), .Z(n14) );
  IV U14 ( .A(n944), .Z(n15) );
  IV U15 ( .A(n1123), .Z(n16) );
  IV U16 ( .A(n1295), .Z(n17) );
  IV U17 ( .A(n1460), .Z(n18) );
  IV U18 ( .A(n1618), .Z(n19) );
  IV U19 ( .A(n1769), .Z(n20) );
  IV U20 ( .A(n1913), .Z(n21) );
  IV U21 ( .A(n2054), .Z(n22) );
  IV U22 ( .A(n2184), .Z(n23) );
  IV U23 ( .A(n2307), .Z(n24) );
  IV U24 ( .A(n2423), .Z(n25) );
  IV U25 ( .A(n2532), .Z(n26) );
  IV U26 ( .A(n2634), .Z(n27) );
  IV U27 ( .A(n2729), .Z(n28) );
  IV U28 ( .A(n2817), .Z(n29) );
  IV U29 ( .A(n2974), .Z(n30) );
  IV U30 ( .A(n3010), .Z(n31) );
  IV U31 ( .A(n3070), .Z(n32) );
  IV U32 ( .A(n3123), .Z(n33) );
  IV U33 ( .A(n3169), .Z(n34) );
  IV U34 ( .A(n3208), .Z(n35) );
  IV U35 ( .A(n3240), .Z(n36) );
  IV U36 ( .A(n3265), .Z(n37) );
  IV U37 ( .A(n3283), .Z(n38) );
  IV U38 ( .A(n2898), .Z(n39) );
  IV U39 ( .A(n2973), .Z(n40) );
  IV U40 ( .A(B[1]), .Z(n41) );
  IV U41 ( .A(B[0]), .Z(n42) );
  XNOR U42 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U43 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  XOR U44 ( .A(n45), .B(n46), .Z(PRODUCT[11]) );
  XNOR U45 ( .A(n47), .B(n4), .Z(n46) );
  XNOR U46 ( .A(n48), .B(n49), .Z(PRODUCT[10]) );
  XNOR U47 ( .A(n50), .B(n51), .Z(n49) );
  XOR U48 ( .A(n52), .B(n53), .Z(PRODUCT[9]) );
  XNOR U49 ( .A(n54), .B(n6), .Z(n53) );
  XNOR U50 ( .A(n55), .B(n56), .Z(PRODUCT[8]) );
  XNOR U51 ( .A(n57), .B(n58), .Z(n56) );
  XOR U52 ( .A(n59), .B(n60), .Z(PRODUCT[7]) );
  XNOR U53 ( .A(n61), .B(n8), .Z(n60) );
  XNOR U54 ( .A(n62), .B(n63), .Z(PRODUCT[6]) );
  XNOR U55 ( .A(n64), .B(n65), .Z(n63) );
  XOR U56 ( .A(n66), .B(n67), .Z(PRODUCT[5]) );
  XNOR U57 ( .A(n68), .B(n10), .Z(n67) );
  XNOR U58 ( .A(n160), .B(n161), .Z(PRODUCT[4]) );
  XNOR U59 ( .A(n162), .B(n163), .Z(n161) );
  XOR U60 ( .A(n159), .B(n164), .Z(PRODUCT[31]) );
  XNOR U61 ( .A(n158), .B(n157), .Z(n164) );
  AND U62 ( .A(n165), .B(n166), .Z(n157) );
  NAND U63 ( .A(n167), .B(n168), .Z(n166) );
  NANDN U64 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U65 ( .A(n170), .B(n169), .Z(n165) );
  ANDN U66 ( .B(B[0]), .A(n3), .Z(n158) );
  XNOR U67 ( .A(n71), .B(n171), .Z(n159) );
  XNOR U68 ( .A(n70), .B(n69), .Z(n171) );
  AND U69 ( .A(n172), .B(n173), .Z(n69) );
  NANDN U70 ( .A(n174), .B(n175), .Z(n173) );
  OR U71 ( .A(n176), .B(n177), .Z(n175) );
  NAND U72 ( .A(n177), .B(n176), .Z(n172) );
  ANDN U73 ( .B(A[30]), .A(n41), .Z(n70) );
  XNOR U74 ( .A(n74), .B(n178), .Z(n71) );
  XNOR U75 ( .A(n73), .B(n72), .Z(n178) );
  AND U76 ( .A(n179), .B(n180), .Z(n72) );
  NANDN U77 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U78 ( .A(n183), .B(n184), .Z(n182) );
  NANDN U79 ( .A(n184), .B(n183), .Z(n179) );
  AND U80 ( .A(A[29]), .B(B[2]), .Z(n73) );
  XNOR U81 ( .A(n77), .B(n185), .Z(n74) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n185) );
  AND U83 ( .A(n186), .B(n187), .Z(n75) );
  NANDN U84 ( .A(n188), .B(n189), .Z(n187) );
  OR U85 ( .A(n190), .B(n191), .Z(n189) );
  NAND U86 ( .A(n191), .B(n190), .Z(n186) );
  AND U87 ( .A(A[28]), .B(B[3]), .Z(n76) );
  XNOR U88 ( .A(n80), .B(n192), .Z(n77) );
  XNOR U89 ( .A(n79), .B(n78), .Z(n192) );
  AND U90 ( .A(n193), .B(n194), .Z(n78) );
  NANDN U91 ( .A(n195), .B(n196), .Z(n194) );
  NANDN U92 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U93 ( .A(n198), .B(n197), .Z(n193) );
  AND U94 ( .A(A[27]), .B(B[4]), .Z(n79) );
  XNOR U95 ( .A(n83), .B(n199), .Z(n80) );
  XNOR U96 ( .A(n82), .B(n81), .Z(n199) );
  AND U97 ( .A(n200), .B(n201), .Z(n81) );
  NANDN U98 ( .A(n202), .B(n203), .Z(n201) );
  OR U99 ( .A(n204), .B(n205), .Z(n203) );
  NAND U100 ( .A(n205), .B(n204), .Z(n200) );
  AND U101 ( .A(A[26]), .B(B[5]), .Z(n82) );
  XNOR U102 ( .A(n86), .B(n206), .Z(n83) );
  XNOR U103 ( .A(n85), .B(n84), .Z(n206) );
  AND U104 ( .A(n207), .B(n208), .Z(n84) );
  NANDN U105 ( .A(n209), .B(n210), .Z(n208) );
  NANDN U106 ( .A(n211), .B(n212), .Z(n210) );
  NANDN U107 ( .A(n212), .B(n211), .Z(n207) );
  AND U108 ( .A(A[25]), .B(B[6]), .Z(n85) );
  XNOR U109 ( .A(n89), .B(n213), .Z(n86) );
  XNOR U110 ( .A(n88), .B(n87), .Z(n213) );
  AND U111 ( .A(n214), .B(n215), .Z(n87) );
  NANDN U112 ( .A(n216), .B(n217), .Z(n215) );
  OR U113 ( .A(n218), .B(n219), .Z(n217) );
  NAND U114 ( .A(n219), .B(n218), .Z(n214) );
  AND U115 ( .A(A[24]), .B(B[7]), .Z(n88) );
  XNOR U116 ( .A(n92), .B(n220), .Z(n89) );
  XNOR U117 ( .A(n91), .B(n90), .Z(n220) );
  AND U118 ( .A(n221), .B(n222), .Z(n90) );
  NANDN U119 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U120 ( .A(n225), .B(n226), .Z(n224) );
  NANDN U121 ( .A(n226), .B(n225), .Z(n221) );
  AND U122 ( .A(A[23]), .B(B[8]), .Z(n91) );
  XNOR U123 ( .A(n95), .B(n227), .Z(n92) );
  XNOR U124 ( .A(n94), .B(n93), .Z(n227) );
  AND U125 ( .A(n228), .B(n229), .Z(n93) );
  NANDN U126 ( .A(n230), .B(n231), .Z(n229) );
  OR U127 ( .A(n232), .B(n233), .Z(n231) );
  NAND U128 ( .A(n233), .B(n232), .Z(n228) );
  AND U129 ( .A(A[22]), .B(B[9]), .Z(n94) );
  XNOR U130 ( .A(n98), .B(n234), .Z(n95) );
  XNOR U131 ( .A(n97), .B(n96), .Z(n234) );
  AND U132 ( .A(n235), .B(n236), .Z(n96) );
  NANDN U133 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U134 ( .A(n239), .B(n240), .Z(n238) );
  NANDN U135 ( .A(n240), .B(n239), .Z(n235) );
  AND U136 ( .A(A[21]), .B(B[10]), .Z(n97) );
  XNOR U137 ( .A(n101), .B(n241), .Z(n98) );
  XNOR U138 ( .A(n100), .B(n99), .Z(n241) );
  AND U139 ( .A(n242), .B(n243), .Z(n99) );
  NANDN U140 ( .A(n244), .B(n245), .Z(n243) );
  OR U141 ( .A(n246), .B(n247), .Z(n245) );
  NAND U142 ( .A(n247), .B(n246), .Z(n242) );
  AND U143 ( .A(A[20]), .B(B[11]), .Z(n100) );
  XNOR U144 ( .A(n104), .B(n248), .Z(n101) );
  XNOR U145 ( .A(n103), .B(n102), .Z(n248) );
  AND U146 ( .A(n249), .B(n250), .Z(n102) );
  NANDN U147 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U148 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U149 ( .A(n254), .B(n253), .Z(n249) );
  AND U150 ( .A(A[19]), .B(B[12]), .Z(n103) );
  XNOR U151 ( .A(n107), .B(n255), .Z(n104) );
  XNOR U152 ( .A(n106), .B(n105), .Z(n255) );
  AND U153 ( .A(n256), .B(n257), .Z(n105) );
  NANDN U154 ( .A(n258), .B(n259), .Z(n257) );
  OR U155 ( .A(n260), .B(n261), .Z(n259) );
  NAND U156 ( .A(n261), .B(n260), .Z(n256) );
  AND U157 ( .A(A[18]), .B(B[13]), .Z(n106) );
  XNOR U158 ( .A(n110), .B(n262), .Z(n107) );
  XNOR U159 ( .A(n109), .B(n108), .Z(n262) );
  AND U160 ( .A(n263), .B(n264), .Z(n108) );
  NANDN U161 ( .A(n265), .B(n266), .Z(n264) );
  NANDN U162 ( .A(n267), .B(n268), .Z(n266) );
  NANDN U163 ( .A(n268), .B(n267), .Z(n263) );
  AND U164 ( .A(A[17]), .B(B[14]), .Z(n109) );
  XNOR U165 ( .A(n113), .B(n269), .Z(n110) );
  XNOR U166 ( .A(n112), .B(n111), .Z(n269) );
  AND U167 ( .A(n270), .B(n271), .Z(n111) );
  NANDN U168 ( .A(n272), .B(n273), .Z(n271) );
  OR U169 ( .A(n274), .B(n275), .Z(n273) );
  NAND U170 ( .A(n275), .B(n274), .Z(n270) );
  AND U171 ( .A(A[16]), .B(B[15]), .Z(n112) );
  XNOR U172 ( .A(n116), .B(n276), .Z(n113) );
  XNOR U173 ( .A(n115), .B(n114), .Z(n276) );
  AND U174 ( .A(n277), .B(n278), .Z(n114) );
  NANDN U175 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U176 ( .A(n281), .B(n282), .Z(n280) );
  NANDN U177 ( .A(n282), .B(n281), .Z(n277) );
  AND U178 ( .A(A[15]), .B(B[16]), .Z(n115) );
  XNOR U179 ( .A(n119), .B(n283), .Z(n116) );
  XNOR U180 ( .A(n118), .B(n117), .Z(n283) );
  AND U181 ( .A(n284), .B(n285), .Z(n117) );
  NANDN U182 ( .A(n286), .B(n287), .Z(n285) );
  OR U183 ( .A(n288), .B(n289), .Z(n287) );
  NAND U184 ( .A(n289), .B(n288), .Z(n284) );
  AND U185 ( .A(A[14]), .B(B[17]), .Z(n118) );
  XNOR U186 ( .A(n122), .B(n290), .Z(n119) );
  XNOR U187 ( .A(n121), .B(n120), .Z(n290) );
  AND U188 ( .A(n291), .B(n292), .Z(n120) );
  NANDN U189 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U190 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U191 ( .A(n296), .B(n295), .Z(n291) );
  AND U192 ( .A(A[13]), .B(B[18]), .Z(n121) );
  XNOR U193 ( .A(n125), .B(n297), .Z(n122) );
  XNOR U194 ( .A(n124), .B(n123), .Z(n297) );
  AND U195 ( .A(n298), .B(n299), .Z(n123) );
  NANDN U196 ( .A(n300), .B(n301), .Z(n299) );
  OR U197 ( .A(n302), .B(n303), .Z(n301) );
  NAND U198 ( .A(n303), .B(n302), .Z(n298) );
  AND U199 ( .A(A[12]), .B(B[19]), .Z(n124) );
  XNOR U200 ( .A(n128), .B(n304), .Z(n125) );
  XNOR U201 ( .A(n127), .B(n126), .Z(n304) );
  AND U202 ( .A(n305), .B(n306), .Z(n126) );
  NANDN U203 ( .A(n307), .B(n308), .Z(n306) );
  NANDN U204 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U205 ( .A(n310), .B(n309), .Z(n305) );
  AND U206 ( .A(A[11]), .B(B[20]), .Z(n127) );
  XNOR U207 ( .A(n131), .B(n311), .Z(n128) );
  XNOR U208 ( .A(n130), .B(n129), .Z(n311) );
  AND U209 ( .A(n312), .B(n313), .Z(n129) );
  NANDN U210 ( .A(n314), .B(n315), .Z(n313) );
  OR U211 ( .A(n316), .B(n317), .Z(n315) );
  NAND U212 ( .A(n317), .B(n316), .Z(n312) );
  AND U213 ( .A(A[10]), .B(B[21]), .Z(n130) );
  XNOR U214 ( .A(n134), .B(n318), .Z(n131) );
  XNOR U215 ( .A(n133), .B(n132), .Z(n318) );
  AND U216 ( .A(n319), .B(n320), .Z(n132) );
  NANDN U217 ( .A(n321), .B(n322), .Z(n320) );
  NANDN U218 ( .A(n323), .B(n324), .Z(n322) );
  NANDN U219 ( .A(n324), .B(n323), .Z(n319) );
  AND U220 ( .A(A[9]), .B(B[22]), .Z(n133) );
  XNOR U221 ( .A(n137), .B(n325), .Z(n134) );
  XNOR U222 ( .A(n136), .B(n135), .Z(n325) );
  AND U223 ( .A(n326), .B(n327), .Z(n135) );
  NANDN U224 ( .A(n328), .B(n329), .Z(n327) );
  OR U225 ( .A(n330), .B(n331), .Z(n329) );
  NAND U226 ( .A(n331), .B(n330), .Z(n326) );
  AND U227 ( .A(A[8]), .B(B[23]), .Z(n136) );
  XNOR U228 ( .A(n140), .B(n332), .Z(n137) );
  XNOR U229 ( .A(n139), .B(n138), .Z(n332) );
  AND U230 ( .A(n333), .B(n334), .Z(n138) );
  NANDN U231 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U232 ( .A(n337), .B(n338), .Z(n336) );
  NANDN U233 ( .A(n338), .B(n337), .Z(n333) );
  AND U234 ( .A(A[7]), .B(B[24]), .Z(n139) );
  XNOR U235 ( .A(n143), .B(n339), .Z(n140) );
  XNOR U236 ( .A(n142), .B(n141), .Z(n339) );
  AND U237 ( .A(n340), .B(n341), .Z(n141) );
  NANDN U238 ( .A(n342), .B(n343), .Z(n341) );
  OR U239 ( .A(n344), .B(n345), .Z(n343) );
  NAND U240 ( .A(n345), .B(n344), .Z(n340) );
  AND U241 ( .A(A[6]), .B(B[25]), .Z(n142) );
  XNOR U242 ( .A(n146), .B(n346), .Z(n143) );
  XNOR U243 ( .A(n145), .B(n144), .Z(n346) );
  AND U244 ( .A(n347), .B(n348), .Z(n144) );
  NANDN U245 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U246 ( .A(n351), .B(n352), .Z(n350) );
  NANDN U247 ( .A(n352), .B(n351), .Z(n347) );
  AND U248 ( .A(A[5]), .B(B[26]), .Z(n145) );
  XNOR U249 ( .A(n149), .B(n353), .Z(n146) );
  XNOR U250 ( .A(n148), .B(n147), .Z(n353) );
  AND U251 ( .A(n354), .B(n355), .Z(n147) );
  NANDN U252 ( .A(n356), .B(n357), .Z(n355) );
  OR U253 ( .A(n358), .B(n359), .Z(n357) );
  NAND U254 ( .A(n359), .B(n358), .Z(n354) );
  AND U255 ( .A(A[4]), .B(B[27]), .Z(n148) );
  XNOR U256 ( .A(n152), .B(n360), .Z(n149) );
  XNOR U257 ( .A(n151), .B(n150), .Z(n360) );
  AND U258 ( .A(n361), .B(n362), .Z(n150) );
  NANDN U259 ( .A(n363), .B(n364), .Z(n362) );
  NAND U260 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U261 ( .A(n366), .B(n12), .Z(n361) );
  AND U262 ( .A(A[3]), .B(B[28]), .Z(n151) );
  XOR U263 ( .A(n154), .B(n367), .Z(n152) );
  XNOR U264 ( .A(n153), .B(n155), .Z(n367) );
  NAND U265 ( .A(A[2]), .B(B[29]), .Z(n155) );
  NANDN U266 ( .A(n368), .B(n369), .Z(n153) );
  AND U267 ( .A(A[0]), .B(B[30]), .Z(n369) );
  XNOR U268 ( .A(n156), .B(n370), .Z(n154) );
  NAND U269 ( .A(B[31]), .B(A[0]), .Z(n370) );
  NAND U270 ( .A(B[30]), .B(A[1]), .Z(n156) );
  XOR U271 ( .A(n170), .B(n371), .Z(PRODUCT[30]) );
  XNOR U272 ( .A(n169), .B(n168), .Z(n371) );
  NAND U273 ( .A(n372), .B(n373), .Z(n168) );
  NANDN U274 ( .A(n374), .B(n375), .Z(n373) );
  OR U275 ( .A(n376), .B(n377), .Z(n375) );
  NAND U276 ( .A(n377), .B(n376), .Z(n372) );
  ANDN U277 ( .B(A[30]), .A(n42), .Z(n169) );
  XNOR U278 ( .A(n177), .B(n378), .Z(n170) );
  XNOR U279 ( .A(n176), .B(n174), .Z(n378) );
  AND U280 ( .A(n379), .B(n380), .Z(n174) );
  NANDN U281 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U282 ( .A(n383), .B(n384), .Z(n382) );
  NANDN U283 ( .A(n384), .B(n383), .Z(n379) );
  ANDN U284 ( .B(A[29]), .A(n41), .Z(n176) );
  XNOR U285 ( .A(n184), .B(n385), .Z(n177) );
  XNOR U286 ( .A(n183), .B(n181), .Z(n385) );
  AND U287 ( .A(n386), .B(n387), .Z(n181) );
  NANDN U288 ( .A(n388), .B(n389), .Z(n387) );
  OR U289 ( .A(n390), .B(n391), .Z(n389) );
  NAND U290 ( .A(n391), .B(n390), .Z(n386) );
  AND U291 ( .A(A[28]), .B(B[2]), .Z(n183) );
  XNOR U292 ( .A(n191), .B(n392), .Z(n184) );
  XNOR U293 ( .A(n190), .B(n188), .Z(n392) );
  AND U294 ( .A(n393), .B(n394), .Z(n188) );
  NANDN U295 ( .A(n395), .B(n396), .Z(n394) );
  NANDN U296 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U297 ( .A(n398), .B(n397), .Z(n393) );
  AND U298 ( .A(A[27]), .B(B[3]), .Z(n190) );
  XNOR U299 ( .A(n198), .B(n399), .Z(n191) );
  XNOR U300 ( .A(n197), .B(n195), .Z(n399) );
  AND U301 ( .A(n400), .B(n401), .Z(n195) );
  NANDN U302 ( .A(n402), .B(n403), .Z(n401) );
  OR U303 ( .A(n404), .B(n405), .Z(n403) );
  NAND U304 ( .A(n405), .B(n404), .Z(n400) );
  AND U305 ( .A(A[26]), .B(B[4]), .Z(n197) );
  XNOR U306 ( .A(n205), .B(n406), .Z(n198) );
  XNOR U307 ( .A(n204), .B(n202), .Z(n406) );
  AND U308 ( .A(n407), .B(n408), .Z(n202) );
  NANDN U309 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U310 ( .A(n411), .B(n412), .Z(n410) );
  NANDN U311 ( .A(n412), .B(n411), .Z(n407) );
  AND U312 ( .A(A[25]), .B(B[5]), .Z(n204) );
  XNOR U313 ( .A(n212), .B(n413), .Z(n205) );
  XNOR U314 ( .A(n211), .B(n209), .Z(n413) );
  AND U315 ( .A(n414), .B(n415), .Z(n209) );
  NANDN U316 ( .A(n416), .B(n417), .Z(n415) );
  OR U317 ( .A(n418), .B(n419), .Z(n417) );
  NAND U318 ( .A(n419), .B(n418), .Z(n414) );
  AND U319 ( .A(A[24]), .B(B[6]), .Z(n211) );
  XNOR U320 ( .A(n219), .B(n420), .Z(n212) );
  XNOR U321 ( .A(n218), .B(n216), .Z(n420) );
  AND U322 ( .A(n421), .B(n422), .Z(n216) );
  NANDN U323 ( .A(n423), .B(n424), .Z(n422) );
  NANDN U324 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U325 ( .A(n426), .B(n425), .Z(n421) );
  AND U326 ( .A(A[23]), .B(B[7]), .Z(n218) );
  XNOR U327 ( .A(n226), .B(n427), .Z(n219) );
  XNOR U328 ( .A(n225), .B(n223), .Z(n427) );
  AND U329 ( .A(n428), .B(n429), .Z(n223) );
  NANDN U330 ( .A(n430), .B(n431), .Z(n429) );
  OR U331 ( .A(n432), .B(n433), .Z(n431) );
  NAND U332 ( .A(n433), .B(n432), .Z(n428) );
  AND U333 ( .A(A[22]), .B(B[8]), .Z(n225) );
  XNOR U334 ( .A(n233), .B(n434), .Z(n226) );
  XNOR U335 ( .A(n232), .B(n230), .Z(n434) );
  AND U336 ( .A(n435), .B(n436), .Z(n230) );
  NANDN U337 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U338 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U339 ( .A(n440), .B(n439), .Z(n435) );
  AND U340 ( .A(A[21]), .B(B[9]), .Z(n232) );
  XNOR U341 ( .A(n240), .B(n441), .Z(n233) );
  XNOR U342 ( .A(n239), .B(n237), .Z(n441) );
  AND U343 ( .A(n442), .B(n443), .Z(n237) );
  NANDN U344 ( .A(n444), .B(n445), .Z(n443) );
  OR U345 ( .A(n446), .B(n447), .Z(n445) );
  NAND U346 ( .A(n447), .B(n446), .Z(n442) );
  AND U347 ( .A(A[20]), .B(B[10]), .Z(n239) );
  XNOR U348 ( .A(n247), .B(n448), .Z(n240) );
  XNOR U349 ( .A(n246), .B(n244), .Z(n448) );
  AND U350 ( .A(n449), .B(n450), .Z(n244) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U352 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U353 ( .A(n454), .B(n453), .Z(n449) );
  AND U354 ( .A(A[19]), .B(B[11]), .Z(n246) );
  XNOR U355 ( .A(n254), .B(n455), .Z(n247) );
  XNOR U356 ( .A(n253), .B(n251), .Z(n455) );
  AND U357 ( .A(n456), .B(n457), .Z(n251) );
  NANDN U358 ( .A(n458), .B(n459), .Z(n457) );
  OR U359 ( .A(n460), .B(n461), .Z(n459) );
  NAND U360 ( .A(n461), .B(n460), .Z(n456) );
  AND U361 ( .A(A[18]), .B(B[12]), .Z(n253) );
  XNOR U362 ( .A(n261), .B(n462), .Z(n254) );
  XNOR U363 ( .A(n260), .B(n258), .Z(n462) );
  AND U364 ( .A(n463), .B(n464), .Z(n258) );
  NANDN U365 ( .A(n465), .B(n466), .Z(n464) );
  NANDN U366 ( .A(n467), .B(n468), .Z(n466) );
  NANDN U367 ( .A(n468), .B(n467), .Z(n463) );
  AND U368 ( .A(A[17]), .B(B[13]), .Z(n260) );
  XNOR U369 ( .A(n268), .B(n469), .Z(n261) );
  XNOR U370 ( .A(n267), .B(n265), .Z(n469) );
  AND U371 ( .A(n470), .B(n471), .Z(n265) );
  NANDN U372 ( .A(n472), .B(n473), .Z(n471) );
  OR U373 ( .A(n474), .B(n475), .Z(n473) );
  NAND U374 ( .A(n475), .B(n474), .Z(n470) );
  AND U375 ( .A(A[16]), .B(B[14]), .Z(n267) );
  XNOR U376 ( .A(n275), .B(n476), .Z(n268) );
  XNOR U377 ( .A(n274), .B(n272), .Z(n476) );
  AND U378 ( .A(n477), .B(n478), .Z(n272) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n482), .B(n481), .Z(n477) );
  AND U382 ( .A(A[15]), .B(B[15]), .Z(n274) );
  XNOR U383 ( .A(n282), .B(n483), .Z(n275) );
  XNOR U384 ( .A(n281), .B(n279), .Z(n483) );
  AND U385 ( .A(n484), .B(n485), .Z(n279) );
  NANDN U386 ( .A(n486), .B(n487), .Z(n485) );
  OR U387 ( .A(n488), .B(n489), .Z(n487) );
  NAND U388 ( .A(n489), .B(n488), .Z(n484) );
  AND U389 ( .A(A[14]), .B(B[16]), .Z(n281) );
  XNOR U390 ( .A(n289), .B(n490), .Z(n282) );
  XNOR U391 ( .A(n288), .B(n286), .Z(n490) );
  AND U392 ( .A(n491), .B(n492), .Z(n286) );
  NANDN U393 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U394 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U395 ( .A(n496), .B(n495), .Z(n491) );
  AND U396 ( .A(A[13]), .B(B[17]), .Z(n288) );
  XNOR U397 ( .A(n296), .B(n497), .Z(n289) );
  XNOR U398 ( .A(n295), .B(n293), .Z(n497) );
  AND U399 ( .A(n498), .B(n499), .Z(n293) );
  NANDN U400 ( .A(n500), .B(n501), .Z(n499) );
  OR U401 ( .A(n502), .B(n503), .Z(n501) );
  NAND U402 ( .A(n503), .B(n502), .Z(n498) );
  AND U403 ( .A(A[12]), .B(B[18]), .Z(n295) );
  XNOR U404 ( .A(n303), .B(n504), .Z(n296) );
  XNOR U405 ( .A(n302), .B(n300), .Z(n504) );
  AND U406 ( .A(n505), .B(n506), .Z(n300) );
  NANDN U407 ( .A(n507), .B(n508), .Z(n506) );
  NANDN U408 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U409 ( .A(n510), .B(n509), .Z(n505) );
  AND U410 ( .A(A[11]), .B(B[19]), .Z(n302) );
  XNOR U411 ( .A(n310), .B(n511), .Z(n303) );
  XNOR U412 ( .A(n309), .B(n307), .Z(n511) );
  AND U413 ( .A(n512), .B(n513), .Z(n307) );
  NANDN U414 ( .A(n514), .B(n515), .Z(n513) );
  OR U415 ( .A(n516), .B(n517), .Z(n515) );
  NAND U416 ( .A(n517), .B(n516), .Z(n512) );
  AND U417 ( .A(A[10]), .B(B[20]), .Z(n309) );
  XNOR U418 ( .A(n317), .B(n518), .Z(n310) );
  XNOR U419 ( .A(n316), .B(n314), .Z(n518) );
  AND U420 ( .A(n519), .B(n520), .Z(n314) );
  NANDN U421 ( .A(n521), .B(n522), .Z(n520) );
  NANDN U422 ( .A(n523), .B(n524), .Z(n522) );
  NANDN U423 ( .A(n524), .B(n523), .Z(n519) );
  AND U424 ( .A(A[9]), .B(B[21]), .Z(n316) );
  XNOR U425 ( .A(n324), .B(n525), .Z(n317) );
  XNOR U426 ( .A(n323), .B(n321), .Z(n525) );
  AND U427 ( .A(n526), .B(n527), .Z(n321) );
  NANDN U428 ( .A(n528), .B(n529), .Z(n527) );
  OR U429 ( .A(n530), .B(n531), .Z(n529) );
  NAND U430 ( .A(n531), .B(n530), .Z(n526) );
  AND U431 ( .A(A[8]), .B(B[22]), .Z(n323) );
  XNOR U432 ( .A(n331), .B(n532), .Z(n324) );
  XNOR U433 ( .A(n330), .B(n328), .Z(n532) );
  AND U434 ( .A(n533), .B(n534), .Z(n328) );
  NANDN U435 ( .A(n535), .B(n536), .Z(n534) );
  NANDN U436 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U437 ( .A(n538), .B(n537), .Z(n533) );
  AND U438 ( .A(A[7]), .B(B[23]), .Z(n330) );
  XNOR U439 ( .A(n338), .B(n539), .Z(n331) );
  XNOR U440 ( .A(n337), .B(n335), .Z(n539) );
  AND U441 ( .A(n540), .B(n541), .Z(n335) );
  NANDN U442 ( .A(n542), .B(n543), .Z(n541) );
  OR U443 ( .A(n544), .B(n545), .Z(n543) );
  NAND U444 ( .A(n545), .B(n544), .Z(n540) );
  AND U445 ( .A(A[6]), .B(B[24]), .Z(n337) );
  XNOR U446 ( .A(n345), .B(n546), .Z(n338) );
  XNOR U447 ( .A(n344), .B(n342), .Z(n546) );
  AND U448 ( .A(n547), .B(n548), .Z(n342) );
  NANDN U449 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U450 ( .A(n551), .B(n552), .Z(n550) );
  NANDN U451 ( .A(n552), .B(n551), .Z(n547) );
  AND U452 ( .A(A[5]), .B(B[25]), .Z(n344) );
  XNOR U453 ( .A(n352), .B(n553), .Z(n345) );
  XNOR U454 ( .A(n351), .B(n349), .Z(n553) );
  AND U455 ( .A(n554), .B(n555), .Z(n349) );
  NANDN U456 ( .A(n556), .B(n557), .Z(n555) );
  OR U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n559), .B(n558), .Z(n554) );
  AND U459 ( .A(A[4]), .B(B[26]), .Z(n351) );
  XNOR U460 ( .A(n359), .B(n560), .Z(n352) );
  XNOR U461 ( .A(n358), .B(n356), .Z(n560) );
  AND U462 ( .A(n561), .B(n562), .Z(n356) );
  NANDN U463 ( .A(n563), .B(n564), .Z(n562) );
  NAND U464 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U465 ( .A(n566), .B(n13), .Z(n561) );
  AND U466 ( .A(A[3]), .B(B[27]), .Z(n358) );
  XOR U467 ( .A(n365), .B(n567), .Z(n359) );
  XNOR U468 ( .A(n363), .B(n366), .Z(n567) );
  NAND U469 ( .A(A[2]), .B(B[28]), .Z(n366) );
  NANDN U470 ( .A(n568), .B(n569), .Z(n363) );
  AND U471 ( .A(A[0]), .B(B[29]), .Z(n569) );
  XNOR U472 ( .A(n368), .B(n570), .Z(n365) );
  NAND U473 ( .A(B[30]), .B(A[0]), .Z(n570) );
  NAND U474 ( .A(B[29]), .B(A[1]), .Z(n368) );
  XOR U475 ( .A(n377), .B(n571), .Z(PRODUCT[29]) );
  XNOR U476 ( .A(n376), .B(n374), .Z(n571) );
  AND U477 ( .A(n572), .B(n573), .Z(n374) );
  NAND U478 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U479 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U480 ( .A(n577), .B(n576), .Z(n572) );
  ANDN U481 ( .B(A[29]), .A(n42), .Z(n376) );
  XNOR U482 ( .A(n384), .B(n578), .Z(n377) );
  XNOR U483 ( .A(n383), .B(n381), .Z(n578) );
  AND U484 ( .A(n579), .B(n580), .Z(n381) );
  NANDN U485 ( .A(n581), .B(n582), .Z(n580) );
  OR U486 ( .A(n583), .B(n584), .Z(n582) );
  NAND U487 ( .A(n584), .B(n583), .Z(n579) );
  ANDN U488 ( .B(A[28]), .A(n41), .Z(n383) );
  XNOR U489 ( .A(n391), .B(n585), .Z(n384) );
  XNOR U490 ( .A(n390), .B(n388), .Z(n585) );
  AND U491 ( .A(n586), .B(n587), .Z(n388) );
  NANDN U492 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U493 ( .A(n590), .B(n591), .Z(n589) );
  NANDN U494 ( .A(n591), .B(n590), .Z(n586) );
  AND U495 ( .A(A[27]), .B(B[2]), .Z(n390) );
  XNOR U496 ( .A(n398), .B(n592), .Z(n391) );
  XNOR U497 ( .A(n397), .B(n395), .Z(n592) );
  AND U498 ( .A(n593), .B(n594), .Z(n395) );
  NANDN U499 ( .A(n595), .B(n596), .Z(n594) );
  OR U500 ( .A(n597), .B(n598), .Z(n596) );
  NAND U501 ( .A(n598), .B(n597), .Z(n593) );
  AND U502 ( .A(A[26]), .B(B[3]), .Z(n397) );
  XNOR U503 ( .A(n405), .B(n599), .Z(n398) );
  XNOR U504 ( .A(n404), .B(n402), .Z(n599) );
  AND U505 ( .A(n600), .B(n601), .Z(n402) );
  NANDN U506 ( .A(n602), .B(n603), .Z(n601) );
  NANDN U507 ( .A(n604), .B(n605), .Z(n603) );
  NANDN U508 ( .A(n605), .B(n604), .Z(n600) );
  AND U509 ( .A(A[25]), .B(B[4]), .Z(n404) );
  XNOR U510 ( .A(n412), .B(n606), .Z(n405) );
  XNOR U511 ( .A(n411), .B(n409), .Z(n606) );
  AND U512 ( .A(n607), .B(n608), .Z(n409) );
  NANDN U513 ( .A(n609), .B(n610), .Z(n608) );
  OR U514 ( .A(n611), .B(n612), .Z(n610) );
  NAND U515 ( .A(n612), .B(n611), .Z(n607) );
  AND U516 ( .A(A[24]), .B(B[5]), .Z(n411) );
  XNOR U517 ( .A(n419), .B(n613), .Z(n412) );
  XNOR U518 ( .A(n418), .B(n416), .Z(n613) );
  AND U519 ( .A(n614), .B(n615), .Z(n416) );
  NANDN U520 ( .A(n616), .B(n617), .Z(n615) );
  NANDN U521 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U522 ( .A(n619), .B(n618), .Z(n614) );
  AND U523 ( .A(A[23]), .B(B[6]), .Z(n418) );
  XNOR U524 ( .A(n426), .B(n620), .Z(n419) );
  XNOR U525 ( .A(n425), .B(n423), .Z(n620) );
  AND U526 ( .A(n621), .B(n622), .Z(n423) );
  NANDN U527 ( .A(n623), .B(n624), .Z(n622) );
  OR U528 ( .A(n625), .B(n626), .Z(n624) );
  NAND U529 ( .A(n626), .B(n625), .Z(n621) );
  AND U530 ( .A(A[22]), .B(B[7]), .Z(n425) );
  XNOR U531 ( .A(n433), .B(n627), .Z(n426) );
  XNOR U532 ( .A(n432), .B(n430), .Z(n627) );
  AND U533 ( .A(n628), .B(n629), .Z(n430) );
  NANDN U534 ( .A(n630), .B(n631), .Z(n629) );
  NANDN U535 ( .A(n632), .B(n633), .Z(n631) );
  NANDN U536 ( .A(n633), .B(n632), .Z(n628) );
  AND U537 ( .A(A[21]), .B(B[8]), .Z(n432) );
  XNOR U538 ( .A(n440), .B(n634), .Z(n433) );
  XNOR U539 ( .A(n439), .B(n437), .Z(n634) );
  AND U540 ( .A(n635), .B(n636), .Z(n437) );
  NANDN U541 ( .A(n637), .B(n638), .Z(n636) );
  OR U542 ( .A(n639), .B(n640), .Z(n638) );
  NAND U543 ( .A(n640), .B(n639), .Z(n635) );
  AND U544 ( .A(A[20]), .B(B[9]), .Z(n439) );
  XNOR U545 ( .A(n447), .B(n641), .Z(n440) );
  XNOR U546 ( .A(n446), .B(n444), .Z(n641) );
  AND U547 ( .A(n642), .B(n643), .Z(n444) );
  NANDN U548 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U549 ( .A(n646), .B(n647), .Z(n645) );
  NANDN U550 ( .A(n647), .B(n646), .Z(n642) );
  AND U551 ( .A(A[19]), .B(B[10]), .Z(n446) );
  XNOR U552 ( .A(n454), .B(n648), .Z(n447) );
  XNOR U553 ( .A(n453), .B(n451), .Z(n648) );
  AND U554 ( .A(n649), .B(n650), .Z(n451) );
  NANDN U555 ( .A(n651), .B(n652), .Z(n650) );
  OR U556 ( .A(n653), .B(n654), .Z(n652) );
  NAND U557 ( .A(n654), .B(n653), .Z(n649) );
  AND U558 ( .A(A[18]), .B(B[11]), .Z(n453) );
  XNOR U559 ( .A(n461), .B(n655), .Z(n454) );
  XNOR U560 ( .A(n460), .B(n458), .Z(n655) );
  AND U561 ( .A(n656), .B(n657), .Z(n458) );
  NANDN U562 ( .A(n658), .B(n659), .Z(n657) );
  NANDN U563 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U564 ( .A(n661), .B(n660), .Z(n656) );
  AND U565 ( .A(A[17]), .B(B[12]), .Z(n460) );
  XNOR U566 ( .A(n468), .B(n662), .Z(n461) );
  XNOR U567 ( .A(n467), .B(n465), .Z(n662) );
  AND U568 ( .A(n663), .B(n664), .Z(n465) );
  NANDN U569 ( .A(n665), .B(n666), .Z(n664) );
  OR U570 ( .A(n667), .B(n668), .Z(n666) );
  NAND U571 ( .A(n668), .B(n667), .Z(n663) );
  AND U572 ( .A(A[16]), .B(B[13]), .Z(n467) );
  XNOR U573 ( .A(n475), .B(n669), .Z(n468) );
  XNOR U574 ( .A(n474), .B(n472), .Z(n669) );
  AND U575 ( .A(n670), .B(n671), .Z(n472) );
  NANDN U576 ( .A(n672), .B(n673), .Z(n671) );
  NANDN U577 ( .A(n674), .B(n675), .Z(n673) );
  NANDN U578 ( .A(n675), .B(n674), .Z(n670) );
  AND U579 ( .A(A[15]), .B(B[14]), .Z(n474) );
  XNOR U580 ( .A(n482), .B(n676), .Z(n475) );
  XNOR U581 ( .A(n481), .B(n479), .Z(n676) );
  AND U582 ( .A(n677), .B(n678), .Z(n479) );
  NANDN U583 ( .A(n679), .B(n680), .Z(n678) );
  OR U584 ( .A(n681), .B(n682), .Z(n680) );
  NAND U585 ( .A(n682), .B(n681), .Z(n677) );
  AND U586 ( .A(A[14]), .B(B[15]), .Z(n481) );
  XNOR U587 ( .A(n489), .B(n683), .Z(n482) );
  XNOR U588 ( .A(n488), .B(n486), .Z(n683) );
  AND U589 ( .A(n684), .B(n685), .Z(n486) );
  NANDN U590 ( .A(n686), .B(n687), .Z(n685) );
  NANDN U591 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U592 ( .A(n689), .B(n688), .Z(n684) );
  AND U593 ( .A(A[13]), .B(B[16]), .Z(n488) );
  XNOR U594 ( .A(n496), .B(n690), .Z(n489) );
  XNOR U595 ( .A(n495), .B(n493), .Z(n690) );
  AND U596 ( .A(n691), .B(n692), .Z(n493) );
  NANDN U597 ( .A(n693), .B(n694), .Z(n692) );
  OR U598 ( .A(n695), .B(n696), .Z(n694) );
  NAND U599 ( .A(n696), .B(n695), .Z(n691) );
  AND U600 ( .A(A[12]), .B(B[17]), .Z(n495) );
  XNOR U601 ( .A(n503), .B(n697), .Z(n496) );
  XNOR U602 ( .A(n502), .B(n500), .Z(n697) );
  AND U603 ( .A(n698), .B(n699), .Z(n500) );
  NANDN U604 ( .A(n700), .B(n701), .Z(n699) );
  NANDN U605 ( .A(n702), .B(n703), .Z(n701) );
  NANDN U606 ( .A(n703), .B(n702), .Z(n698) );
  AND U607 ( .A(A[11]), .B(B[18]), .Z(n502) );
  XNOR U608 ( .A(n510), .B(n704), .Z(n503) );
  XNOR U609 ( .A(n509), .B(n507), .Z(n704) );
  AND U610 ( .A(n705), .B(n706), .Z(n507) );
  NANDN U611 ( .A(n707), .B(n708), .Z(n706) );
  OR U612 ( .A(n709), .B(n710), .Z(n708) );
  NAND U613 ( .A(n710), .B(n709), .Z(n705) );
  AND U614 ( .A(A[10]), .B(B[19]), .Z(n509) );
  XNOR U615 ( .A(n517), .B(n711), .Z(n510) );
  XNOR U616 ( .A(n516), .B(n514), .Z(n711) );
  AND U617 ( .A(n712), .B(n713), .Z(n514) );
  NANDN U618 ( .A(n714), .B(n715), .Z(n713) );
  NANDN U619 ( .A(n716), .B(n717), .Z(n715) );
  NANDN U620 ( .A(n717), .B(n716), .Z(n712) );
  AND U621 ( .A(A[9]), .B(B[20]), .Z(n516) );
  XNOR U622 ( .A(n524), .B(n718), .Z(n517) );
  XNOR U623 ( .A(n523), .B(n521), .Z(n718) );
  AND U624 ( .A(n719), .B(n720), .Z(n521) );
  NANDN U625 ( .A(n721), .B(n722), .Z(n720) );
  OR U626 ( .A(n723), .B(n724), .Z(n722) );
  NAND U627 ( .A(n724), .B(n723), .Z(n719) );
  AND U628 ( .A(A[8]), .B(B[21]), .Z(n523) );
  XNOR U629 ( .A(n531), .B(n725), .Z(n524) );
  XNOR U630 ( .A(n530), .B(n528), .Z(n725) );
  AND U631 ( .A(n726), .B(n727), .Z(n528) );
  NANDN U632 ( .A(n728), .B(n729), .Z(n727) );
  NANDN U633 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U634 ( .A(n731), .B(n730), .Z(n726) );
  AND U635 ( .A(A[7]), .B(B[22]), .Z(n530) );
  XNOR U636 ( .A(n538), .B(n732), .Z(n531) );
  XNOR U637 ( .A(n537), .B(n535), .Z(n732) );
  AND U638 ( .A(n733), .B(n734), .Z(n535) );
  NANDN U639 ( .A(n735), .B(n736), .Z(n734) );
  OR U640 ( .A(n737), .B(n738), .Z(n736) );
  NAND U641 ( .A(n738), .B(n737), .Z(n733) );
  AND U642 ( .A(A[6]), .B(B[23]), .Z(n537) );
  XNOR U643 ( .A(n545), .B(n739), .Z(n538) );
  XNOR U644 ( .A(n544), .B(n542), .Z(n739) );
  AND U645 ( .A(n740), .B(n741), .Z(n542) );
  NANDN U646 ( .A(n742), .B(n743), .Z(n741) );
  NANDN U647 ( .A(n744), .B(n745), .Z(n743) );
  NANDN U648 ( .A(n745), .B(n744), .Z(n740) );
  AND U649 ( .A(A[5]), .B(B[24]), .Z(n544) );
  XNOR U650 ( .A(n552), .B(n746), .Z(n545) );
  XNOR U651 ( .A(n551), .B(n549), .Z(n746) );
  AND U652 ( .A(n747), .B(n748), .Z(n549) );
  NANDN U653 ( .A(n749), .B(n750), .Z(n748) );
  OR U654 ( .A(n751), .B(n752), .Z(n750) );
  NAND U655 ( .A(n752), .B(n751), .Z(n747) );
  AND U656 ( .A(A[4]), .B(B[25]), .Z(n551) );
  XNOR U657 ( .A(n559), .B(n753), .Z(n552) );
  XNOR U658 ( .A(n558), .B(n556), .Z(n753) );
  AND U659 ( .A(n754), .B(n755), .Z(n556) );
  NANDN U660 ( .A(n756), .B(n757), .Z(n755) );
  NAND U661 ( .A(n758), .B(n759), .Z(n757) );
  NANDN U662 ( .A(n759), .B(n14), .Z(n754) );
  AND U663 ( .A(A[3]), .B(B[26]), .Z(n558) );
  XOR U664 ( .A(n565), .B(n760), .Z(n559) );
  XNOR U665 ( .A(n563), .B(n566), .Z(n760) );
  NAND U666 ( .A(A[2]), .B(B[27]), .Z(n566) );
  NANDN U667 ( .A(n761), .B(n762), .Z(n563) );
  AND U668 ( .A(A[0]), .B(B[28]), .Z(n762) );
  XNOR U669 ( .A(n568), .B(n763), .Z(n565) );
  NAND U670 ( .A(A[0]), .B(B[29]), .Z(n763) );
  NAND U671 ( .A(B[28]), .B(A[1]), .Z(n568) );
  XOR U672 ( .A(n577), .B(n764), .Z(PRODUCT[28]) );
  XNOR U673 ( .A(n576), .B(n575), .Z(n764) );
  NAND U674 ( .A(n765), .B(n766), .Z(n575) );
  NANDN U675 ( .A(n767), .B(n768), .Z(n766) );
  OR U676 ( .A(n769), .B(n770), .Z(n768) );
  NAND U677 ( .A(n770), .B(n769), .Z(n765) );
  ANDN U678 ( .B(A[28]), .A(n42), .Z(n576) );
  XNOR U679 ( .A(n584), .B(n771), .Z(n577) );
  XNOR U680 ( .A(n583), .B(n581), .Z(n771) );
  AND U681 ( .A(n772), .B(n773), .Z(n581) );
  NANDN U682 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U683 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U684 ( .A(n777), .B(n776), .Z(n772) );
  ANDN U685 ( .B(A[27]), .A(n41), .Z(n583) );
  XNOR U686 ( .A(n591), .B(n778), .Z(n584) );
  XNOR U687 ( .A(n590), .B(n588), .Z(n778) );
  AND U688 ( .A(n779), .B(n780), .Z(n588) );
  NANDN U689 ( .A(n781), .B(n782), .Z(n780) );
  OR U690 ( .A(n783), .B(n784), .Z(n782) );
  NAND U691 ( .A(n784), .B(n783), .Z(n779) );
  AND U692 ( .A(A[26]), .B(B[2]), .Z(n590) );
  XNOR U693 ( .A(n598), .B(n785), .Z(n591) );
  XNOR U694 ( .A(n597), .B(n595), .Z(n785) );
  AND U695 ( .A(n786), .B(n787), .Z(n595) );
  NANDN U696 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U697 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U698 ( .A(n791), .B(n790), .Z(n786) );
  AND U699 ( .A(A[25]), .B(B[3]), .Z(n597) );
  XNOR U700 ( .A(n605), .B(n792), .Z(n598) );
  XNOR U701 ( .A(n604), .B(n602), .Z(n792) );
  AND U702 ( .A(n793), .B(n794), .Z(n602) );
  NANDN U703 ( .A(n795), .B(n796), .Z(n794) );
  OR U704 ( .A(n797), .B(n798), .Z(n796) );
  NAND U705 ( .A(n798), .B(n797), .Z(n793) );
  AND U706 ( .A(A[24]), .B(B[4]), .Z(n604) );
  XNOR U707 ( .A(n612), .B(n799), .Z(n605) );
  XNOR U708 ( .A(n611), .B(n609), .Z(n799) );
  AND U709 ( .A(n800), .B(n801), .Z(n609) );
  NANDN U710 ( .A(n802), .B(n803), .Z(n801) );
  NANDN U711 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U712 ( .A(n805), .B(n804), .Z(n800) );
  AND U713 ( .A(A[23]), .B(B[5]), .Z(n611) );
  XNOR U714 ( .A(n619), .B(n806), .Z(n612) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n806) );
  AND U716 ( .A(n807), .B(n808), .Z(n616) );
  NANDN U717 ( .A(n809), .B(n810), .Z(n808) );
  OR U718 ( .A(n811), .B(n812), .Z(n810) );
  NAND U719 ( .A(n812), .B(n811), .Z(n807) );
  AND U720 ( .A(A[22]), .B(B[6]), .Z(n618) );
  XNOR U721 ( .A(n626), .B(n813), .Z(n619) );
  XNOR U722 ( .A(n625), .B(n623), .Z(n813) );
  AND U723 ( .A(n814), .B(n815), .Z(n623) );
  NANDN U724 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U725 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U726 ( .A(n819), .B(n818), .Z(n814) );
  AND U727 ( .A(A[21]), .B(B[7]), .Z(n625) );
  XNOR U728 ( .A(n633), .B(n820), .Z(n626) );
  XNOR U729 ( .A(n632), .B(n630), .Z(n820) );
  AND U730 ( .A(n821), .B(n822), .Z(n630) );
  NANDN U731 ( .A(n823), .B(n824), .Z(n822) );
  OR U732 ( .A(n825), .B(n826), .Z(n824) );
  NAND U733 ( .A(n826), .B(n825), .Z(n821) );
  AND U734 ( .A(A[20]), .B(B[8]), .Z(n632) );
  XNOR U735 ( .A(n640), .B(n827), .Z(n633) );
  XNOR U736 ( .A(n639), .B(n637), .Z(n827) );
  AND U737 ( .A(n828), .B(n829), .Z(n637) );
  NANDN U738 ( .A(n830), .B(n831), .Z(n829) );
  NANDN U739 ( .A(n832), .B(n833), .Z(n831) );
  NANDN U740 ( .A(n833), .B(n832), .Z(n828) );
  AND U741 ( .A(A[19]), .B(B[9]), .Z(n639) );
  XNOR U742 ( .A(n647), .B(n834), .Z(n640) );
  XNOR U743 ( .A(n646), .B(n644), .Z(n834) );
  AND U744 ( .A(n835), .B(n836), .Z(n644) );
  NANDN U745 ( .A(n837), .B(n838), .Z(n836) );
  OR U746 ( .A(n839), .B(n840), .Z(n838) );
  NAND U747 ( .A(n840), .B(n839), .Z(n835) );
  AND U748 ( .A(A[18]), .B(B[10]), .Z(n646) );
  XNOR U749 ( .A(n654), .B(n841), .Z(n647) );
  XNOR U750 ( .A(n653), .B(n651), .Z(n841) );
  AND U751 ( .A(n842), .B(n843), .Z(n651) );
  NANDN U752 ( .A(n844), .B(n845), .Z(n843) );
  NANDN U753 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U754 ( .A(n847), .B(n846), .Z(n842) );
  AND U755 ( .A(A[17]), .B(B[11]), .Z(n653) );
  XNOR U756 ( .A(n661), .B(n848), .Z(n654) );
  XNOR U757 ( .A(n660), .B(n658), .Z(n848) );
  AND U758 ( .A(n849), .B(n850), .Z(n658) );
  NANDN U759 ( .A(n851), .B(n852), .Z(n850) );
  OR U760 ( .A(n853), .B(n854), .Z(n852) );
  NAND U761 ( .A(n854), .B(n853), .Z(n849) );
  AND U762 ( .A(A[16]), .B(B[12]), .Z(n660) );
  XNOR U763 ( .A(n668), .B(n855), .Z(n661) );
  XNOR U764 ( .A(n667), .B(n665), .Z(n855) );
  AND U765 ( .A(n856), .B(n857), .Z(n665) );
  NANDN U766 ( .A(n858), .B(n859), .Z(n857) );
  NANDN U767 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U768 ( .A(n861), .B(n860), .Z(n856) );
  AND U769 ( .A(A[15]), .B(B[13]), .Z(n667) );
  XNOR U770 ( .A(n675), .B(n862), .Z(n668) );
  XNOR U771 ( .A(n674), .B(n672), .Z(n862) );
  AND U772 ( .A(n863), .B(n864), .Z(n672) );
  NANDN U773 ( .A(n865), .B(n866), .Z(n864) );
  OR U774 ( .A(n867), .B(n868), .Z(n866) );
  NAND U775 ( .A(n868), .B(n867), .Z(n863) );
  AND U776 ( .A(A[14]), .B(B[14]), .Z(n674) );
  XNOR U777 ( .A(n682), .B(n869), .Z(n675) );
  XNOR U778 ( .A(n681), .B(n679), .Z(n869) );
  AND U779 ( .A(n870), .B(n871), .Z(n679) );
  NANDN U780 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U781 ( .A(n874), .B(n875), .Z(n873) );
  NANDN U782 ( .A(n875), .B(n874), .Z(n870) );
  AND U783 ( .A(A[13]), .B(B[15]), .Z(n681) );
  XNOR U784 ( .A(n689), .B(n876), .Z(n682) );
  XNOR U785 ( .A(n688), .B(n686), .Z(n876) );
  AND U786 ( .A(n877), .B(n878), .Z(n686) );
  NANDN U787 ( .A(n879), .B(n880), .Z(n878) );
  OR U788 ( .A(n881), .B(n882), .Z(n880) );
  NAND U789 ( .A(n882), .B(n881), .Z(n877) );
  AND U790 ( .A(A[12]), .B(B[16]), .Z(n688) );
  XNOR U791 ( .A(n696), .B(n883), .Z(n689) );
  XNOR U792 ( .A(n695), .B(n693), .Z(n883) );
  AND U793 ( .A(n884), .B(n885), .Z(n693) );
  NANDN U794 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U795 ( .A(n888), .B(n889), .Z(n887) );
  NANDN U796 ( .A(n889), .B(n888), .Z(n884) );
  AND U797 ( .A(A[11]), .B(B[17]), .Z(n695) );
  XNOR U798 ( .A(n703), .B(n890), .Z(n696) );
  XNOR U799 ( .A(n702), .B(n700), .Z(n890) );
  AND U800 ( .A(n891), .B(n892), .Z(n700) );
  NANDN U801 ( .A(n893), .B(n894), .Z(n892) );
  OR U802 ( .A(n895), .B(n896), .Z(n894) );
  NAND U803 ( .A(n896), .B(n895), .Z(n891) );
  AND U804 ( .A(A[10]), .B(B[18]), .Z(n702) );
  XNOR U805 ( .A(n710), .B(n897), .Z(n703) );
  XNOR U806 ( .A(n709), .B(n707), .Z(n897) );
  AND U807 ( .A(n898), .B(n899), .Z(n707) );
  NANDN U808 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U809 ( .A(n902), .B(n903), .Z(n901) );
  NANDN U810 ( .A(n903), .B(n902), .Z(n898) );
  AND U811 ( .A(A[9]), .B(B[19]), .Z(n709) );
  XNOR U812 ( .A(n717), .B(n904), .Z(n710) );
  XNOR U813 ( .A(n716), .B(n714), .Z(n904) );
  AND U814 ( .A(n905), .B(n906), .Z(n714) );
  NANDN U815 ( .A(n907), .B(n908), .Z(n906) );
  OR U816 ( .A(n909), .B(n910), .Z(n908) );
  NAND U817 ( .A(n910), .B(n909), .Z(n905) );
  AND U818 ( .A(A[8]), .B(B[20]), .Z(n716) );
  XNOR U819 ( .A(n724), .B(n911), .Z(n717) );
  XNOR U820 ( .A(n723), .B(n721), .Z(n911) );
  AND U821 ( .A(n912), .B(n913), .Z(n721) );
  NANDN U822 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U823 ( .A(n916), .B(n917), .Z(n915) );
  NANDN U824 ( .A(n917), .B(n916), .Z(n912) );
  AND U825 ( .A(A[7]), .B(B[21]), .Z(n723) );
  XNOR U826 ( .A(n731), .B(n918), .Z(n724) );
  XNOR U827 ( .A(n730), .B(n728), .Z(n918) );
  AND U828 ( .A(n919), .B(n920), .Z(n728) );
  NANDN U829 ( .A(n921), .B(n922), .Z(n920) );
  OR U830 ( .A(n923), .B(n924), .Z(n922) );
  NAND U831 ( .A(n924), .B(n923), .Z(n919) );
  AND U832 ( .A(A[6]), .B(B[22]), .Z(n730) );
  XNOR U833 ( .A(n738), .B(n925), .Z(n731) );
  XNOR U834 ( .A(n737), .B(n735), .Z(n925) );
  AND U835 ( .A(n926), .B(n927), .Z(n735) );
  NANDN U836 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U837 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U838 ( .A(n931), .B(n930), .Z(n926) );
  AND U839 ( .A(A[5]), .B(B[23]), .Z(n737) );
  XNOR U840 ( .A(n745), .B(n932), .Z(n738) );
  XNOR U841 ( .A(n744), .B(n742), .Z(n932) );
  AND U842 ( .A(n933), .B(n934), .Z(n742) );
  NANDN U843 ( .A(n935), .B(n936), .Z(n934) );
  OR U844 ( .A(n937), .B(n938), .Z(n936) );
  NAND U845 ( .A(n938), .B(n937), .Z(n933) );
  AND U846 ( .A(A[4]), .B(B[24]), .Z(n744) );
  XNOR U847 ( .A(n752), .B(n939), .Z(n745) );
  XNOR U848 ( .A(n751), .B(n749), .Z(n939) );
  AND U849 ( .A(n940), .B(n941), .Z(n749) );
  NANDN U850 ( .A(n942), .B(n943), .Z(n941) );
  NAND U851 ( .A(n944), .B(n945), .Z(n943) );
  NANDN U852 ( .A(n945), .B(n15), .Z(n940) );
  AND U853 ( .A(A[3]), .B(B[25]), .Z(n751) );
  XOR U854 ( .A(n758), .B(n946), .Z(n752) );
  XNOR U855 ( .A(n756), .B(n759), .Z(n946) );
  NAND U856 ( .A(A[2]), .B(B[26]), .Z(n759) );
  NANDN U857 ( .A(n947), .B(n948), .Z(n756) );
  AND U858 ( .A(A[0]), .B(B[27]), .Z(n948) );
  XNOR U859 ( .A(n761), .B(n949), .Z(n758) );
  NAND U860 ( .A(A[0]), .B(B[28]), .Z(n949) );
  NAND U861 ( .A(B[27]), .B(A[1]), .Z(n761) );
  XOR U862 ( .A(n770), .B(n950), .Z(PRODUCT[27]) );
  XNOR U863 ( .A(n769), .B(n767), .Z(n950) );
  AND U864 ( .A(n951), .B(n952), .Z(n767) );
  NAND U865 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U866 ( .A(n955), .B(n956), .Z(n953) );
  NANDN U867 ( .A(n956), .B(n955), .Z(n951) );
  ANDN U868 ( .B(A[27]), .A(n42), .Z(n769) );
  XNOR U869 ( .A(n777), .B(n957), .Z(n770) );
  XNOR U870 ( .A(n776), .B(n774), .Z(n957) );
  AND U871 ( .A(n958), .B(n959), .Z(n774) );
  NANDN U872 ( .A(n960), .B(n961), .Z(n959) );
  OR U873 ( .A(n962), .B(n963), .Z(n961) );
  NAND U874 ( .A(n963), .B(n962), .Z(n958) );
  ANDN U875 ( .B(A[26]), .A(n41), .Z(n776) );
  XNOR U876 ( .A(n784), .B(n964), .Z(n777) );
  XNOR U877 ( .A(n783), .B(n781), .Z(n964) );
  AND U878 ( .A(n965), .B(n966), .Z(n781) );
  NANDN U879 ( .A(n967), .B(n968), .Z(n966) );
  NANDN U880 ( .A(n969), .B(n970), .Z(n968) );
  NANDN U881 ( .A(n970), .B(n969), .Z(n965) );
  AND U882 ( .A(A[25]), .B(B[2]), .Z(n783) );
  XNOR U883 ( .A(n791), .B(n971), .Z(n784) );
  XNOR U884 ( .A(n790), .B(n788), .Z(n971) );
  AND U885 ( .A(n972), .B(n973), .Z(n788) );
  NANDN U886 ( .A(n974), .B(n975), .Z(n973) );
  OR U887 ( .A(n976), .B(n977), .Z(n975) );
  NAND U888 ( .A(n977), .B(n976), .Z(n972) );
  AND U889 ( .A(A[24]), .B(B[3]), .Z(n790) );
  XNOR U890 ( .A(n798), .B(n978), .Z(n791) );
  XNOR U891 ( .A(n797), .B(n795), .Z(n978) );
  AND U892 ( .A(n979), .B(n980), .Z(n795) );
  NANDN U893 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U894 ( .A(n983), .B(n984), .Z(n982) );
  NANDN U895 ( .A(n984), .B(n983), .Z(n979) );
  AND U896 ( .A(A[23]), .B(B[4]), .Z(n797) );
  XNOR U897 ( .A(n805), .B(n985), .Z(n798) );
  XNOR U898 ( .A(n804), .B(n802), .Z(n985) );
  AND U899 ( .A(n986), .B(n987), .Z(n802) );
  NANDN U900 ( .A(n988), .B(n989), .Z(n987) );
  OR U901 ( .A(n990), .B(n991), .Z(n989) );
  NAND U902 ( .A(n991), .B(n990), .Z(n986) );
  AND U903 ( .A(A[22]), .B(B[5]), .Z(n804) );
  XNOR U904 ( .A(n812), .B(n992), .Z(n805) );
  XNOR U905 ( .A(n811), .B(n809), .Z(n992) );
  AND U906 ( .A(n993), .B(n994), .Z(n809) );
  NANDN U907 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U908 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U909 ( .A(n998), .B(n997), .Z(n993) );
  AND U910 ( .A(A[21]), .B(B[6]), .Z(n811) );
  XNOR U911 ( .A(n819), .B(n999), .Z(n812) );
  XNOR U912 ( .A(n818), .B(n816), .Z(n999) );
  AND U913 ( .A(n1000), .B(n1001), .Z(n816) );
  NANDN U914 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U915 ( .A(n1004), .B(n1005), .Z(n1003) );
  NAND U916 ( .A(n1005), .B(n1004), .Z(n1000) );
  AND U917 ( .A(A[20]), .B(B[7]), .Z(n818) );
  XNOR U918 ( .A(n826), .B(n1006), .Z(n819) );
  XNOR U919 ( .A(n825), .B(n823), .Z(n1006) );
  AND U920 ( .A(n1007), .B(n1008), .Z(n823) );
  NANDN U921 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U922 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U923 ( .A(n1012), .B(n1011), .Z(n1007) );
  AND U924 ( .A(A[19]), .B(B[8]), .Z(n825) );
  XNOR U925 ( .A(n833), .B(n1013), .Z(n826) );
  XNOR U926 ( .A(n832), .B(n830), .Z(n1013) );
  AND U927 ( .A(n1014), .B(n1015), .Z(n830) );
  NANDN U928 ( .A(n1016), .B(n1017), .Z(n1015) );
  OR U929 ( .A(n1018), .B(n1019), .Z(n1017) );
  NAND U930 ( .A(n1019), .B(n1018), .Z(n1014) );
  AND U931 ( .A(A[18]), .B(B[9]), .Z(n832) );
  XNOR U932 ( .A(n840), .B(n1020), .Z(n833) );
  XNOR U933 ( .A(n839), .B(n837), .Z(n1020) );
  AND U934 ( .A(n1021), .B(n1022), .Z(n837) );
  NANDN U935 ( .A(n1023), .B(n1024), .Z(n1022) );
  NANDN U936 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U937 ( .A(n1026), .B(n1025), .Z(n1021) );
  AND U938 ( .A(A[17]), .B(B[10]), .Z(n839) );
  XNOR U939 ( .A(n847), .B(n1027), .Z(n840) );
  XNOR U940 ( .A(n846), .B(n844), .Z(n1027) );
  AND U941 ( .A(n1028), .B(n1029), .Z(n844) );
  NANDN U942 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U943 ( .A(n1032), .B(n1033), .Z(n1031) );
  NAND U944 ( .A(n1033), .B(n1032), .Z(n1028) );
  AND U945 ( .A(A[16]), .B(B[11]), .Z(n846) );
  XNOR U946 ( .A(n854), .B(n1034), .Z(n847) );
  XNOR U947 ( .A(n853), .B(n851), .Z(n1034) );
  AND U948 ( .A(n1035), .B(n1036), .Z(n851) );
  NANDN U949 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U950 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U951 ( .A(n1040), .B(n1039), .Z(n1035) );
  AND U952 ( .A(A[15]), .B(B[12]), .Z(n853) );
  XNOR U953 ( .A(n861), .B(n1041), .Z(n854) );
  XNOR U954 ( .A(n860), .B(n858), .Z(n1041) );
  AND U955 ( .A(n1042), .B(n1043), .Z(n858) );
  NANDN U956 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U957 ( .A(n1046), .B(n1047), .Z(n1045) );
  NAND U958 ( .A(n1047), .B(n1046), .Z(n1042) );
  AND U959 ( .A(A[14]), .B(B[13]), .Z(n860) );
  XNOR U960 ( .A(n868), .B(n1048), .Z(n861) );
  XNOR U961 ( .A(n867), .B(n865), .Z(n1048) );
  AND U962 ( .A(n1049), .B(n1050), .Z(n865) );
  NANDN U963 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U964 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U965 ( .A(n1054), .B(n1053), .Z(n1049) );
  AND U966 ( .A(A[13]), .B(B[14]), .Z(n867) );
  XNOR U967 ( .A(n875), .B(n1055), .Z(n868) );
  XNOR U968 ( .A(n874), .B(n872), .Z(n1055) );
  AND U969 ( .A(n1056), .B(n1057), .Z(n872) );
  NANDN U970 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U971 ( .A(n1060), .B(n1061), .Z(n1059) );
  NAND U972 ( .A(n1061), .B(n1060), .Z(n1056) );
  AND U973 ( .A(A[12]), .B(B[15]), .Z(n874) );
  XNOR U974 ( .A(n882), .B(n1062), .Z(n875) );
  XNOR U975 ( .A(n881), .B(n879), .Z(n1062) );
  AND U976 ( .A(n1063), .B(n1064), .Z(n879) );
  NANDN U977 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U978 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U979 ( .A(n1068), .B(n1067), .Z(n1063) );
  AND U980 ( .A(A[11]), .B(B[16]), .Z(n881) );
  XNOR U981 ( .A(n889), .B(n1069), .Z(n882) );
  XNOR U982 ( .A(n888), .B(n886), .Z(n1069) );
  AND U983 ( .A(n1070), .B(n1071), .Z(n886) );
  NANDN U984 ( .A(n1072), .B(n1073), .Z(n1071) );
  OR U985 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U986 ( .A(n1075), .B(n1074), .Z(n1070) );
  AND U987 ( .A(A[10]), .B(B[17]), .Z(n888) );
  XNOR U988 ( .A(n896), .B(n1076), .Z(n889) );
  XNOR U989 ( .A(n895), .B(n893), .Z(n1076) );
  AND U990 ( .A(n1077), .B(n1078), .Z(n893) );
  NANDN U991 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U992 ( .A(n1081), .B(n1082), .Z(n1080) );
  NANDN U993 ( .A(n1082), .B(n1081), .Z(n1077) );
  AND U994 ( .A(A[9]), .B(B[18]), .Z(n895) );
  XNOR U995 ( .A(n903), .B(n1083), .Z(n896) );
  XNOR U996 ( .A(n902), .B(n900), .Z(n1083) );
  AND U997 ( .A(n1084), .B(n1085), .Z(n900) );
  NANDN U998 ( .A(n1086), .B(n1087), .Z(n1085) );
  OR U999 ( .A(n1088), .B(n1089), .Z(n1087) );
  NAND U1000 ( .A(n1089), .B(n1088), .Z(n1084) );
  AND U1001 ( .A(A[8]), .B(B[19]), .Z(n902) );
  XNOR U1002 ( .A(n910), .B(n1090), .Z(n903) );
  XNOR U1003 ( .A(n909), .B(n907), .Z(n1090) );
  AND U1004 ( .A(n1091), .B(n1092), .Z(n907) );
  NANDN U1005 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1006 ( .A(n1095), .B(n1096), .Z(n1094) );
  NANDN U1007 ( .A(n1096), .B(n1095), .Z(n1091) );
  AND U1008 ( .A(A[7]), .B(B[20]), .Z(n909) );
  XNOR U1009 ( .A(n917), .B(n1097), .Z(n910) );
  XNOR U1010 ( .A(n916), .B(n914), .Z(n1097) );
  AND U1011 ( .A(n1098), .B(n1099), .Z(n914) );
  NANDN U1012 ( .A(n1100), .B(n1101), .Z(n1099) );
  OR U1013 ( .A(n1102), .B(n1103), .Z(n1101) );
  NAND U1014 ( .A(n1103), .B(n1102), .Z(n1098) );
  AND U1015 ( .A(A[6]), .B(B[21]), .Z(n916) );
  XNOR U1016 ( .A(n924), .B(n1104), .Z(n917) );
  XNOR U1017 ( .A(n923), .B(n921), .Z(n1104) );
  AND U1018 ( .A(n1105), .B(n1106), .Z(n921) );
  NANDN U1019 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1020 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U1021 ( .A(n1110), .B(n1109), .Z(n1105) );
  AND U1022 ( .A(A[5]), .B(B[22]), .Z(n923) );
  XNOR U1023 ( .A(n931), .B(n1111), .Z(n924) );
  XNOR U1024 ( .A(n930), .B(n928), .Z(n1111) );
  AND U1025 ( .A(n1112), .B(n1113), .Z(n928) );
  NANDN U1026 ( .A(n1114), .B(n1115), .Z(n1113) );
  OR U1027 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U1028 ( .A(n1117), .B(n1116), .Z(n1112) );
  AND U1029 ( .A(A[4]), .B(B[23]), .Z(n930) );
  XNOR U1030 ( .A(n938), .B(n1118), .Z(n931) );
  XNOR U1031 ( .A(n937), .B(n935), .Z(n1118) );
  AND U1032 ( .A(n1119), .B(n1120), .Z(n935) );
  NANDN U1033 ( .A(n1121), .B(n1122), .Z(n1120) );
  NAND U1034 ( .A(n1123), .B(n1124), .Z(n1122) );
  NANDN U1035 ( .A(n1124), .B(n16), .Z(n1119) );
  AND U1036 ( .A(A[3]), .B(B[24]), .Z(n937) );
  XOR U1037 ( .A(n944), .B(n1125), .Z(n938) );
  XNOR U1038 ( .A(n942), .B(n945), .Z(n1125) );
  NAND U1039 ( .A(A[2]), .B(B[25]), .Z(n945) );
  NANDN U1040 ( .A(n1126), .B(n1127), .Z(n942) );
  AND U1041 ( .A(A[0]), .B(B[26]), .Z(n1127) );
  XNOR U1042 ( .A(n947), .B(n1128), .Z(n944) );
  NAND U1043 ( .A(A[0]), .B(B[27]), .Z(n1128) );
  NAND U1044 ( .A(B[26]), .B(A[1]), .Z(n947) );
  XOR U1045 ( .A(n956), .B(n1129), .Z(PRODUCT[26]) );
  XNOR U1046 ( .A(n955), .B(n954), .Z(n1129) );
  NAND U1047 ( .A(n1130), .B(n1131), .Z(n954) );
  NANDN U1048 ( .A(n1132), .B(n1133), .Z(n1131) );
  OR U1049 ( .A(n1134), .B(n1135), .Z(n1133) );
  NAND U1050 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1051 ( .B(A[26]), .A(n42), .Z(n955) );
  XNOR U1052 ( .A(n963), .B(n1136), .Z(n956) );
  XNOR U1053 ( .A(n962), .B(n960), .Z(n1136) );
  AND U1054 ( .A(n1137), .B(n1138), .Z(n960) );
  NANDN U1055 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1056 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U1057 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1058 ( .B(A[25]), .A(n41), .Z(n962) );
  XNOR U1059 ( .A(n970), .B(n1143), .Z(n963) );
  XNOR U1060 ( .A(n969), .B(n967), .Z(n1143) );
  AND U1061 ( .A(n1144), .B(n1145), .Z(n967) );
  NANDN U1062 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1063 ( .A(n1148), .B(n1149), .Z(n1147) );
  NAND U1064 ( .A(n1149), .B(n1148), .Z(n1144) );
  AND U1065 ( .A(A[24]), .B(B[2]), .Z(n969) );
  XNOR U1066 ( .A(n977), .B(n1150), .Z(n970) );
  XNOR U1067 ( .A(n976), .B(n974), .Z(n1150) );
  AND U1068 ( .A(n1151), .B(n1152), .Z(n974) );
  NANDN U1069 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1070 ( .A(n1155), .B(n1156), .Z(n1154) );
  NANDN U1071 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1072 ( .A(A[23]), .B(B[3]), .Z(n976) );
  XNOR U1073 ( .A(n984), .B(n1157), .Z(n977) );
  XNOR U1074 ( .A(n983), .B(n981), .Z(n1157) );
  AND U1075 ( .A(n1158), .B(n1159), .Z(n981) );
  NANDN U1076 ( .A(n1160), .B(n1161), .Z(n1159) );
  OR U1077 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1078 ( .A(n1163), .B(n1162), .Z(n1158) );
  AND U1079 ( .A(A[22]), .B(B[4]), .Z(n983) );
  XNOR U1080 ( .A(n991), .B(n1164), .Z(n984) );
  XNOR U1081 ( .A(n990), .B(n988), .Z(n1164) );
  AND U1082 ( .A(n1165), .B(n1166), .Z(n988) );
  NANDN U1083 ( .A(n1167), .B(n1168), .Z(n1166) );
  NANDN U1084 ( .A(n1169), .B(n1170), .Z(n1168) );
  NANDN U1085 ( .A(n1170), .B(n1169), .Z(n1165) );
  AND U1086 ( .A(A[21]), .B(B[5]), .Z(n990) );
  XNOR U1087 ( .A(n998), .B(n1171), .Z(n991) );
  XNOR U1088 ( .A(n997), .B(n995), .Z(n1171) );
  AND U1089 ( .A(n1172), .B(n1173), .Z(n995) );
  NANDN U1090 ( .A(n1174), .B(n1175), .Z(n1173) );
  OR U1091 ( .A(n1176), .B(n1177), .Z(n1175) );
  NAND U1092 ( .A(n1177), .B(n1176), .Z(n1172) );
  AND U1093 ( .A(A[20]), .B(B[6]), .Z(n997) );
  XNOR U1094 ( .A(n1005), .B(n1178), .Z(n998) );
  XNOR U1095 ( .A(n1004), .B(n1002), .Z(n1178) );
  AND U1096 ( .A(n1179), .B(n1180), .Z(n1002) );
  NANDN U1097 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1098 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1099 ( .A(n1184), .B(n1183), .Z(n1179) );
  AND U1100 ( .A(A[19]), .B(B[7]), .Z(n1004) );
  XNOR U1101 ( .A(n1012), .B(n1185), .Z(n1005) );
  XNOR U1102 ( .A(n1011), .B(n1009), .Z(n1185) );
  AND U1103 ( .A(n1186), .B(n1187), .Z(n1009) );
  NANDN U1104 ( .A(n1188), .B(n1189), .Z(n1187) );
  OR U1105 ( .A(n1190), .B(n1191), .Z(n1189) );
  NAND U1106 ( .A(n1191), .B(n1190), .Z(n1186) );
  AND U1107 ( .A(A[18]), .B(B[8]), .Z(n1011) );
  XNOR U1108 ( .A(n1019), .B(n1192), .Z(n1012) );
  XNOR U1109 ( .A(n1018), .B(n1016), .Z(n1192) );
  AND U1110 ( .A(n1193), .B(n1194), .Z(n1016) );
  NANDN U1111 ( .A(n1195), .B(n1196), .Z(n1194) );
  NANDN U1112 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1113 ( .A(n1198), .B(n1197), .Z(n1193) );
  AND U1114 ( .A(A[17]), .B(B[9]), .Z(n1018) );
  XNOR U1115 ( .A(n1026), .B(n1199), .Z(n1019) );
  XNOR U1116 ( .A(n1025), .B(n1023), .Z(n1199) );
  AND U1117 ( .A(n1200), .B(n1201), .Z(n1023) );
  NANDN U1118 ( .A(n1202), .B(n1203), .Z(n1201) );
  OR U1119 ( .A(n1204), .B(n1205), .Z(n1203) );
  NAND U1120 ( .A(n1205), .B(n1204), .Z(n1200) );
  AND U1121 ( .A(A[16]), .B(B[10]), .Z(n1025) );
  XNOR U1122 ( .A(n1033), .B(n1206), .Z(n1026) );
  XNOR U1123 ( .A(n1032), .B(n1030), .Z(n1206) );
  AND U1124 ( .A(n1207), .B(n1208), .Z(n1030) );
  NANDN U1125 ( .A(n1209), .B(n1210), .Z(n1208) );
  NANDN U1126 ( .A(n1211), .B(n1212), .Z(n1210) );
  NANDN U1127 ( .A(n1212), .B(n1211), .Z(n1207) );
  AND U1128 ( .A(A[15]), .B(B[11]), .Z(n1032) );
  XNOR U1129 ( .A(n1040), .B(n1213), .Z(n1033) );
  XNOR U1130 ( .A(n1039), .B(n1037), .Z(n1213) );
  AND U1131 ( .A(n1214), .B(n1215), .Z(n1037) );
  NANDN U1132 ( .A(n1216), .B(n1217), .Z(n1215) );
  OR U1133 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1134 ( .A(n1219), .B(n1218), .Z(n1214) );
  AND U1135 ( .A(A[14]), .B(B[12]), .Z(n1039) );
  XNOR U1136 ( .A(n1047), .B(n1220), .Z(n1040) );
  XNOR U1137 ( .A(n1046), .B(n1044), .Z(n1220) );
  AND U1138 ( .A(n1221), .B(n1222), .Z(n1044) );
  NANDN U1139 ( .A(n1223), .B(n1224), .Z(n1222) );
  NANDN U1140 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1141 ( .A(n1226), .B(n1225), .Z(n1221) );
  AND U1142 ( .A(A[13]), .B(B[13]), .Z(n1046) );
  XNOR U1143 ( .A(n1054), .B(n1227), .Z(n1047) );
  XNOR U1144 ( .A(n1053), .B(n1051), .Z(n1227) );
  AND U1145 ( .A(n1228), .B(n1229), .Z(n1051) );
  NANDN U1146 ( .A(n1230), .B(n1231), .Z(n1229) );
  OR U1147 ( .A(n1232), .B(n1233), .Z(n1231) );
  NAND U1148 ( .A(n1233), .B(n1232), .Z(n1228) );
  AND U1149 ( .A(A[12]), .B(B[14]), .Z(n1053) );
  XNOR U1150 ( .A(n1061), .B(n1234), .Z(n1054) );
  XNOR U1151 ( .A(n1060), .B(n1058), .Z(n1234) );
  AND U1152 ( .A(n1235), .B(n1236), .Z(n1058) );
  NANDN U1153 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1154 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1155 ( .A(n1240), .B(n1239), .Z(n1235) );
  AND U1156 ( .A(A[11]), .B(B[15]), .Z(n1060) );
  XNOR U1157 ( .A(n1068), .B(n1241), .Z(n1061) );
  XNOR U1158 ( .A(n1067), .B(n1065), .Z(n1241) );
  AND U1159 ( .A(n1242), .B(n1243), .Z(n1065) );
  NANDN U1160 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U1161 ( .A(n1246), .B(n1247), .Z(n1245) );
  NAND U1162 ( .A(n1247), .B(n1246), .Z(n1242) );
  AND U1163 ( .A(A[10]), .B(B[16]), .Z(n1067) );
  XNOR U1164 ( .A(n1075), .B(n1248), .Z(n1068) );
  XNOR U1165 ( .A(n1074), .B(n1072), .Z(n1248) );
  AND U1166 ( .A(n1249), .B(n1250), .Z(n1072) );
  NANDN U1167 ( .A(n1251), .B(n1252), .Z(n1250) );
  NANDN U1168 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1169 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1170 ( .A(A[9]), .B(B[17]), .Z(n1074) );
  XNOR U1171 ( .A(n1082), .B(n1255), .Z(n1075) );
  XNOR U1172 ( .A(n1081), .B(n1079), .Z(n1255) );
  AND U1173 ( .A(n1256), .B(n1257), .Z(n1079) );
  NANDN U1174 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1175 ( .A(n1260), .B(n1261), .Z(n1259) );
  NAND U1176 ( .A(n1261), .B(n1260), .Z(n1256) );
  AND U1177 ( .A(A[8]), .B(B[18]), .Z(n1081) );
  XNOR U1178 ( .A(n1089), .B(n1262), .Z(n1082) );
  XNOR U1179 ( .A(n1088), .B(n1086), .Z(n1262) );
  AND U1180 ( .A(n1263), .B(n1264), .Z(n1086) );
  NANDN U1181 ( .A(n1265), .B(n1266), .Z(n1264) );
  NANDN U1182 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1183 ( .A(n1268), .B(n1267), .Z(n1263) );
  AND U1184 ( .A(A[7]), .B(B[19]), .Z(n1088) );
  XNOR U1185 ( .A(n1096), .B(n1269), .Z(n1089) );
  XNOR U1186 ( .A(n1095), .B(n1093), .Z(n1269) );
  AND U1187 ( .A(n1270), .B(n1271), .Z(n1093) );
  NANDN U1188 ( .A(n1272), .B(n1273), .Z(n1271) );
  OR U1189 ( .A(n1274), .B(n1275), .Z(n1273) );
  NAND U1190 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1191 ( .A(A[6]), .B(B[20]), .Z(n1095) );
  XNOR U1192 ( .A(n1103), .B(n1276), .Z(n1096) );
  XNOR U1193 ( .A(n1102), .B(n1100), .Z(n1276) );
  AND U1194 ( .A(n1277), .B(n1278), .Z(n1100) );
  NANDN U1195 ( .A(n1279), .B(n1280), .Z(n1278) );
  NANDN U1196 ( .A(n1281), .B(n1282), .Z(n1280) );
  NANDN U1197 ( .A(n1282), .B(n1281), .Z(n1277) );
  AND U1198 ( .A(A[5]), .B(B[21]), .Z(n1102) );
  XNOR U1199 ( .A(n1110), .B(n1283), .Z(n1103) );
  XNOR U1200 ( .A(n1109), .B(n1107), .Z(n1283) );
  AND U1201 ( .A(n1284), .B(n1285), .Z(n1107) );
  NANDN U1202 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1203 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1204 ( .A(n1289), .B(n1288), .Z(n1284) );
  AND U1205 ( .A(A[4]), .B(B[22]), .Z(n1109) );
  XNOR U1206 ( .A(n1117), .B(n1290), .Z(n1110) );
  XNOR U1207 ( .A(n1116), .B(n1114), .Z(n1290) );
  AND U1208 ( .A(n1291), .B(n1292), .Z(n1114) );
  NANDN U1209 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1210 ( .A(n1295), .B(n1296), .Z(n1294) );
  NANDN U1211 ( .A(n1296), .B(n17), .Z(n1291) );
  AND U1212 ( .A(A[3]), .B(B[23]), .Z(n1116) );
  XOR U1213 ( .A(n1123), .B(n1297), .Z(n1117) );
  XNOR U1214 ( .A(n1121), .B(n1124), .Z(n1297) );
  NAND U1215 ( .A(A[2]), .B(B[24]), .Z(n1124) );
  NANDN U1216 ( .A(n1298), .B(n1299), .Z(n1121) );
  AND U1217 ( .A(A[0]), .B(B[25]), .Z(n1299) );
  XNOR U1218 ( .A(n1126), .B(n1300), .Z(n1123) );
  NAND U1219 ( .A(A[0]), .B(B[26]), .Z(n1300) );
  NAND U1220 ( .A(B[25]), .B(A[1]), .Z(n1126) );
  XOR U1221 ( .A(n1135), .B(n1301), .Z(PRODUCT[25]) );
  XNOR U1222 ( .A(n1134), .B(n1132), .Z(n1301) );
  AND U1223 ( .A(n1302), .B(n1303), .Z(n1132) );
  NAND U1224 ( .A(n1304), .B(n1305), .Z(n1303) );
  NANDN U1225 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U1226 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1227 ( .B(A[25]), .A(n42), .Z(n1134) );
  XNOR U1228 ( .A(n1142), .B(n1308), .Z(n1135) );
  XNOR U1229 ( .A(n1141), .B(n1139), .Z(n1308) );
  AND U1230 ( .A(n1309), .B(n1310), .Z(n1139) );
  NANDN U1231 ( .A(n1311), .B(n1312), .Z(n1310) );
  OR U1232 ( .A(n1313), .B(n1314), .Z(n1312) );
  NAND U1233 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1234 ( .B(A[24]), .A(n41), .Z(n1141) );
  XNOR U1235 ( .A(n1149), .B(n1315), .Z(n1142) );
  XNOR U1236 ( .A(n1148), .B(n1146), .Z(n1315) );
  AND U1237 ( .A(n1316), .B(n1317), .Z(n1146) );
  NANDN U1238 ( .A(n1318), .B(n1319), .Z(n1317) );
  NANDN U1239 ( .A(n1320), .B(n1321), .Z(n1319) );
  NANDN U1240 ( .A(n1321), .B(n1320), .Z(n1316) );
  AND U1241 ( .A(A[23]), .B(B[2]), .Z(n1148) );
  XNOR U1242 ( .A(n1156), .B(n1322), .Z(n1149) );
  XNOR U1243 ( .A(n1155), .B(n1153), .Z(n1322) );
  AND U1244 ( .A(n1323), .B(n1324), .Z(n1153) );
  NANDN U1245 ( .A(n1325), .B(n1326), .Z(n1324) );
  OR U1246 ( .A(n1327), .B(n1328), .Z(n1326) );
  NAND U1247 ( .A(n1328), .B(n1327), .Z(n1323) );
  AND U1248 ( .A(A[22]), .B(B[3]), .Z(n1155) );
  XNOR U1249 ( .A(n1163), .B(n1329), .Z(n1156) );
  XNOR U1250 ( .A(n1162), .B(n1160), .Z(n1329) );
  AND U1251 ( .A(n1330), .B(n1331), .Z(n1160) );
  NANDN U1252 ( .A(n1332), .B(n1333), .Z(n1331) );
  NANDN U1253 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1254 ( .A(n1335), .B(n1334), .Z(n1330) );
  AND U1255 ( .A(A[21]), .B(B[4]), .Z(n1162) );
  XNOR U1256 ( .A(n1170), .B(n1336), .Z(n1163) );
  XNOR U1257 ( .A(n1169), .B(n1167), .Z(n1336) );
  AND U1258 ( .A(n1337), .B(n1338), .Z(n1167) );
  NANDN U1259 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1260 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1261 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U1262 ( .A(A[20]), .B(B[5]), .Z(n1169) );
  XNOR U1263 ( .A(n1177), .B(n1343), .Z(n1170) );
  XNOR U1264 ( .A(n1176), .B(n1174), .Z(n1343) );
  AND U1265 ( .A(n1344), .B(n1345), .Z(n1174) );
  NANDN U1266 ( .A(n1346), .B(n1347), .Z(n1345) );
  NANDN U1267 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1268 ( .A(n1349), .B(n1348), .Z(n1344) );
  AND U1269 ( .A(A[19]), .B(B[6]), .Z(n1176) );
  XNOR U1270 ( .A(n1184), .B(n1350), .Z(n1177) );
  XNOR U1271 ( .A(n1183), .B(n1181), .Z(n1350) );
  AND U1272 ( .A(n1351), .B(n1352), .Z(n1181) );
  NANDN U1273 ( .A(n1353), .B(n1354), .Z(n1352) );
  OR U1274 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1275 ( .A(n1356), .B(n1355), .Z(n1351) );
  AND U1276 ( .A(A[18]), .B(B[7]), .Z(n1183) );
  XNOR U1277 ( .A(n1191), .B(n1357), .Z(n1184) );
  XNOR U1278 ( .A(n1190), .B(n1188), .Z(n1357) );
  AND U1279 ( .A(n1358), .B(n1359), .Z(n1188) );
  NANDN U1280 ( .A(n1360), .B(n1361), .Z(n1359) );
  NANDN U1281 ( .A(n1362), .B(n1363), .Z(n1361) );
  NANDN U1282 ( .A(n1363), .B(n1362), .Z(n1358) );
  AND U1283 ( .A(A[17]), .B(B[8]), .Z(n1190) );
  XNOR U1284 ( .A(n1198), .B(n1364), .Z(n1191) );
  XNOR U1285 ( .A(n1197), .B(n1195), .Z(n1364) );
  AND U1286 ( .A(n1365), .B(n1366), .Z(n1195) );
  NANDN U1287 ( .A(n1367), .B(n1368), .Z(n1366) );
  OR U1288 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1289 ( .A(n1370), .B(n1369), .Z(n1365) );
  AND U1290 ( .A(A[16]), .B(B[9]), .Z(n1197) );
  XNOR U1291 ( .A(n1205), .B(n1371), .Z(n1198) );
  XNOR U1292 ( .A(n1204), .B(n1202), .Z(n1371) );
  AND U1293 ( .A(n1372), .B(n1373), .Z(n1202) );
  NANDN U1294 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1295 ( .A(n1376), .B(n1377), .Z(n1375) );
  NANDN U1296 ( .A(n1377), .B(n1376), .Z(n1372) );
  AND U1297 ( .A(A[15]), .B(B[10]), .Z(n1204) );
  XNOR U1298 ( .A(n1212), .B(n1378), .Z(n1205) );
  XNOR U1299 ( .A(n1211), .B(n1209), .Z(n1378) );
  AND U1300 ( .A(n1379), .B(n1380), .Z(n1209) );
  NANDN U1301 ( .A(n1381), .B(n1382), .Z(n1380) );
  OR U1302 ( .A(n1383), .B(n1384), .Z(n1382) );
  NAND U1303 ( .A(n1384), .B(n1383), .Z(n1379) );
  AND U1304 ( .A(A[14]), .B(B[11]), .Z(n1211) );
  XNOR U1305 ( .A(n1219), .B(n1385), .Z(n1212) );
  XNOR U1306 ( .A(n1218), .B(n1216), .Z(n1385) );
  AND U1307 ( .A(n1386), .B(n1387), .Z(n1216) );
  NANDN U1308 ( .A(n1388), .B(n1389), .Z(n1387) );
  NANDN U1309 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U1310 ( .A(n1391), .B(n1390), .Z(n1386) );
  AND U1311 ( .A(A[13]), .B(B[12]), .Z(n1218) );
  XNOR U1312 ( .A(n1226), .B(n1392), .Z(n1219) );
  XNOR U1313 ( .A(n1225), .B(n1223), .Z(n1392) );
  AND U1314 ( .A(n1393), .B(n1394), .Z(n1223) );
  NANDN U1315 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1316 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U1317 ( .A(n1398), .B(n1397), .Z(n1393) );
  AND U1318 ( .A(A[12]), .B(B[13]), .Z(n1225) );
  XNOR U1319 ( .A(n1233), .B(n1399), .Z(n1226) );
  XNOR U1320 ( .A(n1232), .B(n1230), .Z(n1399) );
  AND U1321 ( .A(n1400), .B(n1401), .Z(n1230) );
  NANDN U1322 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1323 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1324 ( .A(n1405), .B(n1404), .Z(n1400) );
  AND U1325 ( .A(A[11]), .B(B[14]), .Z(n1232) );
  XNOR U1326 ( .A(n1240), .B(n1406), .Z(n1233) );
  XNOR U1327 ( .A(n1239), .B(n1237), .Z(n1406) );
  AND U1328 ( .A(n1407), .B(n1408), .Z(n1237) );
  NANDN U1329 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U1330 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1331 ( .A(n1412), .B(n1411), .Z(n1407) );
  AND U1332 ( .A(A[10]), .B(B[15]), .Z(n1239) );
  XNOR U1333 ( .A(n1247), .B(n1413), .Z(n1240) );
  XNOR U1334 ( .A(n1246), .B(n1244), .Z(n1413) );
  AND U1335 ( .A(n1414), .B(n1415), .Z(n1244) );
  NANDN U1336 ( .A(n1416), .B(n1417), .Z(n1415) );
  NANDN U1337 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1338 ( .A(n1419), .B(n1418), .Z(n1414) );
  AND U1339 ( .A(A[9]), .B(B[16]), .Z(n1246) );
  XNOR U1340 ( .A(n1254), .B(n1420), .Z(n1247) );
  XNOR U1341 ( .A(n1253), .B(n1251), .Z(n1420) );
  AND U1342 ( .A(n1421), .B(n1422), .Z(n1251) );
  NANDN U1343 ( .A(n1423), .B(n1424), .Z(n1422) );
  OR U1344 ( .A(n1425), .B(n1426), .Z(n1424) );
  NAND U1345 ( .A(n1426), .B(n1425), .Z(n1421) );
  AND U1346 ( .A(A[8]), .B(B[17]), .Z(n1253) );
  XNOR U1347 ( .A(n1261), .B(n1427), .Z(n1254) );
  XNOR U1348 ( .A(n1260), .B(n1258), .Z(n1427) );
  AND U1349 ( .A(n1428), .B(n1429), .Z(n1258) );
  NANDN U1350 ( .A(n1430), .B(n1431), .Z(n1429) );
  NANDN U1351 ( .A(n1432), .B(n1433), .Z(n1431) );
  NANDN U1352 ( .A(n1433), .B(n1432), .Z(n1428) );
  AND U1353 ( .A(A[7]), .B(B[18]), .Z(n1260) );
  XNOR U1354 ( .A(n1268), .B(n1434), .Z(n1261) );
  XNOR U1355 ( .A(n1267), .B(n1265), .Z(n1434) );
  AND U1356 ( .A(n1435), .B(n1436), .Z(n1265) );
  NANDN U1357 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U1358 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1359 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U1360 ( .A(A[6]), .B(B[19]), .Z(n1267) );
  XNOR U1361 ( .A(n1275), .B(n1441), .Z(n1268) );
  XNOR U1362 ( .A(n1274), .B(n1272), .Z(n1441) );
  AND U1363 ( .A(n1442), .B(n1443), .Z(n1272) );
  NANDN U1364 ( .A(n1444), .B(n1445), .Z(n1443) );
  NANDN U1365 ( .A(n1446), .B(n1447), .Z(n1445) );
  NANDN U1366 ( .A(n1447), .B(n1446), .Z(n1442) );
  AND U1367 ( .A(A[5]), .B(B[20]), .Z(n1274) );
  XNOR U1368 ( .A(n1282), .B(n1448), .Z(n1275) );
  XNOR U1369 ( .A(n1281), .B(n1279), .Z(n1448) );
  AND U1370 ( .A(n1449), .B(n1450), .Z(n1279) );
  NANDN U1371 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U1372 ( .A(n1453), .B(n1454), .Z(n1452) );
  NAND U1373 ( .A(n1454), .B(n1453), .Z(n1449) );
  AND U1374 ( .A(A[4]), .B(B[21]), .Z(n1281) );
  XNOR U1375 ( .A(n1289), .B(n1455), .Z(n1282) );
  XNOR U1376 ( .A(n1288), .B(n1286), .Z(n1455) );
  AND U1377 ( .A(n1456), .B(n1457), .Z(n1286) );
  NANDN U1378 ( .A(n1458), .B(n1459), .Z(n1457) );
  NAND U1379 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1380 ( .A(n1461), .B(n18), .Z(n1456) );
  AND U1381 ( .A(A[3]), .B(B[22]), .Z(n1288) );
  XOR U1382 ( .A(n1295), .B(n1462), .Z(n1289) );
  XNOR U1383 ( .A(n1293), .B(n1296), .Z(n1462) );
  NAND U1384 ( .A(A[2]), .B(B[23]), .Z(n1296) );
  NANDN U1385 ( .A(n1463), .B(n1464), .Z(n1293) );
  AND U1386 ( .A(A[0]), .B(B[24]), .Z(n1464) );
  XNOR U1387 ( .A(n1298), .B(n1465), .Z(n1295) );
  NAND U1388 ( .A(A[0]), .B(B[25]), .Z(n1465) );
  NAND U1389 ( .A(B[24]), .B(A[1]), .Z(n1298) );
  XOR U1390 ( .A(n1307), .B(n1466), .Z(PRODUCT[24]) );
  XNOR U1391 ( .A(n1306), .B(n1305), .Z(n1466) );
  NAND U1392 ( .A(n1467), .B(n1468), .Z(n1305) );
  NANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1394 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1395 ( .A(n1472), .B(n1471), .Z(n1467) );
  ANDN U1396 ( .B(A[24]), .A(n42), .Z(n1306) );
  XNOR U1397 ( .A(n1314), .B(n1473), .Z(n1307) );
  XNOR U1398 ( .A(n1313), .B(n1311), .Z(n1473) );
  AND U1399 ( .A(n1474), .B(n1475), .Z(n1311) );
  NANDN U1400 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1401 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1402 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1403 ( .B(A[23]), .A(n41), .Z(n1313) );
  XNOR U1404 ( .A(n1321), .B(n1480), .Z(n1314) );
  XNOR U1405 ( .A(n1320), .B(n1318), .Z(n1480) );
  AND U1406 ( .A(n1481), .B(n1482), .Z(n1318) );
  NANDN U1407 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1408 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1409 ( .A(n1486), .B(n1485), .Z(n1481) );
  AND U1410 ( .A(A[22]), .B(B[2]), .Z(n1320) );
  XNOR U1411 ( .A(n1328), .B(n1487), .Z(n1321) );
  XNOR U1412 ( .A(n1327), .B(n1325), .Z(n1487) );
  AND U1413 ( .A(n1488), .B(n1489), .Z(n1325) );
  NANDN U1414 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1415 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1416 ( .A(n1493), .B(n1492), .Z(n1488) );
  AND U1417 ( .A(A[21]), .B(B[3]), .Z(n1327) );
  XNOR U1418 ( .A(n1335), .B(n1494), .Z(n1328) );
  XNOR U1419 ( .A(n1334), .B(n1332), .Z(n1494) );
  AND U1420 ( .A(n1495), .B(n1496), .Z(n1332) );
  NANDN U1421 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1422 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1423 ( .A(n1500), .B(n1499), .Z(n1495) );
  AND U1424 ( .A(A[20]), .B(B[4]), .Z(n1334) );
  XNOR U1425 ( .A(n1342), .B(n1501), .Z(n1335) );
  XNOR U1426 ( .A(n1341), .B(n1339), .Z(n1501) );
  AND U1427 ( .A(n1502), .B(n1503), .Z(n1339) );
  NANDN U1428 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1429 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1430 ( .A(n1507), .B(n1506), .Z(n1502) );
  AND U1431 ( .A(A[19]), .B(B[5]), .Z(n1341) );
  XNOR U1432 ( .A(n1349), .B(n1508), .Z(n1342) );
  XNOR U1433 ( .A(n1348), .B(n1346), .Z(n1508) );
  AND U1434 ( .A(n1509), .B(n1510), .Z(n1346) );
  NANDN U1435 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1436 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1437 ( .A(n1514), .B(n1513), .Z(n1509) );
  AND U1438 ( .A(A[18]), .B(B[6]), .Z(n1348) );
  XNOR U1439 ( .A(n1356), .B(n1515), .Z(n1349) );
  XNOR U1440 ( .A(n1355), .B(n1353), .Z(n1515) );
  AND U1441 ( .A(n1516), .B(n1517), .Z(n1353) );
  NANDN U1442 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1443 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1444 ( .A(n1521), .B(n1520), .Z(n1516) );
  AND U1445 ( .A(A[17]), .B(B[7]), .Z(n1355) );
  XNOR U1446 ( .A(n1363), .B(n1522), .Z(n1356) );
  XNOR U1447 ( .A(n1362), .B(n1360), .Z(n1522) );
  AND U1448 ( .A(n1523), .B(n1524), .Z(n1360) );
  NANDN U1449 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1450 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1451 ( .A(n1528), .B(n1527), .Z(n1523) );
  AND U1452 ( .A(A[16]), .B(B[8]), .Z(n1362) );
  XNOR U1453 ( .A(n1370), .B(n1529), .Z(n1363) );
  XNOR U1454 ( .A(n1369), .B(n1367), .Z(n1529) );
  AND U1455 ( .A(n1530), .B(n1531), .Z(n1367) );
  NANDN U1456 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1457 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1458 ( .A(n1535), .B(n1534), .Z(n1530) );
  AND U1459 ( .A(A[15]), .B(B[9]), .Z(n1369) );
  XNOR U1460 ( .A(n1377), .B(n1536), .Z(n1370) );
  XNOR U1461 ( .A(n1376), .B(n1374), .Z(n1536) );
  AND U1462 ( .A(n1537), .B(n1538), .Z(n1374) );
  NANDN U1463 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1464 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1465 ( .A(n1542), .B(n1541), .Z(n1537) );
  AND U1466 ( .A(A[14]), .B(B[10]), .Z(n1376) );
  XNOR U1467 ( .A(n1384), .B(n1543), .Z(n1377) );
  XNOR U1468 ( .A(n1383), .B(n1381), .Z(n1543) );
  AND U1469 ( .A(n1544), .B(n1545), .Z(n1381) );
  NANDN U1470 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1471 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1472 ( .A(n1549), .B(n1548), .Z(n1544) );
  AND U1473 ( .A(A[13]), .B(B[11]), .Z(n1383) );
  XNOR U1474 ( .A(n1391), .B(n1550), .Z(n1384) );
  XNOR U1475 ( .A(n1390), .B(n1388), .Z(n1550) );
  AND U1476 ( .A(n1551), .B(n1552), .Z(n1388) );
  NANDN U1477 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1478 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1479 ( .A(n1556), .B(n1555), .Z(n1551) );
  AND U1480 ( .A(A[12]), .B(B[12]), .Z(n1390) );
  XNOR U1481 ( .A(n1398), .B(n1557), .Z(n1391) );
  XNOR U1482 ( .A(n1397), .B(n1395), .Z(n1557) );
  AND U1483 ( .A(n1558), .B(n1559), .Z(n1395) );
  NANDN U1484 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1485 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1486 ( .A(n1563), .B(n1562), .Z(n1558) );
  AND U1487 ( .A(A[11]), .B(B[13]), .Z(n1397) );
  XNOR U1488 ( .A(n1405), .B(n1564), .Z(n1398) );
  XNOR U1489 ( .A(n1404), .B(n1402), .Z(n1564) );
  AND U1490 ( .A(n1565), .B(n1566), .Z(n1402) );
  NANDN U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1492 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1493 ( .A(n1570), .B(n1569), .Z(n1565) );
  AND U1494 ( .A(A[10]), .B(B[14]), .Z(n1404) );
  XNOR U1495 ( .A(n1412), .B(n1571), .Z(n1405) );
  XNOR U1496 ( .A(n1411), .B(n1409), .Z(n1571) );
  AND U1497 ( .A(n1572), .B(n1573), .Z(n1409) );
  NANDN U1498 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1499 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1500 ( .A(n1577), .B(n1576), .Z(n1572) );
  AND U1501 ( .A(A[9]), .B(B[15]), .Z(n1411) );
  XNOR U1502 ( .A(n1419), .B(n1578), .Z(n1412) );
  XNOR U1503 ( .A(n1418), .B(n1416), .Z(n1578) );
  AND U1504 ( .A(n1579), .B(n1580), .Z(n1416) );
  NANDN U1505 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1506 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1507 ( .A(n1584), .B(n1583), .Z(n1579) );
  AND U1508 ( .A(A[8]), .B(B[16]), .Z(n1418) );
  XNOR U1509 ( .A(n1426), .B(n1585), .Z(n1419) );
  XNOR U1510 ( .A(n1425), .B(n1423), .Z(n1585) );
  AND U1511 ( .A(n1586), .B(n1587), .Z(n1423) );
  NANDN U1512 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1513 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1514 ( .A(n1591), .B(n1590), .Z(n1586) );
  AND U1515 ( .A(A[7]), .B(B[17]), .Z(n1425) );
  XNOR U1516 ( .A(n1433), .B(n1592), .Z(n1426) );
  XNOR U1517 ( .A(n1432), .B(n1430), .Z(n1592) );
  AND U1518 ( .A(n1593), .B(n1594), .Z(n1430) );
  NANDN U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1520 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1521 ( .A(n1598), .B(n1597), .Z(n1593) );
  AND U1522 ( .A(A[6]), .B(B[18]), .Z(n1432) );
  XNOR U1523 ( .A(n1440), .B(n1599), .Z(n1433) );
  XNOR U1524 ( .A(n1439), .B(n1437), .Z(n1599) );
  AND U1525 ( .A(n1600), .B(n1601), .Z(n1437) );
  NANDN U1526 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1527 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1528 ( .A(n1605), .B(n1604), .Z(n1600) );
  AND U1529 ( .A(A[5]), .B(B[19]), .Z(n1439) );
  XNOR U1530 ( .A(n1447), .B(n1606), .Z(n1440) );
  XNOR U1531 ( .A(n1446), .B(n1444), .Z(n1606) );
  AND U1532 ( .A(n1607), .B(n1608), .Z(n1444) );
  NANDN U1533 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1534 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1535 ( .A(n1612), .B(n1611), .Z(n1607) );
  AND U1536 ( .A(A[4]), .B(B[20]), .Z(n1446) );
  XNOR U1537 ( .A(n1454), .B(n1613), .Z(n1447) );
  XNOR U1538 ( .A(n1453), .B(n1451), .Z(n1613) );
  AND U1539 ( .A(n1614), .B(n1615), .Z(n1451) );
  NANDN U1540 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1541 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1542 ( .A(n1619), .B(n19), .Z(n1614) );
  AND U1543 ( .A(A[3]), .B(B[21]), .Z(n1453) );
  XOR U1544 ( .A(n1460), .B(n1620), .Z(n1454) );
  XNOR U1545 ( .A(n1458), .B(n1461), .Z(n1620) );
  NAND U1546 ( .A(A[2]), .B(B[22]), .Z(n1461) );
  NANDN U1547 ( .A(n1621), .B(n1622), .Z(n1458) );
  AND U1548 ( .A(A[0]), .B(B[23]), .Z(n1622) );
  XNOR U1549 ( .A(n1463), .B(n1623), .Z(n1460) );
  NAND U1550 ( .A(A[0]), .B(B[24]), .Z(n1623) );
  NAND U1551 ( .A(B[23]), .B(A[1]), .Z(n1463) );
  XOR U1552 ( .A(n1472), .B(n1624), .Z(PRODUCT[23]) );
  XNOR U1553 ( .A(n1471), .B(n1469), .Z(n1624) );
  AND U1554 ( .A(n1625), .B(n1626), .Z(n1469) );
  NAND U1555 ( .A(n1627), .B(n1628), .Z(n1626) );
  NANDN U1556 ( .A(n1629), .B(n1630), .Z(n1627) );
  NANDN U1557 ( .A(n1630), .B(n1629), .Z(n1625) );
  ANDN U1558 ( .B(A[23]), .A(n42), .Z(n1471) );
  XNOR U1559 ( .A(n1479), .B(n1631), .Z(n1472) );
  XNOR U1560 ( .A(n1478), .B(n1476), .Z(n1631) );
  AND U1561 ( .A(n1632), .B(n1633), .Z(n1476) );
  NANDN U1562 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1563 ( .A(n1636), .B(n1637), .Z(n1635) );
  NAND U1564 ( .A(n1637), .B(n1636), .Z(n1632) );
  ANDN U1565 ( .B(A[22]), .A(n41), .Z(n1478) );
  XNOR U1566 ( .A(n1486), .B(n1638), .Z(n1479) );
  XNOR U1567 ( .A(n1485), .B(n1483), .Z(n1638) );
  AND U1568 ( .A(n1639), .B(n1640), .Z(n1483) );
  NANDN U1569 ( .A(n1641), .B(n1642), .Z(n1640) );
  NANDN U1570 ( .A(n1643), .B(n1644), .Z(n1642) );
  NANDN U1571 ( .A(n1644), .B(n1643), .Z(n1639) );
  AND U1572 ( .A(A[21]), .B(B[2]), .Z(n1485) );
  XNOR U1573 ( .A(n1493), .B(n1645), .Z(n1486) );
  XNOR U1574 ( .A(n1492), .B(n1490), .Z(n1645) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1490) );
  NANDN U1576 ( .A(n1648), .B(n1649), .Z(n1647) );
  OR U1577 ( .A(n1650), .B(n1651), .Z(n1649) );
  NAND U1578 ( .A(n1651), .B(n1650), .Z(n1646) );
  AND U1579 ( .A(A[20]), .B(B[3]), .Z(n1492) );
  XNOR U1580 ( .A(n1500), .B(n1652), .Z(n1493) );
  XNOR U1581 ( .A(n1499), .B(n1497), .Z(n1652) );
  AND U1582 ( .A(n1653), .B(n1654), .Z(n1497) );
  NANDN U1583 ( .A(n1655), .B(n1656), .Z(n1654) );
  NANDN U1584 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U1585 ( .A(n1658), .B(n1657), .Z(n1653) );
  AND U1586 ( .A(A[19]), .B(B[4]), .Z(n1499) );
  XNOR U1587 ( .A(n1507), .B(n1659), .Z(n1500) );
  XNOR U1588 ( .A(n1506), .B(n1504), .Z(n1659) );
  AND U1589 ( .A(n1660), .B(n1661), .Z(n1504) );
  NANDN U1590 ( .A(n1662), .B(n1663), .Z(n1661) );
  OR U1591 ( .A(n1664), .B(n1665), .Z(n1663) );
  NAND U1592 ( .A(n1665), .B(n1664), .Z(n1660) );
  AND U1593 ( .A(A[18]), .B(B[5]), .Z(n1506) );
  XNOR U1594 ( .A(n1514), .B(n1666), .Z(n1507) );
  XNOR U1595 ( .A(n1513), .B(n1511), .Z(n1666) );
  AND U1596 ( .A(n1667), .B(n1668), .Z(n1511) );
  NANDN U1597 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1598 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U1599 ( .A(n1672), .B(n1671), .Z(n1667) );
  AND U1600 ( .A(A[17]), .B(B[6]), .Z(n1513) );
  XNOR U1601 ( .A(n1521), .B(n1673), .Z(n1514) );
  XNOR U1602 ( .A(n1520), .B(n1518), .Z(n1673) );
  AND U1603 ( .A(n1674), .B(n1675), .Z(n1518) );
  NANDN U1604 ( .A(n1676), .B(n1677), .Z(n1675) );
  OR U1605 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1606 ( .A(n1679), .B(n1678), .Z(n1674) );
  AND U1607 ( .A(A[16]), .B(B[7]), .Z(n1520) );
  XNOR U1608 ( .A(n1528), .B(n1680), .Z(n1521) );
  XNOR U1609 ( .A(n1527), .B(n1525), .Z(n1680) );
  AND U1610 ( .A(n1681), .B(n1682), .Z(n1525) );
  NANDN U1611 ( .A(n1683), .B(n1684), .Z(n1682) );
  NANDN U1612 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1613 ( .A(n1686), .B(n1685), .Z(n1681) );
  AND U1614 ( .A(A[15]), .B(B[8]), .Z(n1527) );
  XNOR U1615 ( .A(n1535), .B(n1687), .Z(n1528) );
  XNOR U1616 ( .A(n1534), .B(n1532), .Z(n1687) );
  AND U1617 ( .A(n1688), .B(n1689), .Z(n1532) );
  NANDN U1618 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U1619 ( .A(n1692), .B(n1693), .Z(n1691) );
  NAND U1620 ( .A(n1693), .B(n1692), .Z(n1688) );
  AND U1621 ( .A(A[14]), .B(B[9]), .Z(n1534) );
  XNOR U1622 ( .A(n1542), .B(n1694), .Z(n1535) );
  XNOR U1623 ( .A(n1541), .B(n1539), .Z(n1694) );
  AND U1624 ( .A(n1695), .B(n1696), .Z(n1539) );
  NANDN U1625 ( .A(n1697), .B(n1698), .Z(n1696) );
  NANDN U1626 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U1627 ( .A(n1700), .B(n1699), .Z(n1695) );
  AND U1628 ( .A(A[13]), .B(B[10]), .Z(n1541) );
  XNOR U1629 ( .A(n1549), .B(n1701), .Z(n1542) );
  XNOR U1630 ( .A(n1548), .B(n1546), .Z(n1701) );
  AND U1631 ( .A(n1702), .B(n1703), .Z(n1546) );
  NANDN U1632 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1633 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1634 ( .A(n1707), .B(n1706), .Z(n1702) );
  AND U1635 ( .A(A[12]), .B(B[11]), .Z(n1548) );
  XNOR U1636 ( .A(n1556), .B(n1708), .Z(n1549) );
  XNOR U1637 ( .A(n1555), .B(n1553), .Z(n1708) );
  AND U1638 ( .A(n1709), .B(n1710), .Z(n1553) );
  NANDN U1639 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1640 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1641 ( .A(n1714), .B(n1713), .Z(n1709) );
  AND U1642 ( .A(A[11]), .B(B[12]), .Z(n1555) );
  XNOR U1643 ( .A(n1563), .B(n1715), .Z(n1556) );
  XNOR U1644 ( .A(n1562), .B(n1560), .Z(n1715) );
  AND U1645 ( .A(n1716), .B(n1717), .Z(n1560) );
  NANDN U1646 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1647 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1648 ( .A(n1721), .B(n1720), .Z(n1716) );
  AND U1649 ( .A(A[10]), .B(B[13]), .Z(n1562) );
  XNOR U1650 ( .A(n1570), .B(n1722), .Z(n1563) );
  XNOR U1651 ( .A(n1569), .B(n1567), .Z(n1722) );
  AND U1652 ( .A(n1723), .B(n1724), .Z(n1567) );
  NANDN U1653 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1654 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1655 ( .A(n1728), .B(n1727), .Z(n1723) );
  AND U1656 ( .A(A[9]), .B(B[14]), .Z(n1569) );
  XNOR U1657 ( .A(n1577), .B(n1729), .Z(n1570) );
  XNOR U1658 ( .A(n1576), .B(n1574), .Z(n1729) );
  AND U1659 ( .A(n1730), .B(n1731), .Z(n1574) );
  NANDN U1660 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1661 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1662 ( .A(n1735), .B(n1734), .Z(n1730) );
  AND U1663 ( .A(A[8]), .B(B[15]), .Z(n1576) );
  XNOR U1664 ( .A(n1584), .B(n1736), .Z(n1577) );
  XNOR U1665 ( .A(n1583), .B(n1581), .Z(n1736) );
  AND U1666 ( .A(n1737), .B(n1738), .Z(n1581) );
  NANDN U1667 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1668 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1669 ( .A(n1742), .B(n1741), .Z(n1737) );
  AND U1670 ( .A(A[7]), .B(B[16]), .Z(n1583) );
  XNOR U1671 ( .A(n1591), .B(n1743), .Z(n1584) );
  XNOR U1672 ( .A(n1590), .B(n1588), .Z(n1743) );
  AND U1673 ( .A(n1744), .B(n1745), .Z(n1588) );
  NANDN U1674 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1675 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1676 ( .A(n1749), .B(n1748), .Z(n1744) );
  AND U1677 ( .A(A[6]), .B(B[17]), .Z(n1590) );
  XNOR U1678 ( .A(n1598), .B(n1750), .Z(n1591) );
  XNOR U1679 ( .A(n1597), .B(n1595), .Z(n1750) );
  AND U1680 ( .A(n1751), .B(n1752), .Z(n1595) );
  NANDN U1681 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1682 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1683 ( .A(n1756), .B(n1755), .Z(n1751) );
  AND U1684 ( .A(A[5]), .B(B[18]), .Z(n1597) );
  XNOR U1685 ( .A(n1605), .B(n1757), .Z(n1598) );
  XNOR U1686 ( .A(n1604), .B(n1602), .Z(n1757) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1602) );
  NANDN U1688 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1689 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1690 ( .A(n1763), .B(n1762), .Z(n1758) );
  AND U1691 ( .A(A[4]), .B(B[19]), .Z(n1604) );
  XNOR U1692 ( .A(n1612), .B(n1764), .Z(n1605) );
  XNOR U1693 ( .A(n1611), .B(n1609), .Z(n1764) );
  AND U1694 ( .A(n1765), .B(n1766), .Z(n1609) );
  NANDN U1695 ( .A(n1767), .B(n1768), .Z(n1766) );
  NAND U1696 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1697 ( .A(n1770), .B(n20), .Z(n1765) );
  AND U1698 ( .A(A[3]), .B(B[20]), .Z(n1611) );
  XOR U1699 ( .A(n1618), .B(n1771), .Z(n1612) );
  XNOR U1700 ( .A(n1616), .B(n1619), .Z(n1771) );
  NAND U1701 ( .A(A[2]), .B(B[21]), .Z(n1619) );
  NANDN U1702 ( .A(n1772), .B(n1773), .Z(n1616) );
  AND U1703 ( .A(A[0]), .B(B[22]), .Z(n1773) );
  XNOR U1704 ( .A(n1621), .B(n1774), .Z(n1618) );
  NAND U1705 ( .A(A[0]), .B(B[23]), .Z(n1774) );
  NAND U1706 ( .A(B[22]), .B(A[1]), .Z(n1621) );
  XOR U1707 ( .A(n1630), .B(n1775), .Z(PRODUCT[22]) );
  XNOR U1708 ( .A(n1629), .B(n1628), .Z(n1775) );
  NAND U1709 ( .A(n1776), .B(n1777), .Z(n1628) );
  NANDN U1710 ( .A(n1778), .B(n1779), .Z(n1777) );
  OR U1711 ( .A(n1780), .B(n1781), .Z(n1779) );
  NAND U1712 ( .A(n1781), .B(n1780), .Z(n1776) );
  ANDN U1713 ( .B(A[22]), .A(n42), .Z(n1629) );
  XNOR U1714 ( .A(n1637), .B(n1782), .Z(n1630) );
  XNOR U1715 ( .A(n1636), .B(n1634), .Z(n1782) );
  AND U1716 ( .A(n1783), .B(n1784), .Z(n1634) );
  NANDN U1717 ( .A(n1785), .B(n1786), .Z(n1784) );
  NANDN U1718 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1719 ( .A(n1788), .B(n1787), .Z(n1783) );
  ANDN U1720 ( .B(A[21]), .A(n41), .Z(n1636) );
  XNOR U1721 ( .A(n1644), .B(n1789), .Z(n1637) );
  XNOR U1722 ( .A(n1643), .B(n1641), .Z(n1789) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1641) );
  NANDN U1724 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1725 ( .A(n1794), .B(n1795), .Z(n1793) );
  NAND U1726 ( .A(n1795), .B(n1794), .Z(n1790) );
  AND U1727 ( .A(A[20]), .B(B[2]), .Z(n1643) );
  XNOR U1728 ( .A(n1651), .B(n1796), .Z(n1644) );
  XNOR U1729 ( .A(n1650), .B(n1648), .Z(n1796) );
  AND U1730 ( .A(n1797), .B(n1798), .Z(n1648) );
  NANDN U1731 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1732 ( .A(n1801), .B(n1802), .Z(n1800) );
  NANDN U1733 ( .A(n1802), .B(n1801), .Z(n1797) );
  AND U1734 ( .A(A[19]), .B(B[3]), .Z(n1650) );
  XNOR U1735 ( .A(n1658), .B(n1803), .Z(n1651) );
  XNOR U1736 ( .A(n1657), .B(n1655), .Z(n1803) );
  AND U1737 ( .A(n1804), .B(n1805), .Z(n1655) );
  NANDN U1738 ( .A(n1806), .B(n1807), .Z(n1805) );
  OR U1739 ( .A(n1808), .B(n1809), .Z(n1807) );
  NAND U1740 ( .A(n1809), .B(n1808), .Z(n1804) );
  AND U1741 ( .A(A[18]), .B(B[4]), .Z(n1657) );
  XNOR U1742 ( .A(n1665), .B(n1810), .Z(n1658) );
  XNOR U1743 ( .A(n1664), .B(n1662), .Z(n1810) );
  AND U1744 ( .A(n1811), .B(n1812), .Z(n1662) );
  NANDN U1745 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1746 ( .A(n1815), .B(n1816), .Z(n1814) );
  NANDN U1747 ( .A(n1816), .B(n1815), .Z(n1811) );
  AND U1748 ( .A(A[17]), .B(B[5]), .Z(n1664) );
  XNOR U1749 ( .A(n1672), .B(n1817), .Z(n1665) );
  XNOR U1750 ( .A(n1671), .B(n1669), .Z(n1817) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1669) );
  NANDN U1752 ( .A(n1820), .B(n1821), .Z(n1819) );
  OR U1753 ( .A(n1822), .B(n1823), .Z(n1821) );
  NAND U1754 ( .A(n1823), .B(n1822), .Z(n1818) );
  AND U1755 ( .A(A[16]), .B(B[6]), .Z(n1671) );
  XNOR U1756 ( .A(n1679), .B(n1824), .Z(n1672) );
  XNOR U1757 ( .A(n1678), .B(n1676), .Z(n1824) );
  AND U1758 ( .A(n1825), .B(n1826), .Z(n1676) );
  NANDN U1759 ( .A(n1827), .B(n1828), .Z(n1826) );
  NANDN U1760 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1761 ( .A(n1830), .B(n1829), .Z(n1825) );
  AND U1762 ( .A(A[15]), .B(B[7]), .Z(n1678) );
  XNOR U1763 ( .A(n1686), .B(n1831), .Z(n1679) );
  XNOR U1764 ( .A(n1685), .B(n1683), .Z(n1831) );
  AND U1765 ( .A(n1832), .B(n1833), .Z(n1683) );
  NANDN U1766 ( .A(n1834), .B(n1835), .Z(n1833) );
  OR U1767 ( .A(n1836), .B(n1837), .Z(n1835) );
  NAND U1768 ( .A(n1837), .B(n1836), .Z(n1832) );
  AND U1769 ( .A(A[14]), .B(B[8]), .Z(n1685) );
  XNOR U1770 ( .A(n1693), .B(n1838), .Z(n1686) );
  XNOR U1771 ( .A(n1692), .B(n1690), .Z(n1838) );
  AND U1772 ( .A(n1839), .B(n1840), .Z(n1690) );
  NANDN U1773 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1774 ( .A(n1843), .B(n1844), .Z(n1842) );
  NANDN U1775 ( .A(n1844), .B(n1843), .Z(n1839) );
  AND U1776 ( .A(A[13]), .B(B[9]), .Z(n1692) );
  XNOR U1777 ( .A(n1700), .B(n1845), .Z(n1693) );
  XNOR U1778 ( .A(n1699), .B(n1697), .Z(n1845) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1697) );
  NANDN U1780 ( .A(n1848), .B(n1849), .Z(n1847) );
  OR U1781 ( .A(n1850), .B(n1851), .Z(n1849) );
  NAND U1782 ( .A(n1851), .B(n1850), .Z(n1846) );
  AND U1783 ( .A(A[12]), .B(B[10]), .Z(n1699) );
  XNOR U1784 ( .A(n1707), .B(n1852), .Z(n1700) );
  XNOR U1785 ( .A(n1706), .B(n1704), .Z(n1852) );
  AND U1786 ( .A(n1853), .B(n1854), .Z(n1704) );
  NANDN U1787 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1788 ( .A(n1857), .B(n1858), .Z(n1856) );
  NANDN U1789 ( .A(n1858), .B(n1857), .Z(n1853) );
  AND U1790 ( .A(A[11]), .B(B[11]), .Z(n1706) );
  XNOR U1791 ( .A(n1714), .B(n1859), .Z(n1707) );
  XNOR U1792 ( .A(n1713), .B(n1711), .Z(n1859) );
  AND U1793 ( .A(n1860), .B(n1861), .Z(n1711) );
  NANDN U1794 ( .A(n1862), .B(n1863), .Z(n1861) );
  OR U1795 ( .A(n1864), .B(n1865), .Z(n1863) );
  NAND U1796 ( .A(n1865), .B(n1864), .Z(n1860) );
  AND U1797 ( .A(A[10]), .B(B[12]), .Z(n1713) );
  XNOR U1798 ( .A(n1721), .B(n1866), .Z(n1714) );
  XNOR U1799 ( .A(n1720), .B(n1718), .Z(n1866) );
  AND U1800 ( .A(n1867), .B(n1868), .Z(n1718) );
  NANDN U1801 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1802 ( .A(n1871), .B(n1872), .Z(n1870) );
  NANDN U1803 ( .A(n1872), .B(n1871), .Z(n1867) );
  AND U1804 ( .A(A[9]), .B(B[13]), .Z(n1720) );
  XNOR U1805 ( .A(n1728), .B(n1873), .Z(n1721) );
  XNOR U1806 ( .A(n1727), .B(n1725), .Z(n1873) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1725) );
  NANDN U1808 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1809 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1810 ( .A(n1879), .B(n1878), .Z(n1874) );
  AND U1811 ( .A(A[8]), .B(B[14]), .Z(n1727) );
  XNOR U1812 ( .A(n1735), .B(n1880), .Z(n1728) );
  XNOR U1813 ( .A(n1734), .B(n1732), .Z(n1880) );
  AND U1814 ( .A(n1881), .B(n1882), .Z(n1732) );
  NANDN U1815 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1816 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1817 ( .A(n1886), .B(n1885), .Z(n1881) );
  AND U1818 ( .A(A[7]), .B(B[15]), .Z(n1734) );
  XNOR U1819 ( .A(n1742), .B(n1887), .Z(n1735) );
  XNOR U1820 ( .A(n1741), .B(n1739), .Z(n1887) );
  AND U1821 ( .A(n1888), .B(n1889), .Z(n1739) );
  NANDN U1822 ( .A(n1890), .B(n1891), .Z(n1889) );
  OR U1823 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND U1824 ( .A(n1893), .B(n1892), .Z(n1888) );
  AND U1825 ( .A(A[6]), .B(B[16]), .Z(n1741) );
  XNOR U1826 ( .A(n1749), .B(n1894), .Z(n1742) );
  XNOR U1827 ( .A(n1748), .B(n1746), .Z(n1894) );
  AND U1828 ( .A(n1895), .B(n1896), .Z(n1746) );
  NANDN U1829 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1830 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U1831 ( .A(n1900), .B(n1899), .Z(n1895) );
  AND U1832 ( .A(A[5]), .B(B[17]), .Z(n1748) );
  XNOR U1833 ( .A(n1756), .B(n1901), .Z(n1749) );
  XNOR U1834 ( .A(n1755), .B(n1753), .Z(n1901) );
  AND U1835 ( .A(n1902), .B(n1903), .Z(n1753) );
  NANDN U1836 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U1837 ( .A(n1906), .B(n1907), .Z(n1905) );
  NAND U1838 ( .A(n1907), .B(n1906), .Z(n1902) );
  AND U1839 ( .A(A[4]), .B(B[18]), .Z(n1755) );
  XNOR U1840 ( .A(n1763), .B(n1908), .Z(n1756) );
  XNOR U1841 ( .A(n1762), .B(n1760), .Z(n1908) );
  AND U1842 ( .A(n1909), .B(n1910), .Z(n1760) );
  NANDN U1843 ( .A(n1911), .B(n1912), .Z(n1910) );
  NAND U1844 ( .A(n1913), .B(n1914), .Z(n1912) );
  NANDN U1845 ( .A(n1914), .B(n21), .Z(n1909) );
  AND U1846 ( .A(A[3]), .B(B[19]), .Z(n1762) );
  XOR U1847 ( .A(n1769), .B(n1915), .Z(n1763) );
  XNOR U1848 ( .A(n1767), .B(n1770), .Z(n1915) );
  NAND U1849 ( .A(A[2]), .B(B[20]), .Z(n1770) );
  NANDN U1850 ( .A(n1916), .B(n1917), .Z(n1767) );
  AND U1851 ( .A(A[0]), .B(B[21]), .Z(n1917) );
  XNOR U1852 ( .A(n1772), .B(n1918), .Z(n1769) );
  NAND U1853 ( .A(A[0]), .B(B[22]), .Z(n1918) );
  NAND U1854 ( .A(B[21]), .B(A[1]), .Z(n1772) );
  XOR U1855 ( .A(n1919), .B(n1920), .Z(PRODUCT[3]) );
  XNOR U1856 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1857 ( .A(n1781), .B(n1923), .Z(PRODUCT[21]) );
  XNOR U1858 ( .A(n1780), .B(n1778), .Z(n1923) );
  AND U1859 ( .A(n1924), .B(n1925), .Z(n1778) );
  NAND U1860 ( .A(n1926), .B(n1927), .Z(n1925) );
  NANDN U1861 ( .A(n1928), .B(n1929), .Z(n1926) );
  NANDN U1862 ( .A(n1929), .B(n1928), .Z(n1924) );
  ANDN U1863 ( .B(A[21]), .A(n42), .Z(n1780) );
  XNOR U1864 ( .A(n1788), .B(n1930), .Z(n1781) );
  XNOR U1865 ( .A(n1787), .B(n1785), .Z(n1930) );
  AND U1866 ( .A(n1931), .B(n1932), .Z(n1785) );
  NANDN U1867 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U1868 ( .A(n1935), .B(n1936), .Z(n1934) );
  NAND U1869 ( .A(n1936), .B(n1935), .Z(n1931) );
  ANDN U1870 ( .B(A[20]), .A(n41), .Z(n1787) );
  XNOR U1871 ( .A(n1795), .B(n1937), .Z(n1788) );
  XNOR U1872 ( .A(n1794), .B(n1792), .Z(n1937) );
  AND U1873 ( .A(n1938), .B(n1939), .Z(n1792) );
  NANDN U1874 ( .A(n1940), .B(n1941), .Z(n1939) );
  NANDN U1875 ( .A(n1942), .B(n1943), .Z(n1941) );
  NANDN U1876 ( .A(n1943), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(A[19]), .B(B[2]), .Z(n1794) );
  XNOR U1878 ( .A(n1802), .B(n1944), .Z(n1795) );
  XNOR U1879 ( .A(n1801), .B(n1799), .Z(n1944) );
  AND U1880 ( .A(n1945), .B(n1946), .Z(n1799) );
  NANDN U1881 ( .A(n1947), .B(n1948), .Z(n1946) );
  OR U1882 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND U1883 ( .A(n1950), .B(n1949), .Z(n1945) );
  AND U1884 ( .A(A[18]), .B(B[3]), .Z(n1801) );
  XNOR U1885 ( .A(n1809), .B(n1951), .Z(n1802) );
  XNOR U1886 ( .A(n1808), .B(n1806), .Z(n1951) );
  AND U1887 ( .A(n1952), .B(n1953), .Z(n1806) );
  NANDN U1888 ( .A(n1954), .B(n1955), .Z(n1953) );
  NANDN U1889 ( .A(n1956), .B(n1957), .Z(n1955) );
  NANDN U1890 ( .A(n1957), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(A[17]), .B(B[4]), .Z(n1808) );
  XNOR U1892 ( .A(n1816), .B(n1958), .Z(n1809) );
  XNOR U1893 ( .A(n1815), .B(n1813), .Z(n1958) );
  AND U1894 ( .A(n1959), .B(n1960), .Z(n1813) );
  NANDN U1895 ( .A(n1961), .B(n1962), .Z(n1960) );
  OR U1896 ( .A(n1963), .B(n1964), .Z(n1962) );
  NAND U1897 ( .A(n1964), .B(n1963), .Z(n1959) );
  AND U1898 ( .A(A[16]), .B(B[5]), .Z(n1815) );
  XNOR U1899 ( .A(n1823), .B(n1965), .Z(n1816) );
  XNOR U1900 ( .A(n1822), .B(n1820), .Z(n1965) );
  AND U1901 ( .A(n1966), .B(n1967), .Z(n1820) );
  NANDN U1902 ( .A(n1968), .B(n1969), .Z(n1967) );
  NANDN U1903 ( .A(n1970), .B(n1971), .Z(n1969) );
  NANDN U1904 ( .A(n1971), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(A[15]), .B(B[6]), .Z(n1822) );
  XNOR U1906 ( .A(n1830), .B(n1972), .Z(n1823) );
  XNOR U1907 ( .A(n1829), .B(n1827), .Z(n1972) );
  AND U1908 ( .A(n1973), .B(n1974), .Z(n1827) );
  NANDN U1909 ( .A(n1975), .B(n1976), .Z(n1974) );
  OR U1910 ( .A(n1977), .B(n1978), .Z(n1976) );
  NAND U1911 ( .A(n1978), .B(n1977), .Z(n1973) );
  AND U1912 ( .A(A[14]), .B(B[7]), .Z(n1829) );
  XNOR U1913 ( .A(n1837), .B(n1979), .Z(n1830) );
  XNOR U1914 ( .A(n1836), .B(n1834), .Z(n1979) );
  AND U1915 ( .A(n1980), .B(n1981), .Z(n1834) );
  NANDN U1916 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U1917 ( .A(n1984), .B(n1985), .Z(n1983) );
  NANDN U1918 ( .A(n1985), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(A[13]), .B(B[8]), .Z(n1836) );
  XNOR U1920 ( .A(n1844), .B(n1986), .Z(n1837) );
  XNOR U1921 ( .A(n1843), .B(n1841), .Z(n1986) );
  AND U1922 ( .A(n1987), .B(n1988), .Z(n1841) );
  NANDN U1923 ( .A(n1989), .B(n1990), .Z(n1988) );
  OR U1924 ( .A(n1991), .B(n1992), .Z(n1990) );
  NAND U1925 ( .A(n1992), .B(n1991), .Z(n1987) );
  AND U1926 ( .A(A[12]), .B(B[9]), .Z(n1843) );
  XNOR U1927 ( .A(n1851), .B(n1993), .Z(n1844) );
  XNOR U1928 ( .A(n1850), .B(n1848), .Z(n1993) );
  AND U1929 ( .A(n1994), .B(n1995), .Z(n1848) );
  NANDN U1930 ( .A(n1996), .B(n1997), .Z(n1995) );
  NANDN U1931 ( .A(n1998), .B(n1999), .Z(n1997) );
  NANDN U1932 ( .A(n1999), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(A[11]), .B(B[10]), .Z(n1850) );
  XNOR U1934 ( .A(n1858), .B(n2000), .Z(n1851) );
  XNOR U1935 ( .A(n1857), .B(n1855), .Z(n2000) );
  AND U1936 ( .A(n2001), .B(n2002), .Z(n1855) );
  NANDN U1937 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U1938 ( .A(n2005), .B(n2006), .Z(n2004) );
  NAND U1939 ( .A(n2006), .B(n2005), .Z(n2001) );
  AND U1940 ( .A(A[10]), .B(B[11]), .Z(n1857) );
  XNOR U1941 ( .A(n1865), .B(n2007), .Z(n1858) );
  XNOR U1942 ( .A(n1864), .B(n1862), .Z(n2007) );
  AND U1943 ( .A(n2008), .B(n2009), .Z(n1862) );
  NANDN U1944 ( .A(n2010), .B(n2011), .Z(n2009) );
  NANDN U1945 ( .A(n2012), .B(n2013), .Z(n2011) );
  NANDN U1946 ( .A(n2013), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(A[9]), .B(B[12]), .Z(n1864) );
  XNOR U1948 ( .A(n1872), .B(n2014), .Z(n1865) );
  XNOR U1949 ( .A(n1871), .B(n1869), .Z(n2014) );
  AND U1950 ( .A(n2015), .B(n2016), .Z(n1869) );
  NANDN U1951 ( .A(n2017), .B(n2018), .Z(n2016) );
  OR U1952 ( .A(n2019), .B(n2020), .Z(n2018) );
  NAND U1953 ( .A(n2020), .B(n2019), .Z(n2015) );
  AND U1954 ( .A(A[8]), .B(B[13]), .Z(n1871) );
  XNOR U1955 ( .A(n1879), .B(n2021), .Z(n1872) );
  XNOR U1956 ( .A(n1878), .B(n1876), .Z(n2021) );
  AND U1957 ( .A(n2022), .B(n2023), .Z(n1876) );
  NANDN U1958 ( .A(n2024), .B(n2025), .Z(n2023) );
  NANDN U1959 ( .A(n2026), .B(n2027), .Z(n2025) );
  NANDN U1960 ( .A(n2027), .B(n2026), .Z(n2022) );
  AND U1961 ( .A(A[7]), .B(B[14]), .Z(n1878) );
  XNOR U1962 ( .A(n1886), .B(n2028), .Z(n1879) );
  XNOR U1963 ( .A(n1885), .B(n1883), .Z(n2028) );
  AND U1964 ( .A(n2029), .B(n2030), .Z(n1883) );
  NANDN U1965 ( .A(n2031), .B(n2032), .Z(n2030) );
  OR U1966 ( .A(n2033), .B(n2034), .Z(n2032) );
  NAND U1967 ( .A(n2034), .B(n2033), .Z(n2029) );
  AND U1968 ( .A(A[6]), .B(B[15]), .Z(n1885) );
  XNOR U1969 ( .A(n1893), .B(n2035), .Z(n1886) );
  XNOR U1970 ( .A(n1892), .B(n1890), .Z(n2035) );
  AND U1971 ( .A(n2036), .B(n2037), .Z(n1890) );
  NANDN U1972 ( .A(n2038), .B(n2039), .Z(n2037) );
  NANDN U1973 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U1974 ( .A(n2041), .B(n2040), .Z(n2036) );
  AND U1975 ( .A(A[5]), .B(B[16]), .Z(n1892) );
  XNOR U1976 ( .A(n1900), .B(n2042), .Z(n1893) );
  XNOR U1977 ( .A(n1899), .B(n1897), .Z(n2042) );
  AND U1978 ( .A(n2043), .B(n2044), .Z(n1897) );
  NANDN U1979 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U1980 ( .A(n2047), .B(n2048), .Z(n2046) );
  NAND U1981 ( .A(n2048), .B(n2047), .Z(n2043) );
  AND U1982 ( .A(A[4]), .B(B[17]), .Z(n1899) );
  XNOR U1983 ( .A(n1907), .B(n2049), .Z(n1900) );
  XNOR U1984 ( .A(n1906), .B(n1904), .Z(n2049) );
  AND U1985 ( .A(n2050), .B(n2051), .Z(n1904) );
  NANDN U1986 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND U1987 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U1988 ( .A(n2055), .B(n22), .Z(n2050) );
  AND U1989 ( .A(A[3]), .B(B[18]), .Z(n1906) );
  XOR U1990 ( .A(n1913), .B(n2056), .Z(n1907) );
  XNOR U1991 ( .A(n1911), .B(n1914), .Z(n2056) );
  NAND U1992 ( .A(A[2]), .B(B[19]), .Z(n1914) );
  NANDN U1993 ( .A(n2057), .B(n2058), .Z(n1911) );
  AND U1994 ( .A(A[0]), .B(B[20]), .Z(n2058) );
  XNOR U1995 ( .A(n1916), .B(n2059), .Z(n1913) );
  NAND U1996 ( .A(A[0]), .B(B[21]), .Z(n2059) );
  NAND U1997 ( .A(B[20]), .B(A[1]), .Z(n1916) );
  XOR U1998 ( .A(n1929), .B(n2060), .Z(PRODUCT[20]) );
  XNOR U1999 ( .A(n1928), .B(n1927), .Z(n2060) );
  NAND U2000 ( .A(n2061), .B(n2062), .Z(n1927) );
  NANDN U2001 ( .A(n2063), .B(n2064), .Z(n2062) );
  OR U2002 ( .A(n2065), .B(n2066), .Z(n2064) );
  NAND U2003 ( .A(n2066), .B(n2065), .Z(n2061) );
  ANDN U2004 ( .B(A[20]), .A(n42), .Z(n1928) );
  XNOR U2005 ( .A(n1936), .B(n2067), .Z(n1929) );
  XNOR U2006 ( .A(n1935), .B(n1933), .Z(n2067) );
  AND U2007 ( .A(n2068), .B(n2069), .Z(n1933) );
  NANDN U2008 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2009 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2010 ( .A(n2073), .B(n2072), .Z(n2068) );
  ANDN U2011 ( .B(A[19]), .A(n41), .Z(n1935) );
  XNOR U2012 ( .A(n1943), .B(n2074), .Z(n1936) );
  XNOR U2013 ( .A(n1942), .B(n1940), .Z(n2074) );
  AND U2014 ( .A(n2075), .B(n2076), .Z(n1940) );
  NANDN U2015 ( .A(n2077), .B(n2078), .Z(n2076) );
  OR U2016 ( .A(n2079), .B(n2080), .Z(n2078) );
  NAND U2017 ( .A(n2080), .B(n2079), .Z(n2075) );
  AND U2018 ( .A(A[18]), .B(B[2]), .Z(n1942) );
  XNOR U2019 ( .A(n1950), .B(n2081), .Z(n1943) );
  XNOR U2020 ( .A(n1949), .B(n1947), .Z(n2081) );
  AND U2021 ( .A(n2082), .B(n2083), .Z(n1947) );
  NANDN U2022 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2023 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2024 ( .A(n2087), .B(n2086), .Z(n2082) );
  AND U2025 ( .A(A[17]), .B(B[3]), .Z(n1949) );
  XNOR U2026 ( .A(n1957), .B(n2088), .Z(n1950) );
  XNOR U2027 ( .A(n1956), .B(n1954), .Z(n2088) );
  AND U2028 ( .A(n2089), .B(n2090), .Z(n1954) );
  NANDN U2029 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U2030 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2031 ( .A(n2094), .B(n2093), .Z(n2089) );
  AND U2032 ( .A(A[16]), .B(B[4]), .Z(n1956) );
  XNOR U2033 ( .A(n1964), .B(n2095), .Z(n1957) );
  XNOR U2034 ( .A(n1963), .B(n1961), .Z(n2095) );
  AND U2035 ( .A(n2096), .B(n2097), .Z(n1961) );
  NANDN U2036 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2037 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2038 ( .A(n2101), .B(n2100), .Z(n2096) );
  AND U2039 ( .A(A[15]), .B(B[5]), .Z(n1963) );
  XNOR U2040 ( .A(n1971), .B(n2102), .Z(n1964) );
  XNOR U2041 ( .A(n1970), .B(n1968), .Z(n2102) );
  AND U2042 ( .A(n2103), .B(n2104), .Z(n1968) );
  NANDN U2043 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2044 ( .A(n2107), .B(n2108), .Z(n2106) );
  NAND U2045 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2046 ( .A(A[14]), .B(B[6]), .Z(n1970) );
  XNOR U2047 ( .A(n1978), .B(n2109), .Z(n1971) );
  XNOR U2048 ( .A(n1977), .B(n1975), .Z(n2109) );
  AND U2049 ( .A(n2110), .B(n2111), .Z(n1975) );
  NANDN U2050 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2051 ( .A(n2114), .B(n2115), .Z(n2113) );
  NANDN U2052 ( .A(n2115), .B(n2114), .Z(n2110) );
  AND U2053 ( .A(A[13]), .B(B[7]), .Z(n1977) );
  XNOR U2054 ( .A(n1985), .B(n2116), .Z(n1978) );
  XNOR U2055 ( .A(n1984), .B(n1982), .Z(n2116) );
  AND U2056 ( .A(n2117), .B(n2118), .Z(n1982) );
  NANDN U2057 ( .A(n2119), .B(n2120), .Z(n2118) );
  OR U2058 ( .A(n2121), .B(n2122), .Z(n2120) );
  NAND U2059 ( .A(n2122), .B(n2121), .Z(n2117) );
  AND U2060 ( .A(A[12]), .B(B[8]), .Z(n1984) );
  XNOR U2061 ( .A(n1992), .B(n2123), .Z(n1985) );
  XNOR U2062 ( .A(n1991), .B(n1989), .Z(n2123) );
  AND U2063 ( .A(n2124), .B(n2125), .Z(n1989) );
  NANDN U2064 ( .A(n2126), .B(n2127), .Z(n2125) );
  NANDN U2065 ( .A(n2128), .B(n2129), .Z(n2127) );
  NANDN U2066 ( .A(n2129), .B(n2128), .Z(n2124) );
  AND U2067 ( .A(A[11]), .B(B[9]), .Z(n1991) );
  XNOR U2068 ( .A(n1999), .B(n2130), .Z(n1992) );
  XNOR U2069 ( .A(n1998), .B(n1996), .Z(n2130) );
  AND U2070 ( .A(n2131), .B(n2132), .Z(n1996) );
  NANDN U2071 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2072 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2073 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2074 ( .A(A[10]), .B(B[10]), .Z(n1998) );
  XNOR U2075 ( .A(n2006), .B(n2137), .Z(n1999) );
  XNOR U2076 ( .A(n2005), .B(n2003), .Z(n2137) );
  AND U2077 ( .A(n2138), .B(n2139), .Z(n2003) );
  NANDN U2078 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U2079 ( .A(n2142), .B(n2143), .Z(n2141) );
  NANDN U2080 ( .A(n2143), .B(n2142), .Z(n2138) );
  AND U2081 ( .A(A[9]), .B(B[11]), .Z(n2005) );
  XNOR U2082 ( .A(n2013), .B(n2144), .Z(n2006) );
  XNOR U2083 ( .A(n2012), .B(n2010), .Z(n2144) );
  AND U2084 ( .A(n2145), .B(n2146), .Z(n2010) );
  NANDN U2085 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2086 ( .A(n2149), .B(n2150), .Z(n2148) );
  NAND U2087 ( .A(n2150), .B(n2149), .Z(n2145) );
  AND U2088 ( .A(A[8]), .B(B[12]), .Z(n2012) );
  XNOR U2089 ( .A(n2020), .B(n2151), .Z(n2013) );
  XNOR U2090 ( .A(n2019), .B(n2017), .Z(n2151) );
  AND U2091 ( .A(n2152), .B(n2153), .Z(n2017) );
  NANDN U2092 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2093 ( .A(n2156), .B(n2157), .Z(n2155) );
  NANDN U2094 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2095 ( .A(A[7]), .B(B[13]), .Z(n2019) );
  XNOR U2096 ( .A(n2027), .B(n2158), .Z(n2020) );
  XNOR U2097 ( .A(n2026), .B(n2024), .Z(n2158) );
  AND U2098 ( .A(n2159), .B(n2160), .Z(n2024) );
  NANDN U2099 ( .A(n2161), .B(n2162), .Z(n2160) );
  OR U2100 ( .A(n2163), .B(n2164), .Z(n2162) );
  NAND U2101 ( .A(n2164), .B(n2163), .Z(n2159) );
  AND U2102 ( .A(A[6]), .B(B[14]), .Z(n2026) );
  XNOR U2103 ( .A(n2034), .B(n2165), .Z(n2027) );
  XNOR U2104 ( .A(n2033), .B(n2031), .Z(n2165) );
  AND U2105 ( .A(n2166), .B(n2167), .Z(n2031) );
  NANDN U2106 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  NANDN U2108 ( .A(n2171), .B(n2170), .Z(n2166) );
  AND U2109 ( .A(A[5]), .B(B[15]), .Z(n2033) );
  XNOR U2110 ( .A(n2041), .B(n2172), .Z(n2034) );
  XNOR U2111 ( .A(n2040), .B(n2038), .Z(n2172) );
  AND U2112 ( .A(n2173), .B(n2174), .Z(n2038) );
  NANDN U2113 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2114 ( .A(n2177), .B(n2178), .Z(n2176) );
  NAND U2115 ( .A(n2178), .B(n2177), .Z(n2173) );
  AND U2116 ( .A(A[4]), .B(B[16]), .Z(n2040) );
  XNOR U2117 ( .A(n2048), .B(n2179), .Z(n2041) );
  XNOR U2118 ( .A(n2047), .B(n2045), .Z(n2179) );
  AND U2119 ( .A(n2180), .B(n2181), .Z(n2045) );
  NANDN U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  NAND U2121 ( .A(n2184), .B(n2185), .Z(n2183) );
  NANDN U2122 ( .A(n2185), .B(n23), .Z(n2180) );
  AND U2123 ( .A(A[3]), .B(B[17]), .Z(n2047) );
  XOR U2124 ( .A(n2054), .B(n2186), .Z(n2048) );
  XNOR U2125 ( .A(n2052), .B(n2055), .Z(n2186) );
  NAND U2126 ( .A(A[2]), .B(B[18]), .Z(n2055) );
  NANDN U2127 ( .A(n2187), .B(n2188), .Z(n2052) );
  AND U2128 ( .A(A[0]), .B(B[19]), .Z(n2188) );
  XNOR U2129 ( .A(n2057), .B(n2189), .Z(n2054) );
  NAND U2130 ( .A(A[0]), .B(B[20]), .Z(n2189) );
  NAND U2131 ( .A(B[19]), .B(A[1]), .Z(n2057) );
  XOR U2132 ( .A(n2066), .B(n2190), .Z(PRODUCT[19]) );
  XNOR U2133 ( .A(n2065), .B(n2063), .Z(n2190) );
  AND U2134 ( .A(n2191), .B(n2192), .Z(n2063) );
  NAND U2135 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U2136 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2137 ( .A(n2196), .B(n2195), .Z(n2191) );
  ANDN U2138 ( .B(A[19]), .A(n42), .Z(n2065) );
  XNOR U2139 ( .A(n2073), .B(n2197), .Z(n2066) );
  XNOR U2140 ( .A(n2072), .B(n2070), .Z(n2197) );
  AND U2141 ( .A(n2198), .B(n2199), .Z(n2070) );
  NANDN U2142 ( .A(n2200), .B(n2201), .Z(n2199) );
  OR U2143 ( .A(n2202), .B(n2203), .Z(n2201) );
  NAND U2144 ( .A(n2203), .B(n2202), .Z(n2198) );
  ANDN U2145 ( .B(A[18]), .A(n41), .Z(n2072) );
  XNOR U2146 ( .A(n2080), .B(n2204), .Z(n2073) );
  XNOR U2147 ( .A(n2079), .B(n2077), .Z(n2204) );
  AND U2148 ( .A(n2205), .B(n2206), .Z(n2077) );
  NANDN U2149 ( .A(n2207), .B(n2208), .Z(n2206) );
  NANDN U2150 ( .A(n2209), .B(n2210), .Z(n2208) );
  NANDN U2151 ( .A(n2210), .B(n2209), .Z(n2205) );
  AND U2152 ( .A(A[17]), .B(B[2]), .Z(n2079) );
  XNOR U2153 ( .A(n2087), .B(n2211), .Z(n2080) );
  XNOR U2154 ( .A(n2086), .B(n2084), .Z(n2211) );
  AND U2155 ( .A(n2212), .B(n2213), .Z(n2084) );
  NANDN U2156 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U2157 ( .A(n2216), .B(n2217), .Z(n2215) );
  NAND U2158 ( .A(n2217), .B(n2216), .Z(n2212) );
  AND U2159 ( .A(A[16]), .B(B[3]), .Z(n2086) );
  XNOR U2160 ( .A(n2094), .B(n2218), .Z(n2087) );
  XNOR U2161 ( .A(n2093), .B(n2091), .Z(n2218) );
  AND U2162 ( .A(n2219), .B(n2220), .Z(n2091) );
  NANDN U2163 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U2164 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2165 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U2166 ( .A(A[15]), .B(B[4]), .Z(n2093) );
  XNOR U2167 ( .A(n2101), .B(n2225), .Z(n2094) );
  XNOR U2168 ( .A(n2100), .B(n2098), .Z(n2225) );
  AND U2169 ( .A(n2226), .B(n2227), .Z(n2098) );
  NANDN U2170 ( .A(n2228), .B(n2229), .Z(n2227) );
  OR U2171 ( .A(n2230), .B(n2231), .Z(n2229) );
  NAND U2172 ( .A(n2231), .B(n2230), .Z(n2226) );
  AND U2173 ( .A(A[14]), .B(B[5]), .Z(n2100) );
  XNOR U2174 ( .A(n2108), .B(n2232), .Z(n2101) );
  XNOR U2175 ( .A(n2107), .B(n2105), .Z(n2232) );
  AND U2176 ( .A(n2233), .B(n2234), .Z(n2105) );
  NANDN U2177 ( .A(n2235), .B(n2236), .Z(n2234) );
  NANDN U2178 ( .A(n2237), .B(n2238), .Z(n2236) );
  NANDN U2179 ( .A(n2238), .B(n2237), .Z(n2233) );
  AND U2180 ( .A(A[13]), .B(B[6]), .Z(n2107) );
  XNOR U2181 ( .A(n2115), .B(n2239), .Z(n2108) );
  XNOR U2182 ( .A(n2114), .B(n2112), .Z(n2239) );
  AND U2183 ( .A(n2240), .B(n2241), .Z(n2112) );
  NANDN U2184 ( .A(n2242), .B(n2243), .Z(n2241) );
  OR U2185 ( .A(n2244), .B(n2245), .Z(n2243) );
  NAND U2186 ( .A(n2245), .B(n2244), .Z(n2240) );
  AND U2187 ( .A(A[12]), .B(B[7]), .Z(n2114) );
  XNOR U2188 ( .A(n2122), .B(n2246), .Z(n2115) );
  XNOR U2189 ( .A(n2121), .B(n2119), .Z(n2246) );
  AND U2190 ( .A(n2247), .B(n2248), .Z(n2119) );
  NANDN U2191 ( .A(n2249), .B(n2250), .Z(n2248) );
  NANDN U2192 ( .A(n2251), .B(n2252), .Z(n2250) );
  NANDN U2193 ( .A(n2252), .B(n2251), .Z(n2247) );
  AND U2194 ( .A(A[11]), .B(B[8]), .Z(n2121) );
  XNOR U2195 ( .A(n2129), .B(n2253), .Z(n2122) );
  XNOR U2196 ( .A(n2128), .B(n2126), .Z(n2253) );
  AND U2197 ( .A(n2254), .B(n2255), .Z(n2126) );
  NANDN U2198 ( .A(n2256), .B(n2257), .Z(n2255) );
  OR U2199 ( .A(n2258), .B(n2259), .Z(n2257) );
  NAND U2200 ( .A(n2259), .B(n2258), .Z(n2254) );
  AND U2201 ( .A(A[10]), .B(B[9]), .Z(n2128) );
  XNOR U2202 ( .A(n2136), .B(n2260), .Z(n2129) );
  XNOR U2203 ( .A(n2135), .B(n2133), .Z(n2260) );
  AND U2204 ( .A(n2261), .B(n2262), .Z(n2133) );
  NANDN U2205 ( .A(n2263), .B(n2264), .Z(n2262) );
  NANDN U2206 ( .A(n2265), .B(n2266), .Z(n2264) );
  NANDN U2207 ( .A(n2266), .B(n2265), .Z(n2261) );
  AND U2208 ( .A(A[9]), .B(B[10]), .Z(n2135) );
  XNOR U2209 ( .A(n2143), .B(n2267), .Z(n2136) );
  XNOR U2210 ( .A(n2142), .B(n2140), .Z(n2267) );
  AND U2211 ( .A(n2268), .B(n2269), .Z(n2140) );
  NANDN U2212 ( .A(n2270), .B(n2271), .Z(n2269) );
  OR U2213 ( .A(n2272), .B(n2273), .Z(n2271) );
  NAND U2214 ( .A(n2273), .B(n2272), .Z(n2268) );
  AND U2215 ( .A(A[8]), .B(B[11]), .Z(n2142) );
  XNOR U2216 ( .A(n2150), .B(n2274), .Z(n2143) );
  XNOR U2217 ( .A(n2149), .B(n2147), .Z(n2274) );
  AND U2218 ( .A(n2275), .B(n2276), .Z(n2147) );
  NANDN U2219 ( .A(n2277), .B(n2278), .Z(n2276) );
  NANDN U2220 ( .A(n2279), .B(n2280), .Z(n2278) );
  NANDN U2221 ( .A(n2280), .B(n2279), .Z(n2275) );
  AND U2222 ( .A(A[7]), .B(B[12]), .Z(n2149) );
  XNOR U2223 ( .A(n2157), .B(n2281), .Z(n2150) );
  XNOR U2224 ( .A(n2156), .B(n2154), .Z(n2281) );
  AND U2225 ( .A(n2282), .B(n2283), .Z(n2154) );
  NANDN U2226 ( .A(n2284), .B(n2285), .Z(n2283) );
  OR U2227 ( .A(n2286), .B(n2287), .Z(n2285) );
  NAND U2228 ( .A(n2287), .B(n2286), .Z(n2282) );
  AND U2229 ( .A(A[6]), .B(B[13]), .Z(n2156) );
  XNOR U2230 ( .A(n2164), .B(n2288), .Z(n2157) );
  XNOR U2231 ( .A(n2163), .B(n2161), .Z(n2288) );
  AND U2232 ( .A(n2289), .B(n2290), .Z(n2161) );
  NANDN U2233 ( .A(n2291), .B(n2292), .Z(n2290) );
  NANDN U2234 ( .A(n2293), .B(n2294), .Z(n2292) );
  NANDN U2235 ( .A(n2294), .B(n2293), .Z(n2289) );
  AND U2236 ( .A(A[5]), .B(B[14]), .Z(n2163) );
  XNOR U2237 ( .A(n2171), .B(n2295), .Z(n2164) );
  XNOR U2238 ( .A(n2170), .B(n2168), .Z(n2295) );
  AND U2239 ( .A(n2296), .B(n2297), .Z(n2168) );
  NANDN U2240 ( .A(n2298), .B(n2299), .Z(n2297) );
  OR U2241 ( .A(n2300), .B(n2301), .Z(n2299) );
  NAND U2242 ( .A(n2301), .B(n2300), .Z(n2296) );
  AND U2243 ( .A(A[4]), .B(B[15]), .Z(n2170) );
  XNOR U2244 ( .A(n2178), .B(n2302), .Z(n2171) );
  XNOR U2245 ( .A(n2177), .B(n2175), .Z(n2302) );
  AND U2246 ( .A(n2303), .B(n2304), .Z(n2175) );
  NANDN U2247 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2248 ( .A(n2307), .B(n2308), .Z(n2306) );
  NANDN U2249 ( .A(n2308), .B(n24), .Z(n2303) );
  AND U2250 ( .A(A[3]), .B(B[16]), .Z(n2177) );
  XOR U2251 ( .A(n2184), .B(n2309), .Z(n2178) );
  XNOR U2252 ( .A(n2182), .B(n2185), .Z(n2309) );
  NAND U2253 ( .A(A[2]), .B(B[17]), .Z(n2185) );
  NANDN U2254 ( .A(n2310), .B(n2311), .Z(n2182) );
  AND U2255 ( .A(A[0]), .B(B[18]), .Z(n2311) );
  XNOR U2256 ( .A(n2187), .B(n2312), .Z(n2184) );
  NAND U2257 ( .A(A[0]), .B(B[19]), .Z(n2312) );
  NAND U2258 ( .A(B[18]), .B(A[1]), .Z(n2187) );
  XOR U2259 ( .A(n2196), .B(n2313), .Z(PRODUCT[18]) );
  XNOR U2260 ( .A(n2195), .B(n2194), .Z(n2313) );
  NAND U2261 ( .A(n2314), .B(n2315), .Z(n2194) );
  NANDN U2262 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2263 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2264 ( .A(n2319), .B(n2318), .Z(n2314) );
  ANDN U2265 ( .B(A[18]), .A(n42), .Z(n2195) );
  XNOR U2266 ( .A(n2203), .B(n2320), .Z(n2196) );
  XNOR U2267 ( .A(n2202), .B(n2200), .Z(n2320) );
  AND U2268 ( .A(n2321), .B(n2322), .Z(n2200) );
  NANDN U2269 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2270 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U2271 ( .A(n2326), .B(n2325), .Z(n2321) );
  ANDN U2272 ( .B(A[17]), .A(n41), .Z(n2202) );
  XNOR U2273 ( .A(n2210), .B(n2327), .Z(n2203) );
  XNOR U2274 ( .A(n2209), .B(n2207), .Z(n2327) );
  AND U2275 ( .A(n2328), .B(n2329), .Z(n2207) );
  NANDN U2276 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR U2277 ( .A(n2332), .B(n2333), .Z(n2331) );
  NAND U2278 ( .A(n2333), .B(n2332), .Z(n2328) );
  AND U2279 ( .A(A[16]), .B(B[2]), .Z(n2209) );
  XNOR U2280 ( .A(n2217), .B(n2334), .Z(n2210) );
  XNOR U2281 ( .A(n2216), .B(n2214), .Z(n2334) );
  AND U2282 ( .A(n2335), .B(n2336), .Z(n2214) );
  NANDN U2283 ( .A(n2337), .B(n2338), .Z(n2336) );
  NANDN U2284 ( .A(n2339), .B(n2340), .Z(n2338) );
  NANDN U2285 ( .A(n2340), .B(n2339), .Z(n2335) );
  AND U2286 ( .A(A[15]), .B(B[3]), .Z(n2216) );
  XNOR U2287 ( .A(n2224), .B(n2341), .Z(n2217) );
  XNOR U2288 ( .A(n2223), .B(n2221), .Z(n2341) );
  AND U2289 ( .A(n2342), .B(n2343), .Z(n2221) );
  NANDN U2290 ( .A(n2344), .B(n2345), .Z(n2343) );
  OR U2291 ( .A(n2346), .B(n2347), .Z(n2345) );
  NAND U2292 ( .A(n2347), .B(n2346), .Z(n2342) );
  AND U2293 ( .A(A[14]), .B(B[4]), .Z(n2223) );
  XNOR U2294 ( .A(n2231), .B(n2348), .Z(n2224) );
  XNOR U2295 ( .A(n2230), .B(n2228), .Z(n2348) );
  AND U2296 ( .A(n2349), .B(n2350), .Z(n2228) );
  NANDN U2297 ( .A(n2351), .B(n2352), .Z(n2350) );
  NANDN U2298 ( .A(n2353), .B(n2354), .Z(n2352) );
  NANDN U2299 ( .A(n2354), .B(n2353), .Z(n2349) );
  AND U2300 ( .A(A[13]), .B(B[5]), .Z(n2230) );
  XNOR U2301 ( .A(n2238), .B(n2355), .Z(n2231) );
  XNOR U2302 ( .A(n2237), .B(n2235), .Z(n2355) );
  AND U2303 ( .A(n2356), .B(n2357), .Z(n2235) );
  NANDN U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U2305 ( .A(n2360), .B(n2361), .Z(n2359) );
  NAND U2306 ( .A(n2361), .B(n2360), .Z(n2356) );
  AND U2307 ( .A(A[12]), .B(B[6]), .Z(n2237) );
  XNOR U2308 ( .A(n2245), .B(n2362), .Z(n2238) );
  XNOR U2309 ( .A(n2244), .B(n2242), .Z(n2362) );
  AND U2310 ( .A(n2363), .B(n2364), .Z(n2242) );
  NANDN U2311 ( .A(n2365), .B(n2366), .Z(n2364) );
  NANDN U2312 ( .A(n2367), .B(n2368), .Z(n2366) );
  NANDN U2313 ( .A(n2368), .B(n2367), .Z(n2363) );
  AND U2314 ( .A(A[11]), .B(B[7]), .Z(n2244) );
  XNOR U2315 ( .A(n2252), .B(n2369), .Z(n2245) );
  XNOR U2316 ( .A(n2251), .B(n2249), .Z(n2369) );
  AND U2317 ( .A(n2370), .B(n2371), .Z(n2249) );
  NANDN U2318 ( .A(n2372), .B(n2373), .Z(n2371) );
  OR U2319 ( .A(n2374), .B(n2375), .Z(n2373) );
  NAND U2320 ( .A(n2375), .B(n2374), .Z(n2370) );
  AND U2321 ( .A(A[10]), .B(B[8]), .Z(n2251) );
  XNOR U2322 ( .A(n2259), .B(n2376), .Z(n2252) );
  XNOR U2323 ( .A(n2258), .B(n2256), .Z(n2376) );
  AND U2324 ( .A(n2377), .B(n2378), .Z(n2256) );
  NANDN U2325 ( .A(n2379), .B(n2380), .Z(n2378) );
  NANDN U2326 ( .A(n2381), .B(n2382), .Z(n2380) );
  NANDN U2327 ( .A(n2382), .B(n2381), .Z(n2377) );
  AND U2328 ( .A(A[9]), .B(B[9]), .Z(n2258) );
  XNOR U2329 ( .A(n2266), .B(n2383), .Z(n2259) );
  XNOR U2330 ( .A(n2265), .B(n2263), .Z(n2383) );
  AND U2331 ( .A(n2384), .B(n2385), .Z(n2263) );
  NANDN U2332 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR U2333 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2334 ( .A(n2389), .B(n2388), .Z(n2384) );
  AND U2335 ( .A(A[8]), .B(B[10]), .Z(n2265) );
  XNOR U2336 ( .A(n2273), .B(n2390), .Z(n2266) );
  XNOR U2337 ( .A(n2272), .B(n2270), .Z(n2390) );
  AND U2338 ( .A(n2391), .B(n2392), .Z(n2270) );
  NANDN U2339 ( .A(n2393), .B(n2394), .Z(n2392) );
  NANDN U2340 ( .A(n2395), .B(n2396), .Z(n2394) );
  NANDN U2341 ( .A(n2396), .B(n2395), .Z(n2391) );
  AND U2342 ( .A(A[7]), .B(B[11]), .Z(n2272) );
  XNOR U2343 ( .A(n2280), .B(n2397), .Z(n2273) );
  XNOR U2344 ( .A(n2279), .B(n2277), .Z(n2397) );
  AND U2345 ( .A(n2398), .B(n2399), .Z(n2277) );
  NANDN U2346 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U2347 ( .A(n2402), .B(n2403), .Z(n2401) );
  NAND U2348 ( .A(n2403), .B(n2402), .Z(n2398) );
  AND U2349 ( .A(A[6]), .B(B[12]), .Z(n2279) );
  XNOR U2350 ( .A(n2287), .B(n2404), .Z(n2280) );
  XNOR U2351 ( .A(n2286), .B(n2284), .Z(n2404) );
  AND U2352 ( .A(n2405), .B(n2406), .Z(n2284) );
  NANDN U2353 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2354 ( .A(n2409), .B(n2410), .Z(n2408) );
  NANDN U2355 ( .A(n2410), .B(n2409), .Z(n2405) );
  AND U2356 ( .A(A[5]), .B(B[13]), .Z(n2286) );
  XNOR U2357 ( .A(n2294), .B(n2411), .Z(n2287) );
  XNOR U2358 ( .A(n2293), .B(n2291), .Z(n2411) );
  AND U2359 ( .A(n2412), .B(n2413), .Z(n2291) );
  NANDN U2360 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2361 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2362 ( .A(n2417), .B(n2416), .Z(n2412) );
  AND U2363 ( .A(A[4]), .B(B[14]), .Z(n2293) );
  XNOR U2364 ( .A(n2301), .B(n2418), .Z(n2294) );
  XNOR U2365 ( .A(n2300), .B(n2298), .Z(n2418) );
  AND U2366 ( .A(n2419), .B(n2420), .Z(n2298) );
  NANDN U2367 ( .A(n2421), .B(n2422), .Z(n2420) );
  NAND U2368 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2369 ( .A(n2424), .B(n25), .Z(n2419) );
  AND U2370 ( .A(A[3]), .B(B[15]), .Z(n2300) );
  XOR U2371 ( .A(n2307), .B(n2425), .Z(n2301) );
  XNOR U2372 ( .A(n2305), .B(n2308), .Z(n2425) );
  NAND U2373 ( .A(A[2]), .B(B[16]), .Z(n2308) );
  NANDN U2374 ( .A(n2426), .B(n2427), .Z(n2305) );
  AND U2375 ( .A(A[0]), .B(B[17]), .Z(n2427) );
  XNOR U2376 ( .A(n2310), .B(n2428), .Z(n2307) );
  NAND U2377 ( .A(A[0]), .B(B[18]), .Z(n2428) );
  NAND U2378 ( .A(B[17]), .B(A[1]), .Z(n2310) );
  XOR U2379 ( .A(n2319), .B(n2429), .Z(PRODUCT[17]) );
  XNOR U2380 ( .A(n2318), .B(n2316), .Z(n2429) );
  AND U2381 ( .A(n2430), .B(n2431), .Z(n2316) );
  NAND U2382 ( .A(n2432), .B(n2433), .Z(n2431) );
  NANDN U2383 ( .A(n2434), .B(n2435), .Z(n2432) );
  NANDN U2384 ( .A(n2435), .B(n2434), .Z(n2430) );
  ANDN U2385 ( .B(A[17]), .A(n42), .Z(n2318) );
  XNOR U2386 ( .A(n2326), .B(n2436), .Z(n2319) );
  XNOR U2387 ( .A(n2325), .B(n2323), .Z(n2436) );
  AND U2388 ( .A(n2437), .B(n2438), .Z(n2323) );
  NANDN U2389 ( .A(n2439), .B(n2440), .Z(n2438) );
  OR U2390 ( .A(n2441), .B(n2442), .Z(n2440) );
  NAND U2391 ( .A(n2442), .B(n2441), .Z(n2437) );
  ANDN U2392 ( .B(A[16]), .A(n41), .Z(n2325) );
  XNOR U2393 ( .A(n2333), .B(n2443), .Z(n2326) );
  XNOR U2394 ( .A(n2332), .B(n2330), .Z(n2443) );
  AND U2395 ( .A(n2444), .B(n2445), .Z(n2330) );
  NANDN U2396 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2397 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U2398 ( .A(n2449), .B(n2448), .Z(n2444) );
  AND U2399 ( .A(A[15]), .B(B[2]), .Z(n2332) );
  XNOR U2400 ( .A(n2340), .B(n2450), .Z(n2333) );
  XNOR U2401 ( .A(n2339), .B(n2337), .Z(n2450) );
  AND U2402 ( .A(n2451), .B(n2452), .Z(n2337) );
  NANDN U2403 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2404 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2405 ( .A(n2456), .B(n2455), .Z(n2451) );
  AND U2406 ( .A(A[14]), .B(B[3]), .Z(n2339) );
  XNOR U2407 ( .A(n2347), .B(n2457), .Z(n2340) );
  XNOR U2408 ( .A(n2346), .B(n2344), .Z(n2457) );
  AND U2409 ( .A(n2458), .B(n2459), .Z(n2344) );
  NANDN U2410 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2411 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U2412 ( .A(n2463), .B(n2462), .Z(n2458) );
  AND U2413 ( .A(A[13]), .B(B[4]), .Z(n2346) );
  XNOR U2414 ( .A(n2354), .B(n2464), .Z(n2347) );
  XNOR U2415 ( .A(n2353), .B(n2351), .Z(n2464) );
  AND U2416 ( .A(n2465), .B(n2466), .Z(n2351) );
  NANDN U2417 ( .A(n2467), .B(n2468), .Z(n2466) );
  OR U2418 ( .A(n2469), .B(n2470), .Z(n2468) );
  NAND U2419 ( .A(n2470), .B(n2469), .Z(n2465) );
  AND U2420 ( .A(A[12]), .B(B[5]), .Z(n2353) );
  XNOR U2421 ( .A(n2361), .B(n2471), .Z(n2354) );
  XNOR U2422 ( .A(n2360), .B(n2358), .Z(n2471) );
  AND U2423 ( .A(n2472), .B(n2473), .Z(n2358) );
  NANDN U2424 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2425 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U2426 ( .A(n2477), .B(n2476), .Z(n2472) );
  AND U2427 ( .A(A[11]), .B(B[6]), .Z(n2360) );
  XNOR U2428 ( .A(n2368), .B(n2478), .Z(n2361) );
  XNOR U2429 ( .A(n2367), .B(n2365), .Z(n2478) );
  AND U2430 ( .A(n2479), .B(n2480), .Z(n2365) );
  NANDN U2431 ( .A(n2481), .B(n2482), .Z(n2480) );
  OR U2432 ( .A(n2483), .B(n2484), .Z(n2482) );
  NAND U2433 ( .A(n2484), .B(n2483), .Z(n2479) );
  AND U2434 ( .A(A[10]), .B(B[7]), .Z(n2367) );
  XNOR U2435 ( .A(n2375), .B(n2485), .Z(n2368) );
  XNOR U2436 ( .A(n2374), .B(n2372), .Z(n2485) );
  AND U2437 ( .A(n2486), .B(n2487), .Z(n2372) );
  NANDN U2438 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2439 ( .A(n2490), .B(n2491), .Z(n2489) );
  NANDN U2440 ( .A(n2491), .B(n2490), .Z(n2486) );
  AND U2441 ( .A(A[9]), .B(B[8]), .Z(n2374) );
  XNOR U2442 ( .A(n2382), .B(n2492), .Z(n2375) );
  XNOR U2443 ( .A(n2381), .B(n2379), .Z(n2492) );
  AND U2444 ( .A(n2493), .B(n2494), .Z(n2379) );
  NANDN U2445 ( .A(n2495), .B(n2496), .Z(n2494) );
  OR U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  NAND U2447 ( .A(n2498), .B(n2497), .Z(n2493) );
  AND U2448 ( .A(A[8]), .B(B[9]), .Z(n2381) );
  XNOR U2449 ( .A(n2389), .B(n2499), .Z(n2382) );
  XNOR U2450 ( .A(n2388), .B(n2386), .Z(n2499) );
  AND U2451 ( .A(n2500), .B(n2501), .Z(n2386) );
  NANDN U2452 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2453 ( .A(n2504), .B(n2505), .Z(n2503) );
  NANDN U2454 ( .A(n2505), .B(n2504), .Z(n2500) );
  AND U2455 ( .A(A[7]), .B(B[10]), .Z(n2388) );
  XNOR U2456 ( .A(n2396), .B(n2506), .Z(n2389) );
  XNOR U2457 ( .A(n2395), .B(n2393), .Z(n2506) );
  AND U2458 ( .A(n2507), .B(n2508), .Z(n2393) );
  NANDN U2459 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U2460 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND U2461 ( .A(n2512), .B(n2511), .Z(n2507) );
  AND U2462 ( .A(A[6]), .B(B[11]), .Z(n2395) );
  XNOR U2463 ( .A(n2403), .B(n2513), .Z(n2396) );
  XNOR U2464 ( .A(n2402), .B(n2400), .Z(n2513) );
  AND U2465 ( .A(n2514), .B(n2515), .Z(n2400) );
  NANDN U2466 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2467 ( .A(n2518), .B(n2519), .Z(n2517) );
  NANDN U2468 ( .A(n2519), .B(n2518), .Z(n2514) );
  AND U2469 ( .A(A[5]), .B(B[12]), .Z(n2402) );
  XNOR U2470 ( .A(n2410), .B(n2520), .Z(n2403) );
  XNOR U2471 ( .A(n2409), .B(n2407), .Z(n2520) );
  AND U2472 ( .A(n2521), .B(n2522), .Z(n2407) );
  NANDN U2473 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U2474 ( .A(n2525), .B(n2526), .Z(n2524) );
  NAND U2475 ( .A(n2526), .B(n2525), .Z(n2521) );
  AND U2476 ( .A(A[4]), .B(B[13]), .Z(n2409) );
  XNOR U2477 ( .A(n2417), .B(n2527), .Z(n2410) );
  XNOR U2478 ( .A(n2416), .B(n2414), .Z(n2527) );
  AND U2479 ( .A(n2528), .B(n2529), .Z(n2414) );
  NANDN U2480 ( .A(n2530), .B(n2531), .Z(n2529) );
  NAND U2481 ( .A(n2532), .B(n2533), .Z(n2531) );
  NANDN U2482 ( .A(n2533), .B(n26), .Z(n2528) );
  AND U2483 ( .A(A[3]), .B(B[14]), .Z(n2416) );
  XOR U2484 ( .A(n2423), .B(n2534), .Z(n2417) );
  XNOR U2485 ( .A(n2421), .B(n2424), .Z(n2534) );
  NAND U2486 ( .A(A[2]), .B(B[15]), .Z(n2424) );
  NANDN U2487 ( .A(n2535), .B(n2536), .Z(n2421) );
  AND U2488 ( .A(A[0]), .B(B[16]), .Z(n2536) );
  XNOR U2489 ( .A(n2426), .B(n2537), .Z(n2423) );
  NAND U2490 ( .A(A[0]), .B(B[17]), .Z(n2537) );
  NAND U2491 ( .A(B[16]), .B(A[1]), .Z(n2426) );
  XOR U2492 ( .A(n2435), .B(n2538), .Z(PRODUCT[16]) );
  XNOR U2493 ( .A(n2434), .B(n2433), .Z(n2538) );
  NAND U2494 ( .A(n2539), .B(n2540), .Z(n2433) );
  NANDN U2495 ( .A(n2541), .B(n2542), .Z(n2540) );
  OR U2496 ( .A(n2543), .B(n2544), .Z(n2542) );
  NAND U2497 ( .A(n2544), .B(n2543), .Z(n2539) );
  ANDN U2498 ( .B(A[16]), .A(n42), .Z(n2434) );
  XNOR U2499 ( .A(n2442), .B(n2545), .Z(n2435) );
  XNOR U2500 ( .A(n2441), .B(n2439), .Z(n2545) );
  AND U2501 ( .A(n2546), .B(n2547), .Z(n2439) );
  NANDN U2502 ( .A(n2548), .B(n2549), .Z(n2547) );
  NANDN U2503 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2504 ( .A(n2551), .B(n2550), .Z(n2546) );
  ANDN U2505 ( .B(A[15]), .A(n41), .Z(n2441) );
  XNOR U2506 ( .A(n2449), .B(n2552), .Z(n2442) );
  XNOR U2507 ( .A(n2448), .B(n2446), .Z(n2552) );
  AND U2508 ( .A(n2553), .B(n2554), .Z(n2446) );
  NANDN U2509 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2510 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2511 ( .A(n2558), .B(n2557), .Z(n2553) );
  AND U2512 ( .A(A[14]), .B(B[2]), .Z(n2448) );
  XNOR U2513 ( .A(n2456), .B(n2559), .Z(n2449) );
  XNOR U2514 ( .A(n2455), .B(n2453), .Z(n2559) );
  AND U2515 ( .A(n2560), .B(n2561), .Z(n2453) );
  NANDN U2516 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2517 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2518 ( .A(n2565), .B(n2564), .Z(n2560) );
  AND U2519 ( .A(A[13]), .B(B[3]), .Z(n2455) );
  XNOR U2520 ( .A(n2463), .B(n2566), .Z(n2456) );
  XNOR U2521 ( .A(n2462), .B(n2460), .Z(n2566) );
  AND U2522 ( .A(n2567), .B(n2568), .Z(n2460) );
  NANDN U2523 ( .A(n2569), .B(n2570), .Z(n2568) );
  OR U2524 ( .A(n2571), .B(n2572), .Z(n2570) );
  NAND U2525 ( .A(n2572), .B(n2571), .Z(n2567) );
  AND U2526 ( .A(A[12]), .B(B[4]), .Z(n2462) );
  XNOR U2527 ( .A(n2470), .B(n2573), .Z(n2463) );
  XNOR U2528 ( .A(n2469), .B(n2467), .Z(n2573) );
  AND U2529 ( .A(n2574), .B(n2575), .Z(n2467) );
  NANDN U2530 ( .A(n2576), .B(n2577), .Z(n2575) );
  NANDN U2531 ( .A(n2578), .B(n2579), .Z(n2577) );
  NANDN U2532 ( .A(n2579), .B(n2578), .Z(n2574) );
  AND U2533 ( .A(A[11]), .B(B[5]), .Z(n2469) );
  XNOR U2534 ( .A(n2477), .B(n2580), .Z(n2470) );
  XNOR U2535 ( .A(n2476), .B(n2474), .Z(n2580) );
  AND U2536 ( .A(n2581), .B(n2582), .Z(n2474) );
  NANDN U2537 ( .A(n2583), .B(n2584), .Z(n2582) );
  OR U2538 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2539 ( .A(n2586), .B(n2585), .Z(n2581) );
  AND U2540 ( .A(A[10]), .B(B[6]), .Z(n2476) );
  XNOR U2541 ( .A(n2484), .B(n2587), .Z(n2477) );
  XNOR U2542 ( .A(n2483), .B(n2481), .Z(n2587) );
  AND U2543 ( .A(n2588), .B(n2589), .Z(n2481) );
  NANDN U2544 ( .A(n2590), .B(n2591), .Z(n2589) );
  NANDN U2545 ( .A(n2592), .B(n2593), .Z(n2591) );
  NANDN U2546 ( .A(n2593), .B(n2592), .Z(n2588) );
  AND U2547 ( .A(A[9]), .B(B[7]), .Z(n2483) );
  XNOR U2548 ( .A(n2491), .B(n2594), .Z(n2484) );
  XNOR U2549 ( .A(n2490), .B(n2488), .Z(n2594) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2488) );
  NANDN U2551 ( .A(n2597), .B(n2598), .Z(n2596) );
  OR U2552 ( .A(n2599), .B(n2600), .Z(n2598) );
  NAND U2553 ( .A(n2600), .B(n2599), .Z(n2595) );
  AND U2554 ( .A(A[8]), .B(B[8]), .Z(n2490) );
  XNOR U2555 ( .A(n2498), .B(n2601), .Z(n2491) );
  XNOR U2556 ( .A(n2497), .B(n2495), .Z(n2601) );
  AND U2557 ( .A(n2602), .B(n2603), .Z(n2495) );
  NANDN U2558 ( .A(n2604), .B(n2605), .Z(n2603) );
  NANDN U2559 ( .A(n2606), .B(n2607), .Z(n2605) );
  NANDN U2560 ( .A(n2607), .B(n2606), .Z(n2602) );
  AND U2561 ( .A(A[7]), .B(B[9]), .Z(n2497) );
  XNOR U2562 ( .A(n2505), .B(n2608), .Z(n2498) );
  XNOR U2563 ( .A(n2504), .B(n2502), .Z(n2608) );
  AND U2564 ( .A(n2609), .B(n2610), .Z(n2502) );
  NANDN U2565 ( .A(n2611), .B(n2612), .Z(n2610) );
  OR U2566 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND U2567 ( .A(n2614), .B(n2613), .Z(n2609) );
  AND U2568 ( .A(A[6]), .B(B[10]), .Z(n2504) );
  XNOR U2569 ( .A(n2512), .B(n2615), .Z(n2505) );
  XNOR U2570 ( .A(n2511), .B(n2509), .Z(n2615) );
  AND U2571 ( .A(n2616), .B(n2617), .Z(n2509) );
  NANDN U2572 ( .A(n2618), .B(n2619), .Z(n2617) );
  NANDN U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  NANDN U2574 ( .A(n2621), .B(n2620), .Z(n2616) );
  AND U2575 ( .A(A[5]), .B(B[11]), .Z(n2511) );
  XNOR U2576 ( .A(n2519), .B(n2622), .Z(n2512) );
  XNOR U2577 ( .A(n2518), .B(n2516), .Z(n2622) );
  AND U2578 ( .A(n2623), .B(n2624), .Z(n2516) );
  NANDN U2579 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR U2580 ( .A(n2627), .B(n2628), .Z(n2626) );
  NAND U2581 ( .A(n2628), .B(n2627), .Z(n2623) );
  AND U2582 ( .A(A[4]), .B(B[12]), .Z(n2518) );
  XNOR U2583 ( .A(n2526), .B(n2629), .Z(n2519) );
  XNOR U2584 ( .A(n2525), .B(n2523), .Z(n2629) );
  AND U2585 ( .A(n2630), .B(n2631), .Z(n2523) );
  NANDN U2586 ( .A(n2632), .B(n2633), .Z(n2631) );
  NAND U2587 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U2588 ( .A(n2635), .B(n27), .Z(n2630) );
  AND U2589 ( .A(A[3]), .B(B[13]), .Z(n2525) );
  XOR U2590 ( .A(n2532), .B(n2636), .Z(n2526) );
  XNOR U2591 ( .A(n2530), .B(n2533), .Z(n2636) );
  NAND U2592 ( .A(A[2]), .B(B[14]), .Z(n2533) );
  NANDN U2593 ( .A(n2637), .B(n2638), .Z(n2530) );
  AND U2594 ( .A(A[0]), .B(B[15]), .Z(n2638) );
  XNOR U2595 ( .A(n2535), .B(n2639), .Z(n2532) );
  NAND U2596 ( .A(A[0]), .B(B[16]), .Z(n2639) );
  NAND U2597 ( .A(B[15]), .B(A[1]), .Z(n2535) );
  XOR U2598 ( .A(n2544), .B(n2640), .Z(PRODUCT[15]) );
  XNOR U2599 ( .A(n2543), .B(n2541), .Z(n2640) );
  AND U2600 ( .A(n2641), .B(n2642), .Z(n2541) );
  NAND U2601 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2602 ( .A(n2645), .B(n2646), .Z(n2643) );
  NANDN U2603 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2604 ( .B(A[15]), .A(n42), .Z(n2543) );
  XNOR U2605 ( .A(n2551), .B(n2647), .Z(n2544) );
  XNOR U2606 ( .A(n2550), .B(n2548), .Z(n2647) );
  AND U2607 ( .A(n2648), .B(n2649), .Z(n2548) );
  NANDN U2608 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2609 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2610 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2611 ( .B(A[14]), .A(n41), .Z(n2550) );
  XNOR U2612 ( .A(n2558), .B(n2654), .Z(n2551) );
  XNOR U2613 ( .A(n2557), .B(n2555), .Z(n2654) );
  AND U2614 ( .A(n2655), .B(n2656), .Z(n2555) );
  NANDN U2615 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2616 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2617 ( .A(n2660), .B(n2659), .Z(n2655) );
  AND U2618 ( .A(A[13]), .B(B[2]), .Z(n2557) );
  XNOR U2619 ( .A(n2565), .B(n2661), .Z(n2558) );
  XNOR U2620 ( .A(n2564), .B(n2562), .Z(n2661) );
  AND U2621 ( .A(n2662), .B(n2663), .Z(n2562) );
  NANDN U2622 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2623 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2624 ( .A(n2667), .B(n2666), .Z(n2662) );
  AND U2625 ( .A(A[12]), .B(B[3]), .Z(n2564) );
  XNOR U2626 ( .A(n2572), .B(n2668), .Z(n2565) );
  XNOR U2627 ( .A(n2571), .B(n2569), .Z(n2668) );
  AND U2628 ( .A(n2669), .B(n2670), .Z(n2569) );
  NANDN U2629 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2630 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2631 ( .A(n2674), .B(n2673), .Z(n2669) );
  AND U2632 ( .A(A[11]), .B(B[4]), .Z(n2571) );
  XNOR U2633 ( .A(n2579), .B(n2675), .Z(n2572) );
  XNOR U2634 ( .A(n2578), .B(n2576), .Z(n2675) );
  AND U2635 ( .A(n2676), .B(n2677), .Z(n2576) );
  NANDN U2636 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2637 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2638 ( .A(n2681), .B(n2680), .Z(n2676) );
  AND U2639 ( .A(A[10]), .B(B[5]), .Z(n2578) );
  XNOR U2640 ( .A(n2586), .B(n2682), .Z(n2579) );
  XNOR U2641 ( .A(n2585), .B(n2583), .Z(n2682) );
  AND U2642 ( .A(n2683), .B(n2684), .Z(n2583) );
  NANDN U2643 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2644 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2645 ( .A(n2688), .B(n2687), .Z(n2683) );
  AND U2646 ( .A(A[9]), .B(B[6]), .Z(n2585) );
  XNOR U2647 ( .A(n2593), .B(n2689), .Z(n2586) );
  XNOR U2648 ( .A(n2592), .B(n2590), .Z(n2689) );
  AND U2649 ( .A(n2690), .B(n2691), .Z(n2590) );
  NANDN U2650 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2651 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2652 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U2653 ( .A(A[8]), .B(B[7]), .Z(n2592) );
  XNOR U2654 ( .A(n2600), .B(n2696), .Z(n2593) );
  XNOR U2655 ( .A(n2599), .B(n2597), .Z(n2696) );
  AND U2656 ( .A(n2697), .B(n2698), .Z(n2597) );
  NANDN U2657 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2658 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2659 ( .A(n2702), .B(n2701), .Z(n2697) );
  AND U2660 ( .A(A[7]), .B(B[8]), .Z(n2599) );
  XNOR U2661 ( .A(n2607), .B(n2703), .Z(n2600) );
  XNOR U2662 ( .A(n2606), .B(n2604), .Z(n2703) );
  AND U2663 ( .A(n2704), .B(n2705), .Z(n2604) );
  NANDN U2664 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2665 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2666 ( .A(n2709), .B(n2708), .Z(n2704) );
  AND U2667 ( .A(A[6]), .B(B[9]), .Z(n2606) );
  XNOR U2668 ( .A(n2614), .B(n2710), .Z(n2607) );
  XNOR U2669 ( .A(n2613), .B(n2611), .Z(n2710) );
  AND U2670 ( .A(n2711), .B(n2712), .Z(n2611) );
  NANDN U2671 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2672 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2673 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U2674 ( .A(A[5]), .B(B[10]), .Z(n2613) );
  XNOR U2675 ( .A(n2621), .B(n2717), .Z(n2614) );
  XNOR U2676 ( .A(n2620), .B(n2618), .Z(n2717) );
  AND U2677 ( .A(n2718), .B(n2719), .Z(n2618) );
  NANDN U2678 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2679 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2680 ( .A(n2723), .B(n2722), .Z(n2718) );
  AND U2681 ( .A(A[4]), .B(B[11]), .Z(n2620) );
  XNOR U2682 ( .A(n2628), .B(n2724), .Z(n2621) );
  XNOR U2683 ( .A(n2627), .B(n2625), .Z(n2724) );
  AND U2684 ( .A(n2725), .B(n2726), .Z(n2625) );
  NANDN U2685 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2686 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2687 ( .A(n2730), .B(n28), .Z(n2725) );
  AND U2688 ( .A(A[3]), .B(B[12]), .Z(n2627) );
  XOR U2689 ( .A(n2634), .B(n2731), .Z(n2628) );
  XNOR U2690 ( .A(n2632), .B(n2635), .Z(n2731) );
  NAND U2691 ( .A(A[2]), .B(B[13]), .Z(n2635) );
  NANDN U2692 ( .A(n2732), .B(n2733), .Z(n2632) );
  AND U2693 ( .A(A[0]), .B(B[14]), .Z(n2733) );
  XNOR U2694 ( .A(n2637), .B(n2734), .Z(n2634) );
  NAND U2695 ( .A(A[0]), .B(B[15]), .Z(n2734) );
  NAND U2696 ( .A(B[14]), .B(A[1]), .Z(n2637) );
  XOR U2697 ( .A(n2646), .B(n2735), .Z(PRODUCT[14]) );
  XNOR U2698 ( .A(n2645), .B(n2644), .Z(n2735) );
  NAND U2699 ( .A(n2736), .B(n2737), .Z(n2644) );
  NANDN U2700 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U2701 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND U2702 ( .A(n2741), .B(n2740), .Z(n2736) );
  ANDN U2703 ( .B(A[14]), .A(n42), .Z(n2645) );
  XNOR U2704 ( .A(n2653), .B(n2742), .Z(n2646) );
  XNOR U2705 ( .A(n2652), .B(n2650), .Z(n2742) );
  AND U2706 ( .A(n2743), .B(n2744), .Z(n2650) );
  NANDN U2707 ( .A(n2745), .B(n2746), .Z(n2744) );
  NANDN U2708 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2709 ( .A(n2748), .B(n2747), .Z(n2743) );
  ANDN U2710 ( .B(A[13]), .A(n41), .Z(n2652) );
  XNOR U2711 ( .A(n2660), .B(n2749), .Z(n2653) );
  XNOR U2712 ( .A(n2659), .B(n2657), .Z(n2749) );
  AND U2713 ( .A(n2750), .B(n2751), .Z(n2657) );
  NANDN U2714 ( .A(n2752), .B(n2753), .Z(n2751) );
  OR U2715 ( .A(n2754), .B(n2755), .Z(n2753) );
  NAND U2716 ( .A(n2755), .B(n2754), .Z(n2750) );
  AND U2717 ( .A(A[12]), .B(B[2]), .Z(n2659) );
  XNOR U2718 ( .A(n2667), .B(n2756), .Z(n2660) );
  XNOR U2719 ( .A(n2666), .B(n2664), .Z(n2756) );
  AND U2720 ( .A(n2757), .B(n2758), .Z(n2664) );
  NANDN U2721 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2723 ( .A(n2762), .B(n2761), .Z(n2757) );
  AND U2724 ( .A(A[11]), .B(B[3]), .Z(n2666) );
  XNOR U2725 ( .A(n2674), .B(n2763), .Z(n2667) );
  XNOR U2726 ( .A(n2673), .B(n2671), .Z(n2763) );
  AND U2727 ( .A(n2764), .B(n2765), .Z(n2671) );
  NANDN U2728 ( .A(n2766), .B(n2767), .Z(n2765) );
  OR U2729 ( .A(n2768), .B(n2769), .Z(n2767) );
  NAND U2730 ( .A(n2769), .B(n2768), .Z(n2764) );
  AND U2731 ( .A(A[10]), .B(B[4]), .Z(n2673) );
  XNOR U2732 ( .A(n2681), .B(n2770), .Z(n2674) );
  XNOR U2733 ( .A(n2680), .B(n2678), .Z(n2770) );
  AND U2734 ( .A(n2771), .B(n2772), .Z(n2678) );
  NANDN U2735 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2736 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2737 ( .A(n2776), .B(n2775), .Z(n2771) );
  AND U2738 ( .A(A[9]), .B(B[5]), .Z(n2680) );
  XNOR U2739 ( .A(n2688), .B(n2777), .Z(n2681) );
  XNOR U2740 ( .A(n2687), .B(n2685), .Z(n2777) );
  AND U2741 ( .A(n2778), .B(n2779), .Z(n2685) );
  NANDN U2742 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U2743 ( .A(n2782), .B(n2783), .Z(n2781) );
  NAND U2744 ( .A(n2783), .B(n2782), .Z(n2778) );
  AND U2745 ( .A(A[8]), .B(B[6]), .Z(n2687) );
  XNOR U2746 ( .A(n2695), .B(n2784), .Z(n2688) );
  XNOR U2747 ( .A(n2694), .B(n2692), .Z(n2784) );
  AND U2748 ( .A(n2785), .B(n2786), .Z(n2692) );
  NANDN U2749 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2750 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2751 ( .A(n2790), .B(n2789), .Z(n2785) );
  AND U2752 ( .A(A[7]), .B(B[7]), .Z(n2694) );
  XNOR U2753 ( .A(n2702), .B(n2791), .Z(n2695) );
  XNOR U2754 ( .A(n2701), .B(n2699), .Z(n2791) );
  AND U2755 ( .A(n2792), .B(n2793), .Z(n2699) );
  NANDN U2756 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U2757 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2758 ( .A(n2797), .B(n2796), .Z(n2792) );
  AND U2759 ( .A(A[6]), .B(B[8]), .Z(n2701) );
  XNOR U2760 ( .A(n2709), .B(n2798), .Z(n2702) );
  XNOR U2761 ( .A(n2708), .B(n2706), .Z(n2798) );
  AND U2762 ( .A(n2799), .B(n2800), .Z(n2706) );
  NANDN U2763 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2764 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2765 ( .A(n2804), .B(n2803), .Z(n2799) );
  AND U2766 ( .A(A[5]), .B(B[9]), .Z(n2708) );
  XNOR U2767 ( .A(n2716), .B(n2805), .Z(n2709) );
  XNOR U2768 ( .A(n2715), .B(n2713), .Z(n2805) );
  AND U2769 ( .A(n2806), .B(n2807), .Z(n2713) );
  NANDN U2770 ( .A(n2808), .B(n2809), .Z(n2807) );
  OR U2771 ( .A(n2810), .B(n2811), .Z(n2809) );
  NAND U2772 ( .A(n2811), .B(n2810), .Z(n2806) );
  AND U2773 ( .A(A[4]), .B(B[10]), .Z(n2715) );
  XNOR U2774 ( .A(n2723), .B(n2812), .Z(n2716) );
  XNOR U2775 ( .A(n2722), .B(n2720), .Z(n2812) );
  AND U2776 ( .A(n2813), .B(n2814), .Z(n2720) );
  NANDN U2777 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U2778 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2779 ( .A(n2818), .B(n29), .Z(n2813) );
  AND U2780 ( .A(A[3]), .B(B[11]), .Z(n2722) );
  XOR U2781 ( .A(n2729), .B(n2819), .Z(n2723) );
  XNOR U2782 ( .A(n2727), .B(n2730), .Z(n2819) );
  NAND U2783 ( .A(A[2]), .B(B[12]), .Z(n2730) );
  NANDN U2784 ( .A(n2820), .B(n2821), .Z(n2727) );
  AND U2785 ( .A(A[0]), .B(B[13]), .Z(n2821) );
  XNOR U2786 ( .A(n2732), .B(n2822), .Z(n2729) );
  NAND U2787 ( .A(A[0]), .B(B[14]), .Z(n2822) );
  NAND U2788 ( .A(B[13]), .B(A[1]), .Z(n2732) );
  XOR U2789 ( .A(n2741), .B(n2823), .Z(PRODUCT[13]) );
  XNOR U2790 ( .A(n2740), .B(n2738), .Z(n2823) );
  AND U2791 ( .A(n2824), .B(n2825), .Z(n2738) );
  NANDN U2792 ( .A(n2826), .B(n2827), .Z(n2825) );
  NANDN U2793 ( .A(n2828), .B(n2829), .Z(n2827) );
  NANDN U2794 ( .A(n2829), .B(n2828), .Z(n2824) );
  ANDN U2795 ( .B(A[13]), .A(n42), .Z(n2740) );
  XNOR U2796 ( .A(n2748), .B(n2830), .Z(n2741) );
  XNOR U2797 ( .A(n2747), .B(n2745), .Z(n2830) );
  AND U2798 ( .A(n2831), .B(n2832), .Z(n2745) );
  NANDN U2799 ( .A(n2833), .B(n2834), .Z(n2832) );
  OR U2800 ( .A(n2835), .B(n2836), .Z(n2834) );
  NAND U2801 ( .A(n2836), .B(n2835), .Z(n2831) );
  ANDN U2802 ( .B(A[12]), .A(n41), .Z(n2747) );
  XNOR U2803 ( .A(n2755), .B(n2837), .Z(n2748) );
  XNOR U2804 ( .A(n2754), .B(n2752), .Z(n2837) );
  AND U2805 ( .A(n2838), .B(n2839), .Z(n2752) );
  NANDN U2806 ( .A(n2840), .B(n2841), .Z(n2839) );
  NANDN U2807 ( .A(n2842), .B(n2843), .Z(n2841) );
  NANDN U2808 ( .A(n2843), .B(n2842), .Z(n2838) );
  AND U2809 ( .A(A[11]), .B(B[2]), .Z(n2754) );
  XNOR U2810 ( .A(n2762), .B(n2844), .Z(n2755) );
  XNOR U2811 ( .A(n2761), .B(n2759), .Z(n2844) );
  AND U2812 ( .A(n2845), .B(n2846), .Z(n2759) );
  NANDN U2813 ( .A(n2847), .B(n2848), .Z(n2846) );
  OR U2814 ( .A(n2849), .B(n2850), .Z(n2848) );
  NAND U2815 ( .A(n2850), .B(n2849), .Z(n2845) );
  AND U2816 ( .A(A[10]), .B(B[3]), .Z(n2761) );
  XNOR U2817 ( .A(n2769), .B(n2851), .Z(n2762) );
  XNOR U2818 ( .A(n2768), .B(n2766), .Z(n2851) );
  AND U2819 ( .A(n2852), .B(n2853), .Z(n2766) );
  NANDN U2820 ( .A(n2854), .B(n2855), .Z(n2853) );
  NANDN U2821 ( .A(n2856), .B(n2857), .Z(n2855) );
  NANDN U2822 ( .A(n2857), .B(n2856), .Z(n2852) );
  AND U2823 ( .A(A[9]), .B(B[4]), .Z(n2768) );
  XNOR U2824 ( .A(n2776), .B(n2858), .Z(n2769) );
  XNOR U2825 ( .A(n2775), .B(n2773), .Z(n2858) );
  AND U2826 ( .A(n2859), .B(n2860), .Z(n2773) );
  NANDN U2827 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2828 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2829 ( .A(n2864), .B(n2863), .Z(n2859) );
  AND U2830 ( .A(A[8]), .B(B[5]), .Z(n2775) );
  XNOR U2831 ( .A(n2783), .B(n2865), .Z(n2776) );
  XNOR U2832 ( .A(n2782), .B(n2780), .Z(n2865) );
  AND U2833 ( .A(n2866), .B(n2867), .Z(n2780) );
  NANDN U2834 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2835 ( .A(n2870), .B(n2871), .Z(n2869) );
  NANDN U2836 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U2837 ( .A(A[7]), .B(B[6]), .Z(n2782) );
  XNOR U2838 ( .A(n2790), .B(n2872), .Z(n2783) );
  XNOR U2839 ( .A(n2789), .B(n2787), .Z(n2872) );
  AND U2840 ( .A(n2873), .B(n2874), .Z(n2787) );
  NANDN U2841 ( .A(n2875), .B(n2876), .Z(n2874) );
  OR U2842 ( .A(n2877), .B(n2878), .Z(n2876) );
  NAND U2843 ( .A(n2878), .B(n2877), .Z(n2873) );
  AND U2844 ( .A(A[6]), .B(B[7]), .Z(n2789) );
  XNOR U2845 ( .A(n2797), .B(n2879), .Z(n2790) );
  XNOR U2846 ( .A(n2796), .B(n2794), .Z(n2879) );
  AND U2847 ( .A(n2880), .B(n2881), .Z(n2794) );
  NANDN U2848 ( .A(n2882), .B(n2883), .Z(n2881) );
  NANDN U2849 ( .A(n2884), .B(n2885), .Z(n2883) );
  NANDN U2850 ( .A(n2885), .B(n2884), .Z(n2880) );
  AND U2851 ( .A(A[5]), .B(B[8]), .Z(n2796) );
  XNOR U2852 ( .A(n2804), .B(n2886), .Z(n2797) );
  XNOR U2853 ( .A(n2803), .B(n2801), .Z(n2886) );
  AND U2854 ( .A(n2887), .B(n2888), .Z(n2801) );
  NANDN U2855 ( .A(n2889), .B(n2890), .Z(n2888) );
  OR U2856 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2857 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U2858 ( .A(A[4]), .B(B[9]), .Z(n2803) );
  XNOR U2859 ( .A(n2811), .B(n2893), .Z(n2804) );
  XNOR U2860 ( .A(n2810), .B(n2808), .Z(n2893) );
  AND U2861 ( .A(n2894), .B(n2895), .Z(n2808) );
  NANDN U2862 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2863 ( .A(n2898), .B(n2899), .Z(n2897) );
  NANDN U2864 ( .A(n2899), .B(n39), .Z(n2894) );
  AND U2865 ( .A(A[3]), .B(B[10]), .Z(n2810) );
  XOR U2866 ( .A(n2817), .B(n2900), .Z(n2811) );
  XNOR U2867 ( .A(n2815), .B(n2818), .Z(n2900) );
  NAND U2868 ( .A(A[2]), .B(B[11]), .Z(n2818) );
  NANDN U2869 ( .A(n2901), .B(n2902), .Z(n2815) );
  AND U2870 ( .A(A[0]), .B(B[12]), .Z(n2902) );
  XNOR U2871 ( .A(n2820), .B(n2903), .Z(n2817) );
  NAND U2872 ( .A(A[0]), .B(B[13]), .Z(n2903) );
  NAND U2873 ( .A(B[12]), .B(A[1]), .Z(n2820) );
  XNOR U2874 ( .A(n2828), .B(n2904), .Z(PRODUCT[12]) );
  XNOR U2875 ( .A(n2826), .B(n2829), .Z(n2904) );
  AND U2876 ( .A(n2905), .B(n2906), .Z(n2829) );
  NANDN U2877 ( .A(n47), .B(n2907), .Z(n2906) );
  NANDN U2878 ( .A(n45), .B(n2908), .Z(n2907) );
  NAND U2879 ( .A(B[0]), .B(A[11]), .Z(n47) );
  NAND U2880 ( .A(n4), .B(n45), .Z(n2905) );
  XOR U2881 ( .A(n2909), .B(n2910), .Z(n45) );
  XNOR U2882 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2883 ( .A(n2913), .B(n2914), .Z(n2908) );
  NANDN U2884 ( .A(n50), .B(n2915), .Z(n2914) );
  NANDN U2885 ( .A(n48), .B(n51), .Z(n2915) );
  NAND U2886 ( .A(B[0]), .B(A[10]), .Z(n50) );
  NANDN U2887 ( .A(n51), .B(n48), .Z(n2913) );
  XOR U2888 ( .A(n2916), .B(n2917), .Z(n48) );
  XNOR U2889 ( .A(n2918), .B(n2919), .Z(n2917) );
  AND U2890 ( .A(n2920), .B(n2921), .Z(n51) );
  NANDN U2891 ( .A(n54), .B(n2922), .Z(n2921) );
  NANDN U2892 ( .A(n52), .B(n2923), .Z(n2922) );
  NAND U2893 ( .A(B[0]), .B(A[9]), .Z(n54) );
  NAND U2894 ( .A(n6), .B(n52), .Z(n2920) );
  XOR U2895 ( .A(n2924), .B(n2925), .Z(n52) );
  XNOR U2896 ( .A(n2926), .B(n2927), .Z(n2925) );
  AND U2897 ( .A(n2928), .B(n2929), .Z(n2923) );
  NANDN U2898 ( .A(n57), .B(n2930), .Z(n2929) );
  NANDN U2899 ( .A(n55), .B(n58), .Z(n2930) );
  NAND U2900 ( .A(B[0]), .B(A[8]), .Z(n57) );
  NANDN U2901 ( .A(n58), .B(n55), .Z(n2928) );
  XOR U2902 ( .A(n2931), .B(n2932), .Z(n55) );
  XNOR U2903 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2904 ( .A(n2935), .B(n2936), .Z(n58) );
  NANDN U2905 ( .A(n61), .B(n2937), .Z(n2936) );
  NANDN U2906 ( .A(n59), .B(n2938), .Z(n2937) );
  NAND U2907 ( .A(B[0]), .B(A[7]), .Z(n61) );
  NAND U2908 ( .A(n8), .B(n59), .Z(n2935) );
  XOR U2909 ( .A(n2939), .B(n2940), .Z(n59) );
  XNOR U2910 ( .A(n2941), .B(n2942), .Z(n2940) );
  AND U2911 ( .A(n2943), .B(n2944), .Z(n2938) );
  NANDN U2912 ( .A(n64), .B(n2945), .Z(n2944) );
  NANDN U2913 ( .A(n62), .B(n65), .Z(n2945) );
  NAND U2914 ( .A(B[0]), .B(A[6]), .Z(n64) );
  NANDN U2915 ( .A(n65), .B(n62), .Z(n2943) );
  XOR U2916 ( .A(n2946), .B(n2947), .Z(n62) );
  XNOR U2917 ( .A(n2948), .B(n2949), .Z(n2947) );
  AND U2918 ( .A(n2950), .B(n2951), .Z(n65) );
  NANDN U2919 ( .A(n68), .B(n2952), .Z(n2951) );
  NANDN U2920 ( .A(n66), .B(n2953), .Z(n2952) );
  NAND U2921 ( .A(B[0]), .B(A[5]), .Z(n68) );
  NAND U2922 ( .A(n10), .B(n66), .Z(n2950) );
  XOR U2923 ( .A(n2954), .B(n2955), .Z(n66) );
  XNOR U2924 ( .A(n2956), .B(n2957), .Z(n2955) );
  AND U2925 ( .A(n2958), .B(n2959), .Z(n2953) );
  NANDN U2926 ( .A(n162), .B(n2960), .Z(n2959) );
  NANDN U2927 ( .A(n160), .B(n163), .Z(n2960) );
  NAND U2928 ( .A(B[0]), .B(A[4]), .Z(n162) );
  NANDN U2929 ( .A(n163), .B(n160), .Z(n2958) );
  XOR U2930 ( .A(n2961), .B(n2962), .Z(n160) );
  XNOR U2931 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U2932 ( .A(n2965), .B(n2966), .Z(n163) );
  NANDN U2933 ( .A(n1922), .B(n2967), .Z(n2966) );
  OR U2934 ( .A(n1921), .B(n1919), .Z(n2967) );
  AND U2935 ( .A(n2968), .B(n2969), .Z(n1922) );
  NANDN U2936 ( .A(n2970), .B(n2971), .Z(n2969) );
  OR U2937 ( .A(n2972), .B(n40), .Z(n2971) );
  NAND U2938 ( .A(n40), .B(n2972), .Z(n2968) );
  NAND U2939 ( .A(n1919), .B(n1921), .Z(n2965) );
  ANDN U2940 ( .B(A[3]), .A(n42), .Z(n1921) );
  XOR U2941 ( .A(n2974), .B(n2975), .Z(n1919) );
  XNOR U2942 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2943 ( .A(B[0]), .B(A[12]), .Z(n2826) );
  XOR U2944 ( .A(n2836), .B(n2978), .Z(n2828) );
  XNOR U2945 ( .A(n2835), .B(n2833), .Z(n2978) );
  AND U2946 ( .A(n2979), .B(n2980), .Z(n2833) );
  NANDN U2947 ( .A(n2912), .B(n2981), .Z(n2980) );
  NANDN U2948 ( .A(n2911), .B(n5), .Z(n2981) );
  AND U2949 ( .A(n2982), .B(n2983), .Z(n2912) );
  NANDN U2950 ( .A(n2919), .B(n2984), .Z(n2983) );
  OR U2951 ( .A(n2918), .B(n2916), .Z(n2984) );
  AND U2952 ( .A(n2985), .B(n2986), .Z(n2919) );
  NANDN U2953 ( .A(n2927), .B(n2987), .Z(n2986) );
  NANDN U2954 ( .A(n2926), .B(n7), .Z(n2987) );
  AND U2955 ( .A(n2988), .B(n2989), .Z(n2927) );
  NANDN U2956 ( .A(n2934), .B(n2990), .Z(n2989) );
  OR U2957 ( .A(n2933), .B(n2931), .Z(n2990) );
  AND U2958 ( .A(n2991), .B(n2992), .Z(n2934) );
  NANDN U2959 ( .A(n2942), .B(n2993), .Z(n2992) );
  NANDN U2960 ( .A(n2941), .B(n9), .Z(n2993) );
  AND U2961 ( .A(n2994), .B(n2995), .Z(n2942) );
  NANDN U2962 ( .A(n2949), .B(n2996), .Z(n2995) );
  OR U2963 ( .A(n2948), .B(n2946), .Z(n2996) );
  AND U2964 ( .A(n2997), .B(n2998), .Z(n2949) );
  NANDN U2965 ( .A(n2957), .B(n2999), .Z(n2998) );
  NANDN U2966 ( .A(n2956), .B(n11), .Z(n2999) );
  AND U2967 ( .A(n3000), .B(n3001), .Z(n2957) );
  NANDN U2968 ( .A(n2964), .B(n3002), .Z(n3001) );
  OR U2969 ( .A(n2963), .B(n2961), .Z(n3002) );
  AND U2970 ( .A(n3003), .B(n3004), .Z(n2964) );
  NANDN U2971 ( .A(n2976), .B(n3005), .Z(n3004) );
  NAND U2972 ( .A(n2974), .B(n2977), .Z(n3005) );
  NANDN U2973 ( .A(n3006), .B(n3007), .Z(n2976) );
  AND U2974 ( .A(A[0]), .B(B[2]), .Z(n3007) );
  NANDN U2975 ( .A(n2977), .B(n30), .Z(n3003) );
  XNOR U2976 ( .A(n3008), .B(n3009), .Z(n2974) );
  NAND U2977 ( .A(A[0]), .B(B[3]), .Z(n3009) );
  NAND U2978 ( .A(B[1]), .B(A[2]), .Z(n2977) );
  NAND U2979 ( .A(n2961), .B(n2963), .Z(n3000) );
  ANDN U2980 ( .B(A[3]), .A(n41), .Z(n2963) );
  XOR U2981 ( .A(n3010), .B(n3011), .Z(n2961) );
  XNOR U2982 ( .A(n3012), .B(n3013), .Z(n3011) );
  NAND U2983 ( .A(n2954), .B(n2956), .Z(n2997) );
  ANDN U2984 ( .B(A[4]), .A(n41), .Z(n2956) );
  XOR U2985 ( .A(n3014), .B(n3015), .Z(n2954) );
  XNOR U2986 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U2987 ( .A(n2946), .B(n2948), .Z(n2994) );
  ANDN U2988 ( .B(A[5]), .A(n41), .Z(n2948) );
  XNOR U2989 ( .A(n3018), .B(n3019), .Z(n2946) );
  XNOR U2990 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND U2991 ( .A(n2939), .B(n2941), .Z(n2991) );
  ANDN U2992 ( .B(A[6]), .A(n41), .Z(n2941) );
  XOR U2993 ( .A(n3022), .B(n3023), .Z(n2939) );
  XNOR U2994 ( .A(n3024), .B(n3025), .Z(n3023) );
  NAND U2995 ( .A(n2931), .B(n2933), .Z(n2988) );
  ANDN U2996 ( .B(A[7]), .A(n41), .Z(n2933) );
  XNOR U2997 ( .A(n3026), .B(n3027), .Z(n2931) );
  XNOR U2998 ( .A(n3028), .B(n3029), .Z(n3027) );
  NAND U2999 ( .A(n2924), .B(n2926), .Z(n2985) );
  ANDN U3000 ( .B(A[8]), .A(n41), .Z(n2926) );
  XOR U3001 ( .A(n3030), .B(n3031), .Z(n2924) );
  XNOR U3002 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3003 ( .A(n2916), .B(n2918), .Z(n2982) );
  ANDN U3004 ( .B(A[9]), .A(n41), .Z(n2918) );
  XNOR U3005 ( .A(n3034), .B(n3035), .Z(n2916) );
  XNOR U3006 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3007 ( .A(n2909), .B(n2911), .Z(n2979) );
  ANDN U3008 ( .B(A[10]), .A(n41), .Z(n2911) );
  XOR U3009 ( .A(n3038), .B(n3039), .Z(n2909) );
  XNOR U3010 ( .A(n3040), .B(n3041), .Z(n3039) );
  ANDN U3011 ( .B(A[11]), .A(n41), .Z(n2835) );
  XNOR U3012 ( .A(n2843), .B(n3042), .Z(n2836) );
  XNOR U3013 ( .A(n2842), .B(n2840), .Z(n3042) );
  AND U3014 ( .A(n3043), .B(n3044), .Z(n2840) );
  NANDN U3015 ( .A(n3041), .B(n3045), .Z(n3044) );
  OR U3016 ( .A(n3040), .B(n3038), .Z(n3045) );
  AND U3017 ( .A(n3046), .B(n3047), .Z(n3041) );
  NANDN U3018 ( .A(n3037), .B(n3048), .Z(n3047) );
  NANDN U3019 ( .A(n3036), .B(n3034), .Z(n3048) );
  AND U3020 ( .A(n3049), .B(n3050), .Z(n3037) );
  NANDN U3021 ( .A(n3033), .B(n3051), .Z(n3050) );
  OR U3022 ( .A(n3032), .B(n3030), .Z(n3051) );
  AND U3023 ( .A(n3052), .B(n3053), .Z(n3033) );
  NANDN U3024 ( .A(n3029), .B(n3054), .Z(n3053) );
  NANDN U3025 ( .A(n3028), .B(n3026), .Z(n3054) );
  AND U3026 ( .A(n3055), .B(n3056), .Z(n3029) );
  NANDN U3027 ( .A(n3025), .B(n3057), .Z(n3056) );
  OR U3028 ( .A(n3024), .B(n3022), .Z(n3057) );
  AND U3029 ( .A(n3058), .B(n3059), .Z(n3025) );
  NANDN U3030 ( .A(n3021), .B(n3060), .Z(n3059) );
  NANDN U3031 ( .A(n3020), .B(n3018), .Z(n3060) );
  AND U3032 ( .A(n3061), .B(n3062), .Z(n3021) );
  NANDN U3033 ( .A(n3017), .B(n3063), .Z(n3062) );
  OR U3034 ( .A(n3016), .B(n3014), .Z(n3063) );
  AND U3035 ( .A(n3064), .B(n3065), .Z(n3017) );
  NANDN U3036 ( .A(n3012), .B(n3066), .Z(n3065) );
  NAND U3037 ( .A(n3010), .B(n3013), .Z(n3066) );
  NANDN U3038 ( .A(n3008), .B(n3067), .Z(n3012) );
  AND U3039 ( .A(A[0]), .B(B[3]), .Z(n3067) );
  NAND U3040 ( .A(B[2]), .B(A[1]), .Z(n3008) );
  NANDN U3041 ( .A(n3013), .B(n31), .Z(n3064) );
  XNOR U3042 ( .A(n3068), .B(n3069), .Z(n3010) );
  NAND U3043 ( .A(A[0]), .B(B[4]), .Z(n3069) );
  NAND U3044 ( .A(A[2]), .B(B[2]), .Z(n3013) );
  NAND U3045 ( .A(n3014), .B(n3016), .Z(n3061) );
  AND U3046 ( .A(A[3]), .B(B[2]), .Z(n3016) );
  XOR U3047 ( .A(n3070), .B(n3071), .Z(n3014) );
  XNOR U3048 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3049 ( .A(n3018), .B(n3020), .Z(n3058) );
  AND U3050 ( .A(A[4]), .B(B[2]), .Z(n3020) );
  XNOR U3051 ( .A(n3074), .B(n3075), .Z(n3018) );
  XNOR U3052 ( .A(n3076), .B(n3077), .Z(n3075) );
  NAND U3053 ( .A(n3022), .B(n3024), .Z(n3055) );
  AND U3054 ( .A(A[5]), .B(B[2]), .Z(n3024) );
  XNOR U3055 ( .A(n3078), .B(n3079), .Z(n3022) );
  XNOR U3056 ( .A(n3080), .B(n3081), .Z(n3079) );
  NANDN U3057 ( .A(n3026), .B(n3028), .Z(n3052) );
  AND U3058 ( .A(A[6]), .B(B[2]), .Z(n3028) );
  XNOR U3059 ( .A(n3082), .B(n3083), .Z(n3026) );
  XNOR U3060 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3061 ( .A(n3030), .B(n3032), .Z(n3049) );
  AND U3062 ( .A(A[7]), .B(B[2]), .Z(n3032) );
  XNOR U3063 ( .A(n3086), .B(n3087), .Z(n3030) );
  XNOR U3064 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3065 ( .A(n3034), .B(n3036), .Z(n3046) );
  AND U3066 ( .A(A[8]), .B(B[2]), .Z(n3036) );
  XNOR U3067 ( .A(n3090), .B(n3091), .Z(n3034) );
  XNOR U3068 ( .A(n3092), .B(n3093), .Z(n3091) );
  NAND U3069 ( .A(n3038), .B(n3040), .Z(n3043) );
  AND U3070 ( .A(A[9]), .B(B[2]), .Z(n3040) );
  XNOR U3071 ( .A(n3094), .B(n3095), .Z(n3038) );
  XNOR U3072 ( .A(n3096), .B(n3097), .Z(n3095) );
  AND U3073 ( .A(A[10]), .B(B[2]), .Z(n2842) );
  XNOR U3074 ( .A(n2850), .B(n3098), .Z(n2843) );
  XNOR U3075 ( .A(n2849), .B(n2847), .Z(n3098) );
  AND U3076 ( .A(n3099), .B(n3100), .Z(n2847) );
  NANDN U3077 ( .A(n3097), .B(n3101), .Z(n3100) );
  NANDN U3078 ( .A(n3096), .B(n3094), .Z(n3101) );
  AND U3079 ( .A(n3102), .B(n3103), .Z(n3097) );
  NANDN U3080 ( .A(n3093), .B(n3104), .Z(n3103) );
  OR U3081 ( .A(n3092), .B(n3090), .Z(n3104) );
  AND U3082 ( .A(n3105), .B(n3106), .Z(n3093) );
  NANDN U3083 ( .A(n3089), .B(n3107), .Z(n3106) );
  NANDN U3084 ( .A(n3088), .B(n3086), .Z(n3107) );
  AND U3085 ( .A(n3108), .B(n3109), .Z(n3089) );
  NANDN U3086 ( .A(n3085), .B(n3110), .Z(n3109) );
  OR U3087 ( .A(n3084), .B(n3082), .Z(n3110) );
  AND U3088 ( .A(n3111), .B(n3112), .Z(n3085) );
  NANDN U3089 ( .A(n3081), .B(n3113), .Z(n3112) );
  NANDN U3090 ( .A(n3080), .B(n3078), .Z(n3113) );
  AND U3091 ( .A(n3114), .B(n3115), .Z(n3081) );
  NANDN U3092 ( .A(n3077), .B(n3116), .Z(n3115) );
  OR U3093 ( .A(n3076), .B(n3074), .Z(n3116) );
  AND U3094 ( .A(n3117), .B(n3118), .Z(n3077) );
  NANDN U3095 ( .A(n3072), .B(n3119), .Z(n3118) );
  NAND U3096 ( .A(n3070), .B(n3073), .Z(n3119) );
  NANDN U3097 ( .A(n3068), .B(n3120), .Z(n3072) );
  AND U3098 ( .A(A[0]), .B(B[4]), .Z(n3120) );
  NAND U3099 ( .A(B[3]), .B(A[1]), .Z(n3068) );
  NANDN U3100 ( .A(n3073), .B(n32), .Z(n3117) );
  XNOR U3101 ( .A(n3121), .B(n3122), .Z(n3070) );
  NAND U3102 ( .A(A[0]), .B(B[5]), .Z(n3122) );
  NAND U3103 ( .A(A[2]), .B(B[3]), .Z(n3073) );
  NAND U3104 ( .A(n3074), .B(n3076), .Z(n3114) );
  AND U3105 ( .A(A[3]), .B(B[3]), .Z(n3076) );
  XOR U3106 ( .A(n3123), .B(n3124), .Z(n3074) );
  XNOR U3107 ( .A(n3125), .B(n3126), .Z(n3124) );
  NANDN U3108 ( .A(n3078), .B(n3080), .Z(n3111) );
  AND U3109 ( .A(A[4]), .B(B[3]), .Z(n3080) );
  XNOR U3110 ( .A(n3127), .B(n3128), .Z(n3078) );
  XNOR U3111 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND U3112 ( .A(n3082), .B(n3084), .Z(n3108) );
  AND U3113 ( .A(A[5]), .B(B[3]), .Z(n3084) );
  XNOR U3114 ( .A(n3131), .B(n3132), .Z(n3082) );
  XNOR U3115 ( .A(n3133), .B(n3134), .Z(n3132) );
  NANDN U3116 ( .A(n3086), .B(n3088), .Z(n3105) );
  AND U3117 ( .A(A[6]), .B(B[3]), .Z(n3088) );
  XNOR U3118 ( .A(n3135), .B(n3136), .Z(n3086) );
  XNOR U3119 ( .A(n3137), .B(n3138), .Z(n3136) );
  NAND U3120 ( .A(n3090), .B(n3092), .Z(n3102) );
  AND U3121 ( .A(A[7]), .B(B[3]), .Z(n3092) );
  XNOR U3122 ( .A(n3139), .B(n3140), .Z(n3090) );
  XNOR U3123 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U3124 ( .A(n3094), .B(n3096), .Z(n3099) );
  AND U3125 ( .A(A[8]), .B(B[3]), .Z(n3096) );
  XNOR U3126 ( .A(n3143), .B(n3144), .Z(n3094) );
  XNOR U3127 ( .A(n3145), .B(n3146), .Z(n3144) );
  AND U3128 ( .A(A[9]), .B(B[3]), .Z(n2849) );
  XNOR U3129 ( .A(n2857), .B(n3147), .Z(n2850) );
  XNOR U3130 ( .A(n2856), .B(n2854), .Z(n3147) );
  AND U3131 ( .A(n3148), .B(n3149), .Z(n2854) );
  NANDN U3132 ( .A(n3146), .B(n3150), .Z(n3149) );
  OR U3133 ( .A(n3145), .B(n3143), .Z(n3150) );
  AND U3134 ( .A(n3151), .B(n3152), .Z(n3146) );
  NANDN U3135 ( .A(n3142), .B(n3153), .Z(n3152) );
  NANDN U3136 ( .A(n3141), .B(n3139), .Z(n3153) );
  AND U3137 ( .A(n3154), .B(n3155), .Z(n3142) );
  NANDN U3138 ( .A(n3138), .B(n3156), .Z(n3155) );
  OR U3139 ( .A(n3137), .B(n3135), .Z(n3156) );
  AND U3140 ( .A(n3157), .B(n3158), .Z(n3138) );
  NANDN U3141 ( .A(n3134), .B(n3159), .Z(n3158) );
  NANDN U3142 ( .A(n3133), .B(n3131), .Z(n3159) );
  AND U3143 ( .A(n3160), .B(n3161), .Z(n3134) );
  NANDN U3144 ( .A(n3130), .B(n3162), .Z(n3161) );
  OR U3145 ( .A(n3129), .B(n3127), .Z(n3162) );
  AND U3146 ( .A(n3163), .B(n3164), .Z(n3130) );
  NANDN U3147 ( .A(n3125), .B(n3165), .Z(n3164) );
  NAND U3148 ( .A(n3123), .B(n3126), .Z(n3165) );
  NANDN U3149 ( .A(n3121), .B(n3166), .Z(n3125) );
  AND U3150 ( .A(A[0]), .B(B[5]), .Z(n3166) );
  NAND U3151 ( .A(B[4]), .B(A[1]), .Z(n3121) );
  NANDN U3152 ( .A(n3126), .B(n33), .Z(n3163) );
  XNOR U3153 ( .A(n3167), .B(n3168), .Z(n3123) );
  NAND U3154 ( .A(A[0]), .B(B[6]), .Z(n3168) );
  NAND U3155 ( .A(A[2]), .B(B[4]), .Z(n3126) );
  NAND U3156 ( .A(n3127), .B(n3129), .Z(n3160) );
  AND U3157 ( .A(A[3]), .B(B[4]), .Z(n3129) );
  XOR U3158 ( .A(n3169), .B(n3170), .Z(n3127) );
  XNOR U3159 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3160 ( .A(n3131), .B(n3133), .Z(n3157) );
  AND U3161 ( .A(A[4]), .B(B[4]), .Z(n3133) );
  XNOR U3162 ( .A(n3173), .B(n3174), .Z(n3131) );
  XNOR U3163 ( .A(n3175), .B(n3176), .Z(n3174) );
  NAND U3164 ( .A(n3135), .B(n3137), .Z(n3154) );
  AND U3165 ( .A(A[5]), .B(B[4]), .Z(n3137) );
  XNOR U3166 ( .A(n3177), .B(n3178), .Z(n3135) );
  XNOR U3167 ( .A(n3179), .B(n3180), .Z(n3178) );
  NANDN U3168 ( .A(n3139), .B(n3141), .Z(n3151) );
  AND U3169 ( .A(A[6]), .B(B[4]), .Z(n3141) );
  XNOR U3170 ( .A(n3181), .B(n3182), .Z(n3139) );
  XNOR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3143), .B(n3145), .Z(n3148) );
  AND U3173 ( .A(A[7]), .B(B[4]), .Z(n3145) );
  XNOR U3174 ( .A(n3185), .B(n3186), .Z(n3143) );
  XNOR U3175 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3176 ( .A(A[8]), .B(B[4]), .Z(n2856) );
  XNOR U3177 ( .A(n2864), .B(n3189), .Z(n2857) );
  XNOR U3178 ( .A(n2863), .B(n2861), .Z(n3189) );
  AND U3179 ( .A(n3190), .B(n3191), .Z(n2861) );
  NANDN U3180 ( .A(n3188), .B(n3192), .Z(n3191) );
  NANDN U3181 ( .A(n3187), .B(n3185), .Z(n3192) );
  AND U3182 ( .A(n3193), .B(n3194), .Z(n3188) );
  NANDN U3183 ( .A(n3184), .B(n3195), .Z(n3194) );
  OR U3184 ( .A(n3183), .B(n3181), .Z(n3195) );
  AND U3185 ( .A(n3196), .B(n3197), .Z(n3184) );
  NANDN U3186 ( .A(n3180), .B(n3198), .Z(n3197) );
  NANDN U3187 ( .A(n3179), .B(n3177), .Z(n3198) );
  AND U3188 ( .A(n3199), .B(n3200), .Z(n3180) );
  NANDN U3189 ( .A(n3176), .B(n3201), .Z(n3200) );
  OR U3190 ( .A(n3175), .B(n3173), .Z(n3201) );
  AND U3191 ( .A(n3202), .B(n3203), .Z(n3176) );
  NANDN U3192 ( .A(n3171), .B(n3204), .Z(n3203) );
  NAND U3193 ( .A(n3169), .B(n3172), .Z(n3204) );
  NANDN U3194 ( .A(n3167), .B(n3205), .Z(n3171) );
  AND U3195 ( .A(A[0]), .B(B[6]), .Z(n3205) );
  NAND U3196 ( .A(B[5]), .B(A[1]), .Z(n3167) );
  NANDN U3197 ( .A(n3172), .B(n34), .Z(n3202) );
  XNOR U3198 ( .A(n3206), .B(n3207), .Z(n3169) );
  NAND U3199 ( .A(A[0]), .B(B[7]), .Z(n3207) );
  NAND U3200 ( .A(A[2]), .B(B[5]), .Z(n3172) );
  NAND U3201 ( .A(n3173), .B(n3175), .Z(n3199) );
  AND U3202 ( .A(A[3]), .B(B[5]), .Z(n3175) );
  XOR U3203 ( .A(n3208), .B(n3209), .Z(n3173) );
  XNOR U3204 ( .A(n3210), .B(n3211), .Z(n3209) );
  NANDN U3205 ( .A(n3177), .B(n3179), .Z(n3196) );
  AND U3206 ( .A(A[4]), .B(B[5]), .Z(n3179) );
  XNOR U3207 ( .A(n3212), .B(n3213), .Z(n3177) );
  XNOR U3208 ( .A(n3214), .B(n3215), .Z(n3213) );
  NAND U3209 ( .A(n3181), .B(n3183), .Z(n3193) );
  AND U3210 ( .A(A[5]), .B(B[5]), .Z(n3183) );
  XNOR U3211 ( .A(n3216), .B(n3217), .Z(n3181) );
  XNOR U3212 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3213 ( .A(n3185), .B(n3187), .Z(n3190) );
  AND U3214 ( .A(A[6]), .B(B[5]), .Z(n3187) );
  XNOR U3215 ( .A(n3220), .B(n3221), .Z(n3185) );
  XNOR U3216 ( .A(n3222), .B(n3223), .Z(n3221) );
  AND U3217 ( .A(A[7]), .B(B[5]), .Z(n2863) );
  XNOR U3218 ( .A(n2871), .B(n3224), .Z(n2864) );
  XNOR U3219 ( .A(n2870), .B(n2868), .Z(n3224) );
  AND U3220 ( .A(n3225), .B(n3226), .Z(n2868) );
  NANDN U3221 ( .A(n3223), .B(n3227), .Z(n3226) );
  OR U3222 ( .A(n3222), .B(n3220), .Z(n3227) );
  AND U3223 ( .A(n3228), .B(n3229), .Z(n3223) );
  NANDN U3224 ( .A(n3219), .B(n3230), .Z(n3229) );
  NANDN U3225 ( .A(n3218), .B(n3216), .Z(n3230) );
  AND U3226 ( .A(n3231), .B(n3232), .Z(n3219) );
  NANDN U3227 ( .A(n3215), .B(n3233), .Z(n3232) );
  OR U3228 ( .A(n3214), .B(n3212), .Z(n3233) );
  AND U3229 ( .A(n3234), .B(n3235), .Z(n3215) );
  NANDN U3230 ( .A(n3210), .B(n3236), .Z(n3235) );
  NAND U3231 ( .A(n3208), .B(n3211), .Z(n3236) );
  NANDN U3232 ( .A(n3206), .B(n3237), .Z(n3210) );
  AND U3233 ( .A(A[0]), .B(B[7]), .Z(n3237) );
  NAND U3234 ( .A(B[6]), .B(A[1]), .Z(n3206) );
  NANDN U3235 ( .A(n3211), .B(n35), .Z(n3234) );
  XNOR U3236 ( .A(n3238), .B(n3239), .Z(n3208) );
  NAND U3237 ( .A(A[0]), .B(B[8]), .Z(n3239) );
  NAND U3238 ( .A(A[2]), .B(B[6]), .Z(n3211) );
  NAND U3239 ( .A(n3212), .B(n3214), .Z(n3231) );
  AND U3240 ( .A(A[3]), .B(B[6]), .Z(n3214) );
  XOR U3241 ( .A(n3240), .B(n3241), .Z(n3212) );
  XNOR U3242 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3243 ( .A(n3216), .B(n3218), .Z(n3228) );
  AND U3244 ( .A(A[4]), .B(B[6]), .Z(n3218) );
  XNOR U3245 ( .A(n3244), .B(n3245), .Z(n3216) );
  XNOR U3246 ( .A(n3246), .B(n3247), .Z(n3245) );
  NAND U3247 ( .A(n3220), .B(n3222), .Z(n3225) );
  AND U3248 ( .A(A[5]), .B(B[6]), .Z(n3222) );
  XNOR U3249 ( .A(n3248), .B(n3249), .Z(n3220) );
  XNOR U3250 ( .A(n3250), .B(n3251), .Z(n3249) );
  AND U3251 ( .A(A[6]), .B(B[6]), .Z(n2870) );
  XNOR U3252 ( .A(n2878), .B(n3252), .Z(n2871) );
  XNOR U3253 ( .A(n2877), .B(n2875), .Z(n3252) );
  AND U3254 ( .A(n3253), .B(n3254), .Z(n2875) );
  NANDN U3255 ( .A(n3251), .B(n3255), .Z(n3254) );
  NANDN U3256 ( .A(n3250), .B(n3248), .Z(n3255) );
  AND U3257 ( .A(n3256), .B(n3257), .Z(n3251) );
  NANDN U3258 ( .A(n3247), .B(n3258), .Z(n3257) );
  OR U3259 ( .A(n3246), .B(n3244), .Z(n3258) );
  AND U3260 ( .A(n3259), .B(n3260), .Z(n3247) );
  NANDN U3261 ( .A(n3242), .B(n3261), .Z(n3260) );
  NAND U3262 ( .A(n3240), .B(n3243), .Z(n3261) );
  NANDN U3263 ( .A(n3238), .B(n3262), .Z(n3242) );
  AND U3264 ( .A(A[0]), .B(B[8]), .Z(n3262) );
  NAND U3265 ( .A(B[7]), .B(A[1]), .Z(n3238) );
  NANDN U3266 ( .A(n3243), .B(n36), .Z(n3259) );
  XNOR U3267 ( .A(n3263), .B(n3264), .Z(n3240) );
  NAND U3268 ( .A(A[0]), .B(B[9]), .Z(n3264) );
  NAND U3269 ( .A(A[2]), .B(B[7]), .Z(n3243) );
  NAND U3270 ( .A(n3244), .B(n3246), .Z(n3256) );
  AND U3271 ( .A(A[3]), .B(B[7]), .Z(n3246) );
  XOR U3272 ( .A(n3265), .B(n3266), .Z(n3244) );
  XNOR U3273 ( .A(n3267), .B(n3268), .Z(n3266) );
  NANDN U3274 ( .A(n3248), .B(n3250), .Z(n3253) );
  AND U3275 ( .A(A[4]), .B(B[7]), .Z(n3250) );
  XNOR U3276 ( .A(n3269), .B(n3270), .Z(n3248) );
  XNOR U3277 ( .A(n3271), .B(n3272), .Z(n3270) );
  AND U3278 ( .A(A[5]), .B(B[7]), .Z(n2877) );
  XNOR U3279 ( .A(n2885), .B(n3273), .Z(n2878) );
  XNOR U3280 ( .A(n2884), .B(n2882), .Z(n3273) );
  AND U3281 ( .A(n3274), .B(n3275), .Z(n2882) );
  NANDN U3282 ( .A(n3272), .B(n3276), .Z(n3275) );
  OR U3283 ( .A(n3271), .B(n3269), .Z(n3276) );
  AND U3284 ( .A(n3277), .B(n3278), .Z(n3272) );
  NANDN U3285 ( .A(n3267), .B(n3279), .Z(n3278) );
  NAND U3286 ( .A(n3265), .B(n3268), .Z(n3279) );
  NANDN U3287 ( .A(n3263), .B(n3280), .Z(n3267) );
  AND U3288 ( .A(A[0]), .B(B[9]), .Z(n3280) );
  NAND U3289 ( .A(B[8]), .B(A[1]), .Z(n3263) );
  NANDN U3290 ( .A(n3268), .B(n37), .Z(n3277) );
  XNOR U3291 ( .A(n3281), .B(n3282), .Z(n3265) );
  NAND U3292 ( .A(A[0]), .B(B[10]), .Z(n3282) );
  NAND U3293 ( .A(A[2]), .B(B[8]), .Z(n3268) );
  NAND U3294 ( .A(n3269), .B(n3271), .Z(n3274) );
  AND U3295 ( .A(A[3]), .B(B[8]), .Z(n3271) );
  XOR U3296 ( .A(n3283), .B(n3284), .Z(n3269) );
  XNOR U3297 ( .A(n3285), .B(n3286), .Z(n3284) );
  AND U3298 ( .A(A[4]), .B(B[8]), .Z(n2884) );
  XNOR U3299 ( .A(n2892), .B(n3287), .Z(n2885) );
  XNOR U3300 ( .A(n2891), .B(n2889), .Z(n3287) );
  AND U3301 ( .A(n3288), .B(n3289), .Z(n2889) );
  NANDN U3302 ( .A(n3285), .B(n3290), .Z(n3289) );
  NAND U3303 ( .A(n3283), .B(n3286), .Z(n3290) );
  NANDN U3304 ( .A(n3281), .B(n3291), .Z(n3285) );
  AND U3305 ( .A(A[0]), .B(B[10]), .Z(n3291) );
  NAND U3306 ( .A(B[9]), .B(A[1]), .Z(n3281) );
  NANDN U3307 ( .A(n3286), .B(n38), .Z(n3288) );
  XNOR U3308 ( .A(n3292), .B(n3293), .Z(n3283) );
  NAND U3309 ( .A(A[0]), .B(B[11]), .Z(n3293) );
  NAND U3310 ( .A(A[2]), .B(B[9]), .Z(n3286) );
  AND U3311 ( .A(A[3]), .B(B[9]), .Z(n2891) );
  XOR U3312 ( .A(n2898), .B(n3294), .Z(n2892) );
  XNOR U3313 ( .A(n2896), .B(n2899), .Z(n3294) );
  NAND U3314 ( .A(A[2]), .B(B[10]), .Z(n2899) );
  NANDN U3315 ( .A(n3292), .B(n3295), .Z(n2896) );
  AND U3316 ( .A(A[0]), .B(B[11]), .Z(n3295) );
  NAND U3317 ( .A(B[10]), .B(A[1]), .Z(n3292) );
  XNOR U3318 ( .A(n2901), .B(n3296), .Z(n2898) );
  NAND U3319 ( .A(A[0]), .B(B[12]), .Z(n3296) );
  NAND U3320 ( .A(B[11]), .B(A[1]), .Z(n2901) );
  XNOR U3321 ( .A(n2973), .B(n3297), .Z(PRODUCT[2]) );
  XNOR U3322 ( .A(n2970), .B(n2972), .Z(n3297) );
  ANDN U3323 ( .B(n44), .A(n43), .Z(n2972) );
  NAND U3324 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U3325 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U3326 ( .A(B[0]), .B(A[2]), .Z(n2970) );
  XNOR U3327 ( .A(n3006), .B(n3298), .Z(n2973) );
  NAND U3328 ( .A(A[0]), .B(B[2]), .Z(n3298) );
  NAND U3329 ( .A(B[1]), .B(A[1]), .Z(n3006) );
endmodule


module matrixMult_N_M_1_N16_M32 ( clk, rst, x, y, o );
  input [511:0] x;
  input [8191:0] y;
  output [511:0] o;
  input clk, rst;
  wire   N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507,
         N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617,
         N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650,
         N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661,
         N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672,
         N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683,
         N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694,
         N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705,
         N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716,
         N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727,
         N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782,
         N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793,
         N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815,
         N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826,
         N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859,
         N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892,
         N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903,
         N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936,
         N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947,
         N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969,
         N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980,
         N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991,
         N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002,
         N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012,
         N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022,
         N1023, N1024;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511;

  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[3][0]  ( .D(N225), .CLK(clk), .RST(rst), .Q(o[96]) );
  DFF \oi_reg[3][1]  ( .D(N226), .CLK(clk), .RST(rst), .Q(o[97]) );
  DFF \oi_reg[3][2]  ( .D(N227), .CLK(clk), .RST(rst), .Q(o[98]) );
  DFF \oi_reg[3][3]  ( .D(N228), .CLK(clk), .RST(rst), .Q(o[99]) );
  DFF \oi_reg[3][4]  ( .D(N229), .CLK(clk), .RST(rst), .Q(o[100]) );
  DFF \oi_reg[3][5]  ( .D(N230), .CLK(clk), .RST(rst), .Q(o[101]) );
  DFF \oi_reg[3][6]  ( .D(N231), .CLK(clk), .RST(rst), .Q(o[102]) );
  DFF \oi_reg[3][7]  ( .D(N232), .CLK(clk), .RST(rst), .Q(o[103]) );
  DFF \oi_reg[3][8]  ( .D(N233), .CLK(clk), .RST(rst), .Q(o[104]) );
  DFF \oi_reg[3][9]  ( .D(N234), .CLK(clk), .RST(rst), .Q(o[105]) );
  DFF \oi_reg[3][10]  ( .D(N235), .CLK(clk), .RST(rst), .Q(o[106]) );
  DFF \oi_reg[3][11]  ( .D(N236), .CLK(clk), .RST(rst), .Q(o[107]) );
  DFF \oi_reg[3][12]  ( .D(N237), .CLK(clk), .RST(rst), .Q(o[108]) );
  DFF \oi_reg[3][13]  ( .D(N238), .CLK(clk), .RST(rst), .Q(o[109]) );
  DFF \oi_reg[3][14]  ( .D(N239), .CLK(clk), .RST(rst), .Q(o[110]) );
  DFF \oi_reg[3][15]  ( .D(N240), .CLK(clk), .RST(rst), .Q(o[111]) );
  DFF \oi_reg[3][16]  ( .D(N241), .CLK(clk), .RST(rst), .Q(o[112]) );
  DFF \oi_reg[3][17]  ( .D(N242), .CLK(clk), .RST(rst), .Q(o[113]) );
  DFF \oi_reg[3][18]  ( .D(N243), .CLK(clk), .RST(rst), .Q(o[114]) );
  DFF \oi_reg[3][19]  ( .D(N244), .CLK(clk), .RST(rst), .Q(o[115]) );
  DFF \oi_reg[3][20]  ( .D(N245), .CLK(clk), .RST(rst), .Q(o[116]) );
  DFF \oi_reg[3][21]  ( .D(N246), .CLK(clk), .RST(rst), .Q(o[117]) );
  DFF \oi_reg[3][22]  ( .D(N247), .CLK(clk), .RST(rst), .Q(o[118]) );
  DFF \oi_reg[3][23]  ( .D(N248), .CLK(clk), .RST(rst), .Q(o[119]) );
  DFF \oi_reg[3][24]  ( .D(N249), .CLK(clk), .RST(rst), .Q(o[120]) );
  DFF \oi_reg[3][25]  ( .D(N250), .CLK(clk), .RST(rst), .Q(o[121]) );
  DFF \oi_reg[3][26]  ( .D(N251), .CLK(clk), .RST(rst), .Q(o[122]) );
  DFF \oi_reg[3][27]  ( .D(N252), .CLK(clk), .RST(rst), .Q(o[123]) );
  DFF \oi_reg[3][28]  ( .D(N253), .CLK(clk), .RST(rst), .Q(o[124]) );
  DFF \oi_reg[3][29]  ( .D(N254), .CLK(clk), .RST(rst), .Q(o[125]) );
  DFF \oi_reg[3][30]  ( .D(N255), .CLK(clk), .RST(rst), .Q(o[126]) );
  DFF \oi_reg[3][31]  ( .D(N256), .CLK(clk), .RST(rst), .Q(o[127]) );
  DFF \oi_reg[4][0]  ( .D(N289), .CLK(clk), .RST(rst), .Q(o[128]) );
  DFF \oi_reg[4][1]  ( .D(N290), .CLK(clk), .RST(rst), .Q(o[129]) );
  DFF \oi_reg[4][2]  ( .D(N291), .CLK(clk), .RST(rst), .Q(o[130]) );
  DFF \oi_reg[4][3]  ( .D(N292), .CLK(clk), .RST(rst), .Q(o[131]) );
  DFF \oi_reg[4][4]  ( .D(N293), .CLK(clk), .RST(rst), .Q(o[132]) );
  DFF \oi_reg[4][5]  ( .D(N294), .CLK(clk), .RST(rst), .Q(o[133]) );
  DFF \oi_reg[4][6]  ( .D(N295), .CLK(clk), .RST(rst), .Q(o[134]) );
  DFF \oi_reg[4][7]  ( .D(N296), .CLK(clk), .RST(rst), .Q(o[135]) );
  DFF \oi_reg[4][8]  ( .D(N297), .CLK(clk), .RST(rst), .Q(o[136]) );
  DFF \oi_reg[4][9]  ( .D(N298), .CLK(clk), .RST(rst), .Q(o[137]) );
  DFF \oi_reg[4][10]  ( .D(N299), .CLK(clk), .RST(rst), .Q(o[138]) );
  DFF \oi_reg[4][11]  ( .D(N300), .CLK(clk), .RST(rst), .Q(o[139]) );
  DFF \oi_reg[4][12]  ( .D(N301), .CLK(clk), .RST(rst), .Q(o[140]) );
  DFF \oi_reg[4][13]  ( .D(N302), .CLK(clk), .RST(rst), .Q(o[141]) );
  DFF \oi_reg[4][14]  ( .D(N303), .CLK(clk), .RST(rst), .Q(o[142]) );
  DFF \oi_reg[4][15]  ( .D(N304), .CLK(clk), .RST(rst), .Q(o[143]) );
  DFF \oi_reg[4][16]  ( .D(N305), .CLK(clk), .RST(rst), .Q(o[144]) );
  DFF \oi_reg[4][17]  ( .D(N306), .CLK(clk), .RST(rst), .Q(o[145]) );
  DFF \oi_reg[4][18]  ( .D(N307), .CLK(clk), .RST(rst), .Q(o[146]) );
  DFF \oi_reg[4][19]  ( .D(N308), .CLK(clk), .RST(rst), .Q(o[147]) );
  DFF \oi_reg[4][20]  ( .D(N309), .CLK(clk), .RST(rst), .Q(o[148]) );
  DFF \oi_reg[4][21]  ( .D(N310), .CLK(clk), .RST(rst), .Q(o[149]) );
  DFF \oi_reg[4][22]  ( .D(N311), .CLK(clk), .RST(rst), .Q(o[150]) );
  DFF \oi_reg[4][23]  ( .D(N312), .CLK(clk), .RST(rst), .Q(o[151]) );
  DFF \oi_reg[4][24]  ( .D(N313), .CLK(clk), .RST(rst), .Q(o[152]) );
  DFF \oi_reg[4][25]  ( .D(N314), .CLK(clk), .RST(rst), .Q(o[153]) );
  DFF \oi_reg[4][26]  ( .D(N315), .CLK(clk), .RST(rst), .Q(o[154]) );
  DFF \oi_reg[4][27]  ( .D(N316), .CLK(clk), .RST(rst), .Q(o[155]) );
  DFF \oi_reg[4][28]  ( .D(N317), .CLK(clk), .RST(rst), .Q(o[156]) );
  DFF \oi_reg[4][29]  ( .D(N318), .CLK(clk), .RST(rst), .Q(o[157]) );
  DFF \oi_reg[4][30]  ( .D(N319), .CLK(clk), .RST(rst), .Q(o[158]) );
  DFF \oi_reg[4][31]  ( .D(N320), .CLK(clk), .RST(rst), .Q(o[159]) );
  DFF \oi_reg[5][0]  ( .D(N353), .CLK(clk), .RST(rst), .Q(o[160]) );
  DFF \oi_reg[5][1]  ( .D(N354), .CLK(clk), .RST(rst), .Q(o[161]) );
  DFF \oi_reg[5][2]  ( .D(N355), .CLK(clk), .RST(rst), .Q(o[162]) );
  DFF \oi_reg[5][3]  ( .D(N356), .CLK(clk), .RST(rst), .Q(o[163]) );
  DFF \oi_reg[5][4]  ( .D(N357), .CLK(clk), .RST(rst), .Q(o[164]) );
  DFF \oi_reg[5][5]  ( .D(N358), .CLK(clk), .RST(rst), .Q(o[165]) );
  DFF \oi_reg[5][6]  ( .D(N359), .CLK(clk), .RST(rst), .Q(o[166]) );
  DFF \oi_reg[5][7]  ( .D(N360), .CLK(clk), .RST(rst), .Q(o[167]) );
  DFF \oi_reg[5][8]  ( .D(N361), .CLK(clk), .RST(rst), .Q(o[168]) );
  DFF \oi_reg[5][9]  ( .D(N362), .CLK(clk), .RST(rst), .Q(o[169]) );
  DFF \oi_reg[5][10]  ( .D(N363), .CLK(clk), .RST(rst), .Q(o[170]) );
  DFF \oi_reg[5][11]  ( .D(N364), .CLK(clk), .RST(rst), .Q(o[171]) );
  DFF \oi_reg[5][12]  ( .D(N365), .CLK(clk), .RST(rst), .Q(o[172]) );
  DFF \oi_reg[5][13]  ( .D(N366), .CLK(clk), .RST(rst), .Q(o[173]) );
  DFF \oi_reg[5][14]  ( .D(N367), .CLK(clk), .RST(rst), .Q(o[174]) );
  DFF \oi_reg[5][15]  ( .D(N368), .CLK(clk), .RST(rst), .Q(o[175]) );
  DFF \oi_reg[5][16]  ( .D(N369), .CLK(clk), .RST(rst), .Q(o[176]) );
  DFF \oi_reg[5][17]  ( .D(N370), .CLK(clk), .RST(rst), .Q(o[177]) );
  DFF \oi_reg[5][18]  ( .D(N371), .CLK(clk), .RST(rst), .Q(o[178]) );
  DFF \oi_reg[5][19]  ( .D(N372), .CLK(clk), .RST(rst), .Q(o[179]) );
  DFF \oi_reg[5][20]  ( .D(N373), .CLK(clk), .RST(rst), .Q(o[180]) );
  DFF \oi_reg[5][21]  ( .D(N374), .CLK(clk), .RST(rst), .Q(o[181]) );
  DFF \oi_reg[5][22]  ( .D(N375), .CLK(clk), .RST(rst), .Q(o[182]) );
  DFF \oi_reg[5][23]  ( .D(N376), .CLK(clk), .RST(rst), .Q(o[183]) );
  DFF \oi_reg[5][24]  ( .D(N377), .CLK(clk), .RST(rst), .Q(o[184]) );
  DFF \oi_reg[5][25]  ( .D(N378), .CLK(clk), .RST(rst), .Q(o[185]) );
  DFF \oi_reg[5][26]  ( .D(N379), .CLK(clk), .RST(rst), .Q(o[186]) );
  DFF \oi_reg[5][27]  ( .D(N380), .CLK(clk), .RST(rst), .Q(o[187]) );
  DFF \oi_reg[5][28]  ( .D(N381), .CLK(clk), .RST(rst), .Q(o[188]) );
  DFF \oi_reg[5][29]  ( .D(N382), .CLK(clk), .RST(rst), .Q(o[189]) );
  DFF \oi_reg[5][30]  ( .D(N383), .CLK(clk), .RST(rst), .Q(o[190]) );
  DFF \oi_reg[5][31]  ( .D(N384), .CLK(clk), .RST(rst), .Q(o[191]) );
  DFF \oi_reg[6][0]  ( .D(N417), .CLK(clk), .RST(rst), .Q(o[192]) );
  DFF \oi_reg[6][1]  ( .D(N418), .CLK(clk), .RST(rst), .Q(o[193]) );
  DFF \oi_reg[6][2]  ( .D(N419), .CLK(clk), .RST(rst), .Q(o[194]) );
  DFF \oi_reg[6][3]  ( .D(N420), .CLK(clk), .RST(rst), .Q(o[195]) );
  DFF \oi_reg[6][4]  ( .D(N421), .CLK(clk), .RST(rst), .Q(o[196]) );
  DFF \oi_reg[6][5]  ( .D(N422), .CLK(clk), .RST(rst), .Q(o[197]) );
  DFF \oi_reg[6][6]  ( .D(N423), .CLK(clk), .RST(rst), .Q(o[198]) );
  DFF \oi_reg[6][7]  ( .D(N424), .CLK(clk), .RST(rst), .Q(o[199]) );
  DFF \oi_reg[6][8]  ( .D(N425), .CLK(clk), .RST(rst), .Q(o[200]) );
  DFF \oi_reg[6][9]  ( .D(N426), .CLK(clk), .RST(rst), .Q(o[201]) );
  DFF \oi_reg[6][10]  ( .D(N427), .CLK(clk), .RST(rst), .Q(o[202]) );
  DFF \oi_reg[6][11]  ( .D(N428), .CLK(clk), .RST(rst), .Q(o[203]) );
  DFF \oi_reg[6][12]  ( .D(N429), .CLK(clk), .RST(rst), .Q(o[204]) );
  DFF \oi_reg[6][13]  ( .D(N430), .CLK(clk), .RST(rst), .Q(o[205]) );
  DFF \oi_reg[6][14]  ( .D(N431), .CLK(clk), .RST(rst), .Q(o[206]) );
  DFF \oi_reg[6][15]  ( .D(N432), .CLK(clk), .RST(rst), .Q(o[207]) );
  DFF \oi_reg[6][16]  ( .D(N433), .CLK(clk), .RST(rst), .Q(o[208]) );
  DFF \oi_reg[6][17]  ( .D(N434), .CLK(clk), .RST(rst), .Q(o[209]) );
  DFF \oi_reg[6][18]  ( .D(N435), .CLK(clk), .RST(rst), .Q(o[210]) );
  DFF \oi_reg[6][19]  ( .D(N436), .CLK(clk), .RST(rst), .Q(o[211]) );
  DFF \oi_reg[6][20]  ( .D(N437), .CLK(clk), .RST(rst), .Q(o[212]) );
  DFF \oi_reg[6][21]  ( .D(N438), .CLK(clk), .RST(rst), .Q(o[213]) );
  DFF \oi_reg[6][22]  ( .D(N439), .CLK(clk), .RST(rst), .Q(o[214]) );
  DFF \oi_reg[6][23]  ( .D(N440), .CLK(clk), .RST(rst), .Q(o[215]) );
  DFF \oi_reg[6][24]  ( .D(N441), .CLK(clk), .RST(rst), .Q(o[216]) );
  DFF \oi_reg[6][25]  ( .D(N442), .CLK(clk), .RST(rst), .Q(o[217]) );
  DFF \oi_reg[6][26]  ( .D(N443), .CLK(clk), .RST(rst), .Q(o[218]) );
  DFF \oi_reg[6][27]  ( .D(N444), .CLK(clk), .RST(rst), .Q(o[219]) );
  DFF \oi_reg[6][28]  ( .D(N445), .CLK(clk), .RST(rst), .Q(o[220]) );
  DFF \oi_reg[6][29]  ( .D(N446), .CLK(clk), .RST(rst), .Q(o[221]) );
  DFF \oi_reg[6][30]  ( .D(N447), .CLK(clk), .RST(rst), .Q(o[222]) );
  DFF \oi_reg[6][31]  ( .D(N448), .CLK(clk), .RST(rst), .Q(o[223]) );
  DFF \oi_reg[7][0]  ( .D(N481), .CLK(clk), .RST(rst), .Q(o[224]) );
  DFF \oi_reg[7][1]  ( .D(N482), .CLK(clk), .RST(rst), .Q(o[225]) );
  DFF \oi_reg[7][2]  ( .D(N483), .CLK(clk), .RST(rst), .Q(o[226]) );
  DFF \oi_reg[7][3]  ( .D(N484), .CLK(clk), .RST(rst), .Q(o[227]) );
  DFF \oi_reg[7][4]  ( .D(N485), .CLK(clk), .RST(rst), .Q(o[228]) );
  DFF \oi_reg[7][5]  ( .D(N486), .CLK(clk), .RST(rst), .Q(o[229]) );
  DFF \oi_reg[7][6]  ( .D(N487), .CLK(clk), .RST(rst), .Q(o[230]) );
  DFF \oi_reg[7][7]  ( .D(N488), .CLK(clk), .RST(rst), .Q(o[231]) );
  DFF \oi_reg[7][8]  ( .D(N489), .CLK(clk), .RST(rst), .Q(o[232]) );
  DFF \oi_reg[7][9]  ( .D(N490), .CLK(clk), .RST(rst), .Q(o[233]) );
  DFF \oi_reg[7][10]  ( .D(N491), .CLK(clk), .RST(rst), .Q(o[234]) );
  DFF \oi_reg[7][11]  ( .D(N492), .CLK(clk), .RST(rst), .Q(o[235]) );
  DFF \oi_reg[7][12]  ( .D(N493), .CLK(clk), .RST(rst), .Q(o[236]) );
  DFF \oi_reg[7][13]  ( .D(N494), .CLK(clk), .RST(rst), .Q(o[237]) );
  DFF \oi_reg[7][14]  ( .D(N495), .CLK(clk), .RST(rst), .Q(o[238]) );
  DFF \oi_reg[7][15]  ( .D(N496), .CLK(clk), .RST(rst), .Q(o[239]) );
  DFF \oi_reg[7][16]  ( .D(N497), .CLK(clk), .RST(rst), .Q(o[240]) );
  DFF \oi_reg[7][17]  ( .D(N498), .CLK(clk), .RST(rst), .Q(o[241]) );
  DFF \oi_reg[7][18]  ( .D(N499), .CLK(clk), .RST(rst), .Q(o[242]) );
  DFF \oi_reg[7][19]  ( .D(N500), .CLK(clk), .RST(rst), .Q(o[243]) );
  DFF \oi_reg[7][20]  ( .D(N501), .CLK(clk), .RST(rst), .Q(o[244]) );
  DFF \oi_reg[7][21]  ( .D(N502), .CLK(clk), .RST(rst), .Q(o[245]) );
  DFF \oi_reg[7][22]  ( .D(N503), .CLK(clk), .RST(rst), .Q(o[246]) );
  DFF \oi_reg[7][23]  ( .D(N504), .CLK(clk), .RST(rst), .Q(o[247]) );
  DFF \oi_reg[7][24]  ( .D(N505), .CLK(clk), .RST(rst), .Q(o[248]) );
  DFF \oi_reg[7][25]  ( .D(N506), .CLK(clk), .RST(rst), .Q(o[249]) );
  DFF \oi_reg[7][26]  ( .D(N507), .CLK(clk), .RST(rst), .Q(o[250]) );
  DFF \oi_reg[7][27]  ( .D(N508), .CLK(clk), .RST(rst), .Q(o[251]) );
  DFF \oi_reg[7][28]  ( .D(N509), .CLK(clk), .RST(rst), .Q(o[252]) );
  DFF \oi_reg[7][29]  ( .D(N510), .CLK(clk), .RST(rst), .Q(o[253]) );
  DFF \oi_reg[7][30]  ( .D(N511), .CLK(clk), .RST(rst), .Q(o[254]) );
  DFF \oi_reg[7][31]  ( .D(N512), .CLK(clk), .RST(rst), .Q(o[255]) );
  DFF \oi_reg[8][0]  ( .D(N545), .CLK(clk), .RST(rst), .Q(o[256]) );
  DFF \oi_reg[8][1]  ( .D(N546), .CLK(clk), .RST(rst), .Q(o[257]) );
  DFF \oi_reg[8][2]  ( .D(N547), .CLK(clk), .RST(rst), .Q(o[258]) );
  DFF \oi_reg[8][3]  ( .D(N548), .CLK(clk), .RST(rst), .Q(o[259]) );
  DFF \oi_reg[8][4]  ( .D(N549), .CLK(clk), .RST(rst), .Q(o[260]) );
  DFF \oi_reg[8][5]  ( .D(N550), .CLK(clk), .RST(rst), .Q(o[261]) );
  DFF \oi_reg[8][6]  ( .D(N551), .CLK(clk), .RST(rst), .Q(o[262]) );
  DFF \oi_reg[8][7]  ( .D(N552), .CLK(clk), .RST(rst), .Q(o[263]) );
  DFF \oi_reg[8][8]  ( .D(N553), .CLK(clk), .RST(rst), .Q(o[264]) );
  DFF \oi_reg[8][9]  ( .D(N554), .CLK(clk), .RST(rst), .Q(o[265]) );
  DFF \oi_reg[8][10]  ( .D(N555), .CLK(clk), .RST(rst), .Q(o[266]) );
  DFF \oi_reg[8][11]  ( .D(N556), .CLK(clk), .RST(rst), .Q(o[267]) );
  DFF \oi_reg[8][12]  ( .D(N557), .CLK(clk), .RST(rst), .Q(o[268]) );
  DFF \oi_reg[8][13]  ( .D(N558), .CLK(clk), .RST(rst), .Q(o[269]) );
  DFF \oi_reg[8][14]  ( .D(N559), .CLK(clk), .RST(rst), .Q(o[270]) );
  DFF \oi_reg[8][15]  ( .D(N560), .CLK(clk), .RST(rst), .Q(o[271]) );
  DFF \oi_reg[8][16]  ( .D(N561), .CLK(clk), .RST(rst), .Q(o[272]) );
  DFF \oi_reg[8][17]  ( .D(N562), .CLK(clk), .RST(rst), .Q(o[273]) );
  DFF \oi_reg[8][18]  ( .D(N563), .CLK(clk), .RST(rst), .Q(o[274]) );
  DFF \oi_reg[8][19]  ( .D(N564), .CLK(clk), .RST(rst), .Q(o[275]) );
  DFF \oi_reg[8][20]  ( .D(N565), .CLK(clk), .RST(rst), .Q(o[276]) );
  DFF \oi_reg[8][21]  ( .D(N566), .CLK(clk), .RST(rst), .Q(o[277]) );
  DFF \oi_reg[8][22]  ( .D(N567), .CLK(clk), .RST(rst), .Q(o[278]) );
  DFF \oi_reg[8][23]  ( .D(N568), .CLK(clk), .RST(rst), .Q(o[279]) );
  DFF \oi_reg[8][24]  ( .D(N569), .CLK(clk), .RST(rst), .Q(o[280]) );
  DFF \oi_reg[8][25]  ( .D(N570), .CLK(clk), .RST(rst), .Q(o[281]) );
  DFF \oi_reg[8][26]  ( .D(N571), .CLK(clk), .RST(rst), .Q(o[282]) );
  DFF \oi_reg[8][27]  ( .D(N572), .CLK(clk), .RST(rst), .Q(o[283]) );
  DFF \oi_reg[8][28]  ( .D(N573), .CLK(clk), .RST(rst), .Q(o[284]) );
  DFF \oi_reg[8][29]  ( .D(N574), .CLK(clk), .RST(rst), .Q(o[285]) );
  DFF \oi_reg[8][30]  ( .D(N575), .CLK(clk), .RST(rst), .Q(o[286]) );
  DFF \oi_reg[8][31]  ( .D(N576), .CLK(clk), .RST(rst), .Q(o[287]) );
  DFF \oi_reg[9][0]  ( .D(N609), .CLK(clk), .RST(rst), .Q(o[288]) );
  DFF \oi_reg[9][1]  ( .D(N610), .CLK(clk), .RST(rst), .Q(o[289]) );
  DFF \oi_reg[9][2]  ( .D(N611), .CLK(clk), .RST(rst), .Q(o[290]) );
  DFF \oi_reg[9][3]  ( .D(N612), .CLK(clk), .RST(rst), .Q(o[291]) );
  DFF \oi_reg[9][4]  ( .D(N613), .CLK(clk), .RST(rst), .Q(o[292]) );
  DFF \oi_reg[9][5]  ( .D(N614), .CLK(clk), .RST(rst), .Q(o[293]) );
  DFF \oi_reg[9][6]  ( .D(N615), .CLK(clk), .RST(rst), .Q(o[294]) );
  DFF \oi_reg[9][7]  ( .D(N616), .CLK(clk), .RST(rst), .Q(o[295]) );
  DFF \oi_reg[9][8]  ( .D(N617), .CLK(clk), .RST(rst), .Q(o[296]) );
  DFF \oi_reg[9][9]  ( .D(N618), .CLK(clk), .RST(rst), .Q(o[297]) );
  DFF \oi_reg[9][10]  ( .D(N619), .CLK(clk), .RST(rst), .Q(o[298]) );
  DFF \oi_reg[9][11]  ( .D(N620), .CLK(clk), .RST(rst), .Q(o[299]) );
  DFF \oi_reg[9][12]  ( .D(N621), .CLK(clk), .RST(rst), .Q(o[300]) );
  DFF \oi_reg[9][13]  ( .D(N622), .CLK(clk), .RST(rst), .Q(o[301]) );
  DFF \oi_reg[9][14]  ( .D(N623), .CLK(clk), .RST(rst), .Q(o[302]) );
  DFF \oi_reg[9][15]  ( .D(N624), .CLK(clk), .RST(rst), .Q(o[303]) );
  DFF \oi_reg[9][16]  ( .D(N625), .CLK(clk), .RST(rst), .Q(o[304]) );
  DFF \oi_reg[9][17]  ( .D(N626), .CLK(clk), .RST(rst), .Q(o[305]) );
  DFF \oi_reg[9][18]  ( .D(N627), .CLK(clk), .RST(rst), .Q(o[306]) );
  DFF \oi_reg[9][19]  ( .D(N628), .CLK(clk), .RST(rst), .Q(o[307]) );
  DFF \oi_reg[9][20]  ( .D(N629), .CLK(clk), .RST(rst), .Q(o[308]) );
  DFF \oi_reg[9][21]  ( .D(N630), .CLK(clk), .RST(rst), .Q(o[309]) );
  DFF \oi_reg[9][22]  ( .D(N631), .CLK(clk), .RST(rst), .Q(o[310]) );
  DFF \oi_reg[9][23]  ( .D(N632), .CLK(clk), .RST(rst), .Q(o[311]) );
  DFF \oi_reg[9][24]  ( .D(N633), .CLK(clk), .RST(rst), .Q(o[312]) );
  DFF \oi_reg[9][25]  ( .D(N634), .CLK(clk), .RST(rst), .Q(o[313]) );
  DFF \oi_reg[9][26]  ( .D(N635), .CLK(clk), .RST(rst), .Q(o[314]) );
  DFF \oi_reg[9][27]  ( .D(N636), .CLK(clk), .RST(rst), .Q(o[315]) );
  DFF \oi_reg[9][28]  ( .D(N637), .CLK(clk), .RST(rst), .Q(o[316]) );
  DFF \oi_reg[9][29]  ( .D(N638), .CLK(clk), .RST(rst), .Q(o[317]) );
  DFF \oi_reg[9][30]  ( .D(N639), .CLK(clk), .RST(rst), .Q(o[318]) );
  DFF \oi_reg[9][31]  ( .D(N640), .CLK(clk), .RST(rst), .Q(o[319]) );
  DFF \oi_reg[10][0]  ( .D(N673), .CLK(clk), .RST(rst), .Q(o[320]) );
  DFF \oi_reg[10][1]  ( .D(N674), .CLK(clk), .RST(rst), .Q(o[321]) );
  DFF \oi_reg[10][2]  ( .D(N675), .CLK(clk), .RST(rst), .Q(o[322]) );
  DFF \oi_reg[10][3]  ( .D(N676), .CLK(clk), .RST(rst), .Q(o[323]) );
  DFF \oi_reg[10][4]  ( .D(N677), .CLK(clk), .RST(rst), .Q(o[324]) );
  DFF \oi_reg[10][5]  ( .D(N678), .CLK(clk), .RST(rst), .Q(o[325]) );
  DFF \oi_reg[10][6]  ( .D(N679), .CLK(clk), .RST(rst), .Q(o[326]) );
  DFF \oi_reg[10][7]  ( .D(N680), .CLK(clk), .RST(rst), .Q(o[327]) );
  DFF \oi_reg[10][8]  ( .D(N681), .CLK(clk), .RST(rst), .Q(o[328]) );
  DFF \oi_reg[10][9]  ( .D(N682), .CLK(clk), .RST(rst), .Q(o[329]) );
  DFF \oi_reg[10][10]  ( .D(N683), .CLK(clk), .RST(rst), .Q(o[330]) );
  DFF \oi_reg[10][11]  ( .D(N684), .CLK(clk), .RST(rst), .Q(o[331]) );
  DFF \oi_reg[10][12]  ( .D(N685), .CLK(clk), .RST(rst), .Q(o[332]) );
  DFF \oi_reg[10][13]  ( .D(N686), .CLK(clk), .RST(rst), .Q(o[333]) );
  DFF \oi_reg[10][14]  ( .D(N687), .CLK(clk), .RST(rst), .Q(o[334]) );
  DFF \oi_reg[10][15]  ( .D(N688), .CLK(clk), .RST(rst), .Q(o[335]) );
  DFF \oi_reg[10][16]  ( .D(N689), .CLK(clk), .RST(rst), .Q(o[336]) );
  DFF \oi_reg[10][17]  ( .D(N690), .CLK(clk), .RST(rst), .Q(o[337]) );
  DFF \oi_reg[10][18]  ( .D(N691), .CLK(clk), .RST(rst), .Q(o[338]) );
  DFF \oi_reg[10][19]  ( .D(N692), .CLK(clk), .RST(rst), .Q(o[339]) );
  DFF \oi_reg[10][20]  ( .D(N693), .CLK(clk), .RST(rst), .Q(o[340]) );
  DFF \oi_reg[10][21]  ( .D(N694), .CLK(clk), .RST(rst), .Q(o[341]) );
  DFF \oi_reg[10][22]  ( .D(N695), .CLK(clk), .RST(rst), .Q(o[342]) );
  DFF \oi_reg[10][23]  ( .D(N696), .CLK(clk), .RST(rst), .Q(o[343]) );
  DFF \oi_reg[10][24]  ( .D(N697), .CLK(clk), .RST(rst), .Q(o[344]) );
  DFF \oi_reg[10][25]  ( .D(N698), .CLK(clk), .RST(rst), .Q(o[345]) );
  DFF \oi_reg[10][26]  ( .D(N699), .CLK(clk), .RST(rst), .Q(o[346]) );
  DFF \oi_reg[10][27]  ( .D(N700), .CLK(clk), .RST(rst), .Q(o[347]) );
  DFF \oi_reg[10][28]  ( .D(N701), .CLK(clk), .RST(rst), .Q(o[348]) );
  DFF \oi_reg[10][29]  ( .D(N702), .CLK(clk), .RST(rst), .Q(o[349]) );
  DFF \oi_reg[10][30]  ( .D(N703), .CLK(clk), .RST(rst), .Q(o[350]) );
  DFF \oi_reg[10][31]  ( .D(N704), .CLK(clk), .RST(rst), .Q(o[351]) );
  DFF \oi_reg[11][0]  ( .D(N737), .CLK(clk), .RST(rst), .Q(o[352]) );
  DFF \oi_reg[11][1]  ( .D(N738), .CLK(clk), .RST(rst), .Q(o[353]) );
  DFF \oi_reg[11][2]  ( .D(N739), .CLK(clk), .RST(rst), .Q(o[354]) );
  DFF \oi_reg[11][3]  ( .D(N740), .CLK(clk), .RST(rst), .Q(o[355]) );
  DFF \oi_reg[11][4]  ( .D(N741), .CLK(clk), .RST(rst), .Q(o[356]) );
  DFF \oi_reg[11][5]  ( .D(N742), .CLK(clk), .RST(rst), .Q(o[357]) );
  DFF \oi_reg[11][6]  ( .D(N743), .CLK(clk), .RST(rst), .Q(o[358]) );
  DFF \oi_reg[11][7]  ( .D(N744), .CLK(clk), .RST(rst), .Q(o[359]) );
  DFF \oi_reg[11][8]  ( .D(N745), .CLK(clk), .RST(rst), .Q(o[360]) );
  DFF \oi_reg[11][9]  ( .D(N746), .CLK(clk), .RST(rst), .Q(o[361]) );
  DFF \oi_reg[11][10]  ( .D(N747), .CLK(clk), .RST(rst), .Q(o[362]) );
  DFF \oi_reg[11][11]  ( .D(N748), .CLK(clk), .RST(rst), .Q(o[363]) );
  DFF \oi_reg[11][12]  ( .D(N749), .CLK(clk), .RST(rst), .Q(o[364]) );
  DFF \oi_reg[11][13]  ( .D(N750), .CLK(clk), .RST(rst), .Q(o[365]) );
  DFF \oi_reg[11][14]  ( .D(N751), .CLK(clk), .RST(rst), .Q(o[366]) );
  DFF \oi_reg[11][15]  ( .D(N752), .CLK(clk), .RST(rst), .Q(o[367]) );
  DFF \oi_reg[11][16]  ( .D(N753), .CLK(clk), .RST(rst), .Q(o[368]) );
  DFF \oi_reg[11][17]  ( .D(N754), .CLK(clk), .RST(rst), .Q(o[369]) );
  DFF \oi_reg[11][18]  ( .D(N755), .CLK(clk), .RST(rst), .Q(o[370]) );
  DFF \oi_reg[11][19]  ( .D(N756), .CLK(clk), .RST(rst), .Q(o[371]) );
  DFF \oi_reg[11][20]  ( .D(N757), .CLK(clk), .RST(rst), .Q(o[372]) );
  DFF \oi_reg[11][21]  ( .D(N758), .CLK(clk), .RST(rst), .Q(o[373]) );
  DFF \oi_reg[11][22]  ( .D(N759), .CLK(clk), .RST(rst), .Q(o[374]) );
  DFF \oi_reg[11][23]  ( .D(N760), .CLK(clk), .RST(rst), .Q(o[375]) );
  DFF \oi_reg[11][24]  ( .D(N761), .CLK(clk), .RST(rst), .Q(o[376]) );
  DFF \oi_reg[11][25]  ( .D(N762), .CLK(clk), .RST(rst), .Q(o[377]) );
  DFF \oi_reg[11][26]  ( .D(N763), .CLK(clk), .RST(rst), .Q(o[378]) );
  DFF \oi_reg[11][27]  ( .D(N764), .CLK(clk), .RST(rst), .Q(o[379]) );
  DFF \oi_reg[11][28]  ( .D(N765), .CLK(clk), .RST(rst), .Q(o[380]) );
  DFF \oi_reg[11][29]  ( .D(N766), .CLK(clk), .RST(rst), .Q(o[381]) );
  DFF \oi_reg[11][30]  ( .D(N767), .CLK(clk), .RST(rst), .Q(o[382]) );
  DFF \oi_reg[11][31]  ( .D(N768), .CLK(clk), .RST(rst), .Q(o[383]) );
  DFF \oi_reg[12][0]  ( .D(N801), .CLK(clk), .RST(rst), .Q(o[384]) );
  DFF \oi_reg[12][1]  ( .D(N802), .CLK(clk), .RST(rst), .Q(o[385]) );
  DFF \oi_reg[12][2]  ( .D(N803), .CLK(clk), .RST(rst), .Q(o[386]) );
  DFF \oi_reg[12][3]  ( .D(N804), .CLK(clk), .RST(rst), .Q(o[387]) );
  DFF \oi_reg[12][4]  ( .D(N805), .CLK(clk), .RST(rst), .Q(o[388]) );
  DFF \oi_reg[12][5]  ( .D(N806), .CLK(clk), .RST(rst), .Q(o[389]) );
  DFF \oi_reg[12][6]  ( .D(N807), .CLK(clk), .RST(rst), .Q(o[390]) );
  DFF \oi_reg[12][7]  ( .D(N808), .CLK(clk), .RST(rst), .Q(o[391]) );
  DFF \oi_reg[12][8]  ( .D(N809), .CLK(clk), .RST(rst), .Q(o[392]) );
  DFF \oi_reg[12][9]  ( .D(N810), .CLK(clk), .RST(rst), .Q(o[393]) );
  DFF \oi_reg[12][10]  ( .D(N811), .CLK(clk), .RST(rst), .Q(o[394]) );
  DFF \oi_reg[12][11]  ( .D(N812), .CLK(clk), .RST(rst), .Q(o[395]) );
  DFF \oi_reg[12][12]  ( .D(N813), .CLK(clk), .RST(rst), .Q(o[396]) );
  DFF \oi_reg[12][13]  ( .D(N814), .CLK(clk), .RST(rst), .Q(o[397]) );
  DFF \oi_reg[12][14]  ( .D(N815), .CLK(clk), .RST(rst), .Q(o[398]) );
  DFF \oi_reg[12][15]  ( .D(N816), .CLK(clk), .RST(rst), .Q(o[399]) );
  DFF \oi_reg[12][16]  ( .D(N817), .CLK(clk), .RST(rst), .Q(o[400]) );
  DFF \oi_reg[12][17]  ( .D(N818), .CLK(clk), .RST(rst), .Q(o[401]) );
  DFF \oi_reg[12][18]  ( .D(N819), .CLK(clk), .RST(rst), .Q(o[402]) );
  DFF \oi_reg[12][19]  ( .D(N820), .CLK(clk), .RST(rst), .Q(o[403]) );
  DFF \oi_reg[12][20]  ( .D(N821), .CLK(clk), .RST(rst), .Q(o[404]) );
  DFF \oi_reg[12][21]  ( .D(N822), .CLK(clk), .RST(rst), .Q(o[405]) );
  DFF \oi_reg[12][22]  ( .D(N823), .CLK(clk), .RST(rst), .Q(o[406]) );
  DFF \oi_reg[12][23]  ( .D(N824), .CLK(clk), .RST(rst), .Q(o[407]) );
  DFF \oi_reg[12][24]  ( .D(N825), .CLK(clk), .RST(rst), .Q(o[408]) );
  DFF \oi_reg[12][25]  ( .D(N826), .CLK(clk), .RST(rst), .Q(o[409]) );
  DFF \oi_reg[12][26]  ( .D(N827), .CLK(clk), .RST(rst), .Q(o[410]) );
  DFF \oi_reg[12][27]  ( .D(N828), .CLK(clk), .RST(rst), .Q(o[411]) );
  DFF \oi_reg[12][28]  ( .D(N829), .CLK(clk), .RST(rst), .Q(o[412]) );
  DFF \oi_reg[12][29]  ( .D(N830), .CLK(clk), .RST(rst), .Q(o[413]) );
  DFF \oi_reg[12][30]  ( .D(N831), .CLK(clk), .RST(rst), .Q(o[414]) );
  DFF \oi_reg[12][31]  ( .D(N832), .CLK(clk), .RST(rst), .Q(o[415]) );
  DFF \oi_reg[13][0]  ( .D(N865), .CLK(clk), .RST(rst), .Q(o[416]) );
  DFF \oi_reg[13][1]  ( .D(N866), .CLK(clk), .RST(rst), .Q(o[417]) );
  DFF \oi_reg[13][2]  ( .D(N867), .CLK(clk), .RST(rst), .Q(o[418]) );
  DFF \oi_reg[13][3]  ( .D(N868), .CLK(clk), .RST(rst), .Q(o[419]) );
  DFF \oi_reg[13][4]  ( .D(N869), .CLK(clk), .RST(rst), .Q(o[420]) );
  DFF \oi_reg[13][5]  ( .D(N870), .CLK(clk), .RST(rst), .Q(o[421]) );
  DFF \oi_reg[13][6]  ( .D(N871), .CLK(clk), .RST(rst), .Q(o[422]) );
  DFF \oi_reg[13][7]  ( .D(N872), .CLK(clk), .RST(rst), .Q(o[423]) );
  DFF \oi_reg[13][8]  ( .D(N873), .CLK(clk), .RST(rst), .Q(o[424]) );
  DFF \oi_reg[13][9]  ( .D(N874), .CLK(clk), .RST(rst), .Q(o[425]) );
  DFF \oi_reg[13][10]  ( .D(N875), .CLK(clk), .RST(rst), .Q(o[426]) );
  DFF \oi_reg[13][11]  ( .D(N876), .CLK(clk), .RST(rst), .Q(o[427]) );
  DFF \oi_reg[13][12]  ( .D(N877), .CLK(clk), .RST(rst), .Q(o[428]) );
  DFF \oi_reg[13][13]  ( .D(N878), .CLK(clk), .RST(rst), .Q(o[429]) );
  DFF \oi_reg[13][14]  ( .D(N879), .CLK(clk), .RST(rst), .Q(o[430]) );
  DFF \oi_reg[13][15]  ( .D(N880), .CLK(clk), .RST(rst), .Q(o[431]) );
  DFF \oi_reg[13][16]  ( .D(N881), .CLK(clk), .RST(rst), .Q(o[432]) );
  DFF \oi_reg[13][17]  ( .D(N882), .CLK(clk), .RST(rst), .Q(o[433]) );
  DFF \oi_reg[13][18]  ( .D(N883), .CLK(clk), .RST(rst), .Q(o[434]) );
  DFF \oi_reg[13][19]  ( .D(N884), .CLK(clk), .RST(rst), .Q(o[435]) );
  DFF \oi_reg[13][20]  ( .D(N885), .CLK(clk), .RST(rst), .Q(o[436]) );
  DFF \oi_reg[13][21]  ( .D(N886), .CLK(clk), .RST(rst), .Q(o[437]) );
  DFF \oi_reg[13][22]  ( .D(N887), .CLK(clk), .RST(rst), .Q(o[438]) );
  DFF \oi_reg[13][23]  ( .D(N888), .CLK(clk), .RST(rst), .Q(o[439]) );
  DFF \oi_reg[13][24]  ( .D(N889), .CLK(clk), .RST(rst), .Q(o[440]) );
  DFF \oi_reg[13][25]  ( .D(N890), .CLK(clk), .RST(rst), .Q(o[441]) );
  DFF \oi_reg[13][26]  ( .D(N891), .CLK(clk), .RST(rst), .Q(o[442]) );
  DFF \oi_reg[13][27]  ( .D(N892), .CLK(clk), .RST(rst), .Q(o[443]) );
  DFF \oi_reg[13][28]  ( .D(N893), .CLK(clk), .RST(rst), .Q(o[444]) );
  DFF \oi_reg[13][29]  ( .D(N894), .CLK(clk), .RST(rst), .Q(o[445]) );
  DFF \oi_reg[13][30]  ( .D(N895), .CLK(clk), .RST(rst), .Q(o[446]) );
  DFF \oi_reg[13][31]  ( .D(N896), .CLK(clk), .RST(rst), .Q(o[447]) );
  DFF \oi_reg[14][0]  ( .D(N929), .CLK(clk), .RST(rst), .Q(o[448]) );
  DFF \oi_reg[14][1]  ( .D(N930), .CLK(clk), .RST(rst), .Q(o[449]) );
  DFF \oi_reg[14][2]  ( .D(N931), .CLK(clk), .RST(rst), .Q(o[450]) );
  DFF \oi_reg[14][3]  ( .D(N932), .CLK(clk), .RST(rst), .Q(o[451]) );
  DFF \oi_reg[14][4]  ( .D(N933), .CLK(clk), .RST(rst), .Q(o[452]) );
  DFF \oi_reg[14][5]  ( .D(N934), .CLK(clk), .RST(rst), .Q(o[453]) );
  DFF \oi_reg[14][6]  ( .D(N935), .CLK(clk), .RST(rst), .Q(o[454]) );
  DFF \oi_reg[14][7]  ( .D(N936), .CLK(clk), .RST(rst), .Q(o[455]) );
  DFF \oi_reg[14][8]  ( .D(N937), .CLK(clk), .RST(rst), .Q(o[456]) );
  DFF \oi_reg[14][9]  ( .D(N938), .CLK(clk), .RST(rst), .Q(o[457]) );
  DFF \oi_reg[14][10]  ( .D(N939), .CLK(clk), .RST(rst), .Q(o[458]) );
  DFF \oi_reg[14][11]  ( .D(N940), .CLK(clk), .RST(rst), .Q(o[459]) );
  DFF \oi_reg[14][12]  ( .D(N941), .CLK(clk), .RST(rst), .Q(o[460]) );
  DFF \oi_reg[14][13]  ( .D(N942), .CLK(clk), .RST(rst), .Q(o[461]) );
  DFF \oi_reg[14][14]  ( .D(N943), .CLK(clk), .RST(rst), .Q(o[462]) );
  DFF \oi_reg[14][15]  ( .D(N944), .CLK(clk), .RST(rst), .Q(o[463]) );
  DFF \oi_reg[14][16]  ( .D(N945), .CLK(clk), .RST(rst), .Q(o[464]) );
  DFF \oi_reg[14][17]  ( .D(N946), .CLK(clk), .RST(rst), .Q(o[465]) );
  DFF \oi_reg[14][18]  ( .D(N947), .CLK(clk), .RST(rst), .Q(o[466]) );
  DFF \oi_reg[14][19]  ( .D(N948), .CLK(clk), .RST(rst), .Q(o[467]) );
  DFF \oi_reg[14][20]  ( .D(N949), .CLK(clk), .RST(rst), .Q(o[468]) );
  DFF \oi_reg[14][21]  ( .D(N950), .CLK(clk), .RST(rst), .Q(o[469]) );
  DFF \oi_reg[14][22]  ( .D(N951), .CLK(clk), .RST(rst), .Q(o[470]) );
  DFF \oi_reg[14][23]  ( .D(N952), .CLK(clk), .RST(rst), .Q(o[471]) );
  DFF \oi_reg[14][24]  ( .D(N953), .CLK(clk), .RST(rst), .Q(o[472]) );
  DFF \oi_reg[14][25]  ( .D(N954), .CLK(clk), .RST(rst), .Q(o[473]) );
  DFF \oi_reg[14][26]  ( .D(N955), .CLK(clk), .RST(rst), .Q(o[474]) );
  DFF \oi_reg[14][27]  ( .D(N956), .CLK(clk), .RST(rst), .Q(o[475]) );
  DFF \oi_reg[14][28]  ( .D(N957), .CLK(clk), .RST(rst), .Q(o[476]) );
  DFF \oi_reg[14][29]  ( .D(N958), .CLK(clk), .RST(rst), .Q(o[477]) );
  DFF \oi_reg[14][30]  ( .D(N959), .CLK(clk), .RST(rst), .Q(o[478]) );
  DFF \oi_reg[14][31]  ( .D(N960), .CLK(clk), .RST(rst), .Q(o[479]) );
  DFF \oi_reg[15][0]  ( .D(N993), .CLK(clk), .RST(rst), .Q(o[480]) );
  DFF \oi_reg[15][1]  ( .D(N994), .CLK(clk), .RST(rst), .Q(o[481]) );
  DFF \oi_reg[15][2]  ( .D(N995), .CLK(clk), .RST(rst), .Q(o[482]) );
  DFF \oi_reg[15][3]  ( .D(N996), .CLK(clk), .RST(rst), .Q(o[483]) );
  DFF \oi_reg[15][4]  ( .D(N997), .CLK(clk), .RST(rst), .Q(o[484]) );
  DFF \oi_reg[15][5]  ( .D(N998), .CLK(clk), .RST(rst), .Q(o[485]) );
  DFF \oi_reg[15][6]  ( .D(N999), .CLK(clk), .RST(rst), .Q(o[486]) );
  DFF \oi_reg[15][7]  ( .D(N1000), .CLK(clk), .RST(rst), .Q(o[487]) );
  DFF \oi_reg[15][8]  ( .D(N1001), .CLK(clk), .RST(rst), .Q(o[488]) );
  DFF \oi_reg[15][9]  ( .D(N1002), .CLK(clk), .RST(rst), .Q(o[489]) );
  DFF \oi_reg[15][10]  ( .D(N1003), .CLK(clk), .RST(rst), .Q(o[490]) );
  DFF \oi_reg[15][11]  ( .D(N1004), .CLK(clk), .RST(rst), .Q(o[491]) );
  DFF \oi_reg[15][12]  ( .D(N1005), .CLK(clk), .RST(rst), .Q(o[492]) );
  DFF \oi_reg[15][13]  ( .D(N1006), .CLK(clk), .RST(rst), .Q(o[493]) );
  DFF \oi_reg[15][14]  ( .D(N1007), .CLK(clk), .RST(rst), .Q(o[494]) );
  DFF \oi_reg[15][15]  ( .D(N1008), .CLK(clk), .RST(rst), .Q(o[495]) );
  DFF \oi_reg[15][16]  ( .D(N1009), .CLK(clk), .RST(rst), .Q(o[496]) );
  DFF \oi_reg[15][17]  ( .D(N1010), .CLK(clk), .RST(rst), .Q(o[497]) );
  DFF \oi_reg[15][18]  ( .D(N1011), .CLK(clk), .RST(rst), .Q(o[498]) );
  DFF \oi_reg[15][19]  ( .D(N1012), .CLK(clk), .RST(rst), .Q(o[499]) );
  DFF \oi_reg[15][20]  ( .D(N1013), .CLK(clk), .RST(rst), .Q(o[500]) );
  DFF \oi_reg[15][21]  ( .D(N1014), .CLK(clk), .RST(rst), .Q(o[501]) );
  DFF \oi_reg[15][22]  ( .D(N1015), .CLK(clk), .RST(rst), .Q(o[502]) );
  DFF \oi_reg[15][23]  ( .D(N1016), .CLK(clk), .RST(rst), .Q(o[503]) );
  DFF \oi_reg[15][24]  ( .D(N1017), .CLK(clk), .RST(rst), .Q(o[504]) );
  DFF \oi_reg[15][25]  ( .D(N1018), .CLK(clk), .RST(rst), .Q(o[505]) );
  DFF \oi_reg[15][26]  ( .D(N1019), .CLK(clk), .RST(rst), .Q(o[506]) );
  DFF \oi_reg[15][27]  ( .D(N1020), .CLK(clk), .RST(rst), .Q(o[507]) );
  DFF \oi_reg[15][28]  ( .D(N1021), .CLK(clk), .RST(rst), .Q(o[508]) );
  DFF \oi_reg[15][29]  ( .D(N1022), .CLK(clk), .RST(rst), .Q(o[509]) );
  DFF \oi_reg[15][30]  ( .D(N1023), .CLK(clk), .RST(rst), .Q(o[510]) );
  DFF \oi_reg[15][31]  ( .D(N1024), .CLK(clk), .RST(rst), .Q(o[511]) );
  matrixMult_N_M_1_N16_M32_DW01_add_0 add_54_I16_G16 ( .A(o[511:480]), .B({
        N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, 
        N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, 
        N968, N967, N966, N965, N964, N963, N962, N961}), .CI(1'b0), .SUM({
        N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, 
        N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, 
        N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, 
        N993}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_0 mult_54_I16_G16 ( .A(x[511:480]), .B(
        y[8191:8160]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, N992, N991, N990, N989, N988, N987, N986, 
        N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, 
        N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, 
        N961}) );
  matrixMult_N_M_1_N16_M32_DW01_add_2 add_54_I16_G15 ( .A(o[479:448]), .B({
        N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, 
        N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, 
        N904, N903, N902, N901, N900, N899, N898, N897}), .CI(1'b0), .SUM({
        N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, 
        N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, 
        N936, N935, N934, N933, N932, N931, N930, N929}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_1 mult_54_I16_G15 ( .A(x[511:480]), .B(
        y[8159:8128]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, N928, N927, N926, N925, N924, N923, N922, 
        N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, 
        N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, 
        N897}) );
  matrixMult_N_M_1_N16_M32_DW01_add_4 add_54_I16_G14 ( .A(o[447:416]), .B({
        N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, 
        N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, 
        N840, N839, N838, N837, N836, N835, N834, N833}), .CI(1'b0), .SUM({
        N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, 
        N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, 
        N872, N871, N870, N869, N868, N867, N866, N865}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_2 mult_54_I16_G14 ( .A(x[511:480]), .B(
        y[8127:8096]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, N864, N863, N862, N861, N860, N859, N858, 
        N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, 
        N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, 
        N833}) );
  matrixMult_N_M_1_N16_M32_DW01_add_6 add_54_I16_G13 ( .A(o[415:384]), .B({
        N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, 
        N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, 
        N776, N775, N774, N773, N772, N771, N770, N769}), .CI(1'b0), .SUM({
        N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, 
        N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, 
        N808, N807, N806, N805, N804, N803, N802, N801}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_3 mult_54_I16_G13 ( .A(x[511:480]), .B(
        y[8095:8064]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, N800, N799, N798, N797, N796, N795, N794, 
        N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, 
        N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, 
        N769}) );
  matrixMult_N_M_1_N16_M32_DW01_add_8 add_54_I16_G12 ( .A(o[383:352]), .B({
        N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, 
        N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, 
        N712, N711, N710, N709, N708, N707, N706, N705}), .CI(1'b0), .SUM({
        N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, 
        N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, 
        N744, N743, N742, N741, N740, N739, N738, N737}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_4 mult_54_I16_G12 ( .A(x[511:480]), .B(
        y[8063:8032]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, N736, N735, N734, N733, N732, N731, N730, 
        N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, 
        N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, 
        N705}) );
  matrixMult_N_M_1_N16_M32_DW01_add_10 add_54_I16_G11 ( .A(o[351:320]), .B({
        N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, 
        N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, 
        N648, N647, N646, N645, N644, N643, N642, N641}), .CI(1'b0), .SUM({
        N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, 
        N680, N679, N678, N677, N676, N675, N674, N673}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_5 mult_54_I16_G11 ( .A(x[511:480]), .B(
        y[8031:8000]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, 
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, 
        SYNOPSYS_UNCONNECTED__191, N672, N671, N670, N669, N668, N667, N666, 
        N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, 
        N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, 
        N641}) );
  matrixMult_N_M_1_N16_M32_DW01_add_12 add_54_I16_G10 ( .A(o[319:288]), .B({
        N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, N581, N580, N579, N578, N577}), .CI(1'b0), .SUM({
        N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, 
        N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, 
        N616, N615, N614, N613, N612, N611, N610, N609}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_6 mult_54_I16_G10 ( .A(x[511:480]), .B(
        y[7999:7968]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__192, 
        SYNOPSYS_UNCONNECTED__193, SYNOPSYS_UNCONNECTED__194, 
        SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, 
        SYNOPSYS_UNCONNECTED__197, SYNOPSYS_UNCONNECTED__198, 
        SYNOPSYS_UNCONNECTED__199, SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, 
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, 
        SYNOPSYS_UNCONNECTED__211, SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213, SYNOPSYS_UNCONNECTED__214, 
        SYNOPSYS_UNCONNECTED__215, SYNOPSYS_UNCONNECTED__216, 
        SYNOPSYS_UNCONNECTED__217, SYNOPSYS_UNCONNECTED__218, 
        SYNOPSYS_UNCONNECTED__219, SYNOPSYS_UNCONNECTED__220, 
        SYNOPSYS_UNCONNECTED__221, SYNOPSYS_UNCONNECTED__222, 
        SYNOPSYS_UNCONNECTED__223, N608, N607, N606, N605, N604, N603, N602, 
        N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, 
        N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, 
        N577}) );
  matrixMult_N_M_1_N16_M32_DW01_add_14 add_54_I16_G9 ( .A(o[287:256]), .B({
        N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, 
        N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, 
        N520, N519, N518, N517, N516, N515, N514, N513}), .CI(1'b0), .SUM({
        N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, 
        N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, 
        N552, N551, N550, N549, N548, N547, N546, N545}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_7 mult_54_I16_G9 ( .A(x[511:480]), .B(
        y[7967:7936]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, 
        SYNOPSYS_UNCONNECTED__227, SYNOPSYS_UNCONNECTED__228, 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, SYNOPSYS_UNCONNECTED__232, 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, 
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, 
        SYNOPSYS_UNCONNECTED__247, SYNOPSYS_UNCONNECTED__248, 
        SYNOPSYS_UNCONNECTED__249, SYNOPSYS_UNCONNECTED__250, 
        SYNOPSYS_UNCONNECTED__251, SYNOPSYS_UNCONNECTED__252, 
        SYNOPSYS_UNCONNECTED__253, SYNOPSYS_UNCONNECTED__254, 
        SYNOPSYS_UNCONNECTED__255, N544, N543, N542, N541, N540, N539, N538, 
        N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, 
        N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, 
        N513}) );
  matrixMult_N_M_1_N16_M32_DW01_add_16 add_54_I16_G8 ( .A(o[255:224]), .B({
        N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, 
        N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, 
        N456, N455, N454, N453, N452, N451, N450, N449}), .CI(1'b0), .SUM({
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N485, N484, N483, N482, N481}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_8 mult_54_I16_G8 ( .A(x[511:480]), .B(
        y[7935:7904]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__256, 
        SYNOPSYS_UNCONNECTED__257, SYNOPSYS_UNCONNECTED__258, 
        SYNOPSYS_UNCONNECTED__259, SYNOPSYS_UNCONNECTED__260, 
        SYNOPSYS_UNCONNECTED__261, SYNOPSYS_UNCONNECTED__262, 
        SYNOPSYS_UNCONNECTED__263, SYNOPSYS_UNCONNECTED__264, 
        SYNOPSYS_UNCONNECTED__265, SYNOPSYS_UNCONNECTED__266, 
        SYNOPSYS_UNCONNECTED__267, SYNOPSYS_UNCONNECTED__268, 
        SYNOPSYS_UNCONNECTED__269, SYNOPSYS_UNCONNECTED__270, 
        SYNOPSYS_UNCONNECTED__271, SYNOPSYS_UNCONNECTED__272, 
        SYNOPSYS_UNCONNECTED__273, SYNOPSYS_UNCONNECTED__274, 
        SYNOPSYS_UNCONNECTED__275, SYNOPSYS_UNCONNECTED__276, 
        SYNOPSYS_UNCONNECTED__277, SYNOPSYS_UNCONNECTED__278, 
        SYNOPSYS_UNCONNECTED__279, SYNOPSYS_UNCONNECTED__280, 
        SYNOPSYS_UNCONNECTED__281, SYNOPSYS_UNCONNECTED__282, 
        SYNOPSYS_UNCONNECTED__283, SYNOPSYS_UNCONNECTED__284, 
        SYNOPSYS_UNCONNECTED__285, SYNOPSYS_UNCONNECTED__286, 
        SYNOPSYS_UNCONNECTED__287, N480, N479, N478, N477, N476, N475, N474, 
        N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, 
        N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, 
        N449}) );
  matrixMult_N_M_1_N16_M32_DW01_add_18 add_54_I16_G7 ( .A(o[223:192]), .B({
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385}), .CI(1'b0), .SUM({
        N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, 
        N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, 
        N424, N423, N422, N421, N420, N419, N418, N417}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_9 mult_54_I16_G7 ( .A(x[511:480]), .B(
        y[7903:7872]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__288, 
        SYNOPSYS_UNCONNECTED__289, SYNOPSYS_UNCONNECTED__290, 
        SYNOPSYS_UNCONNECTED__291, SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, SYNOPSYS_UNCONNECTED__296, 
        SYNOPSYS_UNCONNECTED__297, SYNOPSYS_UNCONNECTED__298, 
        SYNOPSYS_UNCONNECTED__299, SYNOPSYS_UNCONNECTED__300, 
        SYNOPSYS_UNCONNECTED__301, SYNOPSYS_UNCONNECTED__302, 
        SYNOPSYS_UNCONNECTED__303, SYNOPSYS_UNCONNECTED__304, 
        SYNOPSYS_UNCONNECTED__305, SYNOPSYS_UNCONNECTED__306, 
        SYNOPSYS_UNCONNECTED__307, SYNOPSYS_UNCONNECTED__308, 
        SYNOPSYS_UNCONNECTED__309, SYNOPSYS_UNCONNECTED__310, 
        SYNOPSYS_UNCONNECTED__311, SYNOPSYS_UNCONNECTED__312, 
        SYNOPSYS_UNCONNECTED__313, SYNOPSYS_UNCONNECTED__314, 
        SYNOPSYS_UNCONNECTED__315, SYNOPSYS_UNCONNECTED__316, 
        SYNOPSYS_UNCONNECTED__317, SYNOPSYS_UNCONNECTED__318, 
        SYNOPSYS_UNCONNECTED__319, N416, N415, N414, N413, N412, N411, N410, 
        N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, 
        N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, 
        N385}) );
  matrixMult_N_M_1_N16_M32_DW01_add_20 add_54_I16_G6 ( .A(o[191:160]), .B({
        N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, 
        N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, 
        N328, N327, N326, N325, N324, N323, N322, N321}), .CI(1'b0), .SUM({
        N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, 
        N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, 
        N360, N359, N358, N357, N356, N355, N354, N353}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_10 mult_54_I16_G6 ( .A(x[511:480]), .B(
        y[7871:7840]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__320, 
        SYNOPSYS_UNCONNECTED__321, SYNOPSYS_UNCONNECTED__322, 
        SYNOPSYS_UNCONNECTED__323, SYNOPSYS_UNCONNECTED__324, 
        SYNOPSYS_UNCONNECTED__325, SYNOPSYS_UNCONNECTED__326, 
        SYNOPSYS_UNCONNECTED__327, SYNOPSYS_UNCONNECTED__328, 
        SYNOPSYS_UNCONNECTED__329, SYNOPSYS_UNCONNECTED__330, 
        SYNOPSYS_UNCONNECTED__331, SYNOPSYS_UNCONNECTED__332, 
        SYNOPSYS_UNCONNECTED__333, SYNOPSYS_UNCONNECTED__334, 
        SYNOPSYS_UNCONNECTED__335, SYNOPSYS_UNCONNECTED__336, 
        SYNOPSYS_UNCONNECTED__337, SYNOPSYS_UNCONNECTED__338, 
        SYNOPSYS_UNCONNECTED__339, SYNOPSYS_UNCONNECTED__340, 
        SYNOPSYS_UNCONNECTED__341, SYNOPSYS_UNCONNECTED__342, 
        SYNOPSYS_UNCONNECTED__343, SYNOPSYS_UNCONNECTED__344, 
        SYNOPSYS_UNCONNECTED__345, SYNOPSYS_UNCONNECTED__346, 
        SYNOPSYS_UNCONNECTED__347, SYNOPSYS_UNCONNECTED__348, 
        SYNOPSYS_UNCONNECTED__349, SYNOPSYS_UNCONNECTED__350, 
        SYNOPSYS_UNCONNECTED__351, N352, N351, N350, N349, N348, N347, N346, 
        N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, 
        N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, 
        N321}) );
  matrixMult_N_M_1_N16_M32_DW01_add_22 add_54_I16_G5 ( .A(o[159:128]), .B({
        N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, 
        N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257}), .CI(1'b0), .SUM({
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_11 mult_54_I16_G5 ( .A(x[511:480]), .B(
        y[7839:7808]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__352, 
        SYNOPSYS_UNCONNECTED__353, SYNOPSYS_UNCONNECTED__354, 
        SYNOPSYS_UNCONNECTED__355, SYNOPSYS_UNCONNECTED__356, 
        SYNOPSYS_UNCONNECTED__357, SYNOPSYS_UNCONNECTED__358, 
        SYNOPSYS_UNCONNECTED__359, SYNOPSYS_UNCONNECTED__360, 
        SYNOPSYS_UNCONNECTED__361, SYNOPSYS_UNCONNECTED__362, 
        SYNOPSYS_UNCONNECTED__363, SYNOPSYS_UNCONNECTED__364, 
        SYNOPSYS_UNCONNECTED__365, SYNOPSYS_UNCONNECTED__366, 
        SYNOPSYS_UNCONNECTED__367, SYNOPSYS_UNCONNECTED__368, 
        SYNOPSYS_UNCONNECTED__369, SYNOPSYS_UNCONNECTED__370, 
        SYNOPSYS_UNCONNECTED__371, SYNOPSYS_UNCONNECTED__372, 
        SYNOPSYS_UNCONNECTED__373, SYNOPSYS_UNCONNECTED__374, 
        SYNOPSYS_UNCONNECTED__375, SYNOPSYS_UNCONNECTED__376, 
        SYNOPSYS_UNCONNECTED__377, SYNOPSYS_UNCONNECTED__378, 
        SYNOPSYS_UNCONNECTED__379, SYNOPSYS_UNCONNECTED__380, 
        SYNOPSYS_UNCONNECTED__381, SYNOPSYS_UNCONNECTED__382, 
        SYNOPSYS_UNCONNECTED__383, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, 
        N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, 
        N257}) );
  matrixMult_N_M_1_N16_M32_DW01_add_24 add_54_I16_G4 ( .A(o[127:96]), .B({N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193}), .CI(1'b0), .SUM({N256, 
        N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, 
        N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, 
        N231, N230, N229, N228, N227, N226, N225}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_12 mult_54_I16_G4 ( .A(x[511:480]), .B(
        y[7807:7776]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__384, 
        SYNOPSYS_UNCONNECTED__385, SYNOPSYS_UNCONNECTED__386, 
        SYNOPSYS_UNCONNECTED__387, SYNOPSYS_UNCONNECTED__388, 
        SYNOPSYS_UNCONNECTED__389, SYNOPSYS_UNCONNECTED__390, 
        SYNOPSYS_UNCONNECTED__391, SYNOPSYS_UNCONNECTED__392, 
        SYNOPSYS_UNCONNECTED__393, SYNOPSYS_UNCONNECTED__394, 
        SYNOPSYS_UNCONNECTED__395, SYNOPSYS_UNCONNECTED__396, 
        SYNOPSYS_UNCONNECTED__397, SYNOPSYS_UNCONNECTED__398, 
        SYNOPSYS_UNCONNECTED__399, SYNOPSYS_UNCONNECTED__400, 
        SYNOPSYS_UNCONNECTED__401, SYNOPSYS_UNCONNECTED__402, 
        SYNOPSYS_UNCONNECTED__403, SYNOPSYS_UNCONNECTED__404, 
        SYNOPSYS_UNCONNECTED__405, SYNOPSYS_UNCONNECTED__406, 
        SYNOPSYS_UNCONNECTED__407, SYNOPSYS_UNCONNECTED__408, 
        SYNOPSYS_UNCONNECTED__409, SYNOPSYS_UNCONNECTED__410, 
        SYNOPSYS_UNCONNECTED__411, SYNOPSYS_UNCONNECTED__412, 
        SYNOPSYS_UNCONNECTED__413, SYNOPSYS_UNCONNECTED__414, 
        SYNOPSYS_UNCONNECTED__415, N224, N223, N222, N221, N220, N219, N218, 
        N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193}) );
  matrixMult_N_M_1_N16_M32_DW01_add_26 add_54_I16_G3 ( .A(o[95:64]), .B({N160, 
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, 
        N135, N134, N133, N132, N131, N130, N129}), .CI(1'b0), .SUM({N192, 
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_13 mult_54_I16_G3 ( .A(x[511:480]), .B(
        y[7775:7744]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__416, 
        SYNOPSYS_UNCONNECTED__417, SYNOPSYS_UNCONNECTED__418, 
        SYNOPSYS_UNCONNECTED__419, SYNOPSYS_UNCONNECTED__420, 
        SYNOPSYS_UNCONNECTED__421, SYNOPSYS_UNCONNECTED__422, 
        SYNOPSYS_UNCONNECTED__423, SYNOPSYS_UNCONNECTED__424, 
        SYNOPSYS_UNCONNECTED__425, SYNOPSYS_UNCONNECTED__426, 
        SYNOPSYS_UNCONNECTED__427, SYNOPSYS_UNCONNECTED__428, 
        SYNOPSYS_UNCONNECTED__429, SYNOPSYS_UNCONNECTED__430, 
        SYNOPSYS_UNCONNECTED__431, SYNOPSYS_UNCONNECTED__432, 
        SYNOPSYS_UNCONNECTED__433, SYNOPSYS_UNCONNECTED__434, 
        SYNOPSYS_UNCONNECTED__435, SYNOPSYS_UNCONNECTED__436, 
        SYNOPSYS_UNCONNECTED__437, SYNOPSYS_UNCONNECTED__438, 
        SYNOPSYS_UNCONNECTED__439, SYNOPSYS_UNCONNECTED__440, 
        SYNOPSYS_UNCONNECTED__441, SYNOPSYS_UNCONNECTED__442, 
        SYNOPSYS_UNCONNECTED__443, SYNOPSYS_UNCONNECTED__444, 
        SYNOPSYS_UNCONNECTED__445, SYNOPSYS_UNCONNECTED__446, 
        SYNOPSYS_UNCONNECTED__447, N160, N159, N158, N157, N156, N155, N154, 
        N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, 
        N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, 
        N129}) );
  matrixMult_N_M_1_N16_M32_DW01_add_28 add_54_I16_G2 ( .A(o[63:32]), .B({N96, 
        N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, 
        N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, 
        N67, N66, N65}), .CI(1'b0), .SUM({N128, N127, N126, N125, N124, N123, 
        N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_14 mult_54_I16_G2 ( .A(x[511:480]), .B(
        y[7743:7712]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__448, 
        SYNOPSYS_UNCONNECTED__449, SYNOPSYS_UNCONNECTED__450, 
        SYNOPSYS_UNCONNECTED__451, SYNOPSYS_UNCONNECTED__452, 
        SYNOPSYS_UNCONNECTED__453, SYNOPSYS_UNCONNECTED__454, 
        SYNOPSYS_UNCONNECTED__455, SYNOPSYS_UNCONNECTED__456, 
        SYNOPSYS_UNCONNECTED__457, SYNOPSYS_UNCONNECTED__458, 
        SYNOPSYS_UNCONNECTED__459, SYNOPSYS_UNCONNECTED__460, 
        SYNOPSYS_UNCONNECTED__461, SYNOPSYS_UNCONNECTED__462, 
        SYNOPSYS_UNCONNECTED__463, SYNOPSYS_UNCONNECTED__464, 
        SYNOPSYS_UNCONNECTED__465, SYNOPSYS_UNCONNECTED__466, 
        SYNOPSYS_UNCONNECTED__467, SYNOPSYS_UNCONNECTED__468, 
        SYNOPSYS_UNCONNECTED__469, SYNOPSYS_UNCONNECTED__470, 
        SYNOPSYS_UNCONNECTED__471, SYNOPSYS_UNCONNECTED__472, 
        SYNOPSYS_UNCONNECTED__473, SYNOPSYS_UNCONNECTED__474, 
        SYNOPSYS_UNCONNECTED__475, SYNOPSYS_UNCONNECTED__476, 
        SYNOPSYS_UNCONNECTED__477, SYNOPSYS_UNCONNECTED__478, 
        SYNOPSYS_UNCONNECTED__479, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65}) );
  matrixMult_N_M_1_N16_M32_DW01_add_30 add_54_I16 ( .A(o[31:0]), .B({N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}), .CI(1'b0), .SUM({N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33}) );
  matrixMult_N_M_1_N16_M32_DW02_mult_15 mult_54_I16 ( .A(x[511:480]), .B(
        y[7711:7680]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__480, 
        SYNOPSYS_UNCONNECTED__481, SYNOPSYS_UNCONNECTED__482, 
        SYNOPSYS_UNCONNECTED__483, SYNOPSYS_UNCONNECTED__484, 
        SYNOPSYS_UNCONNECTED__485, SYNOPSYS_UNCONNECTED__486, 
        SYNOPSYS_UNCONNECTED__487, SYNOPSYS_UNCONNECTED__488, 
        SYNOPSYS_UNCONNECTED__489, SYNOPSYS_UNCONNECTED__490, 
        SYNOPSYS_UNCONNECTED__491, SYNOPSYS_UNCONNECTED__492, 
        SYNOPSYS_UNCONNECTED__493, SYNOPSYS_UNCONNECTED__494, 
        SYNOPSYS_UNCONNECTED__495, SYNOPSYS_UNCONNECTED__496, 
        SYNOPSYS_UNCONNECTED__497, SYNOPSYS_UNCONNECTED__498, 
        SYNOPSYS_UNCONNECTED__499, SYNOPSYS_UNCONNECTED__500, 
        SYNOPSYS_UNCONNECTED__501, SYNOPSYS_UNCONNECTED__502, 
        SYNOPSYS_UNCONNECTED__503, SYNOPSYS_UNCONNECTED__504, 
        SYNOPSYS_UNCONNECTED__505, SYNOPSYS_UNCONNECTED__506, 
        SYNOPSYS_UNCONNECTED__507, SYNOPSYS_UNCONNECTED__508, 
        SYNOPSYS_UNCONNECTED__509, SYNOPSYS_UNCONNECTED__510, 
        SYNOPSYS_UNCONNECTED__511, N32, N31, N30, N29, N28, N27, N26, N25, N24, 
        N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, 
        N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
endmodule

