
module stackMachine_N64 ( clk, rst, x, opcode, o );
  input [63:0] x;
  input [2:0] opcode;
  output [63:0] o;
  input clk, rst;
  wire   \stack[7][63] , \stack[7][62] , \stack[7][61] , \stack[7][60] ,
         \stack[7][59] , \stack[7][58] , \stack[7][57] , \stack[7][56] ,
         \stack[7][55] , \stack[7][54] , \stack[7][53] , \stack[7][52] ,
         \stack[7][51] , \stack[7][50] , \stack[7][49] , \stack[7][48] ,
         \stack[7][47] , \stack[7][46] , \stack[7][45] , \stack[7][44] ,
         \stack[7][43] , \stack[7][42] , \stack[7][41] , \stack[7][40] ,
         \stack[7][39] , \stack[7][38] , \stack[7][37] , \stack[7][36] ,
         \stack[7][35] , \stack[7][34] , \stack[7][33] , \stack[7][32] ,
         \stack[7][31] , \stack[7][30] , \stack[7][29] , \stack[7][28] ,
         \stack[7][27] , \stack[7][26] , \stack[7][25] , \stack[7][24] ,
         \stack[7][23] , \stack[7][22] , \stack[7][21] , \stack[7][20] ,
         \stack[7][19] , \stack[7][18] , \stack[7][17] , \stack[7][16] ,
         \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][63] , \stack[6][62] , \stack[6][61] , \stack[6][60] ,
         \stack[6][59] , \stack[6][58] , \stack[6][57] , \stack[6][56] ,
         \stack[6][55] , \stack[6][54] , \stack[6][53] , \stack[6][52] ,
         \stack[6][51] , \stack[6][50] , \stack[6][49] , \stack[6][48] ,
         \stack[6][47] , \stack[6][46] , \stack[6][45] , \stack[6][44] ,
         \stack[6][43] , \stack[6][42] , \stack[6][41] , \stack[6][40] ,
         \stack[6][39] , \stack[6][38] , \stack[6][37] , \stack[6][36] ,
         \stack[6][35] , \stack[6][34] , \stack[6][33] , \stack[6][32] ,
         \stack[6][31] , \stack[6][30] , \stack[6][29] , \stack[6][28] ,
         \stack[6][27] , \stack[6][26] , \stack[6][25] , \stack[6][24] ,
         \stack[6][23] , \stack[6][22] , \stack[6][21] , \stack[6][20] ,
         \stack[6][19] , \stack[6][18] , \stack[6][17] , \stack[6][16] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][63] , \stack[5][62] , \stack[5][61] , \stack[5][60] ,
         \stack[5][59] , \stack[5][58] , \stack[5][57] , \stack[5][56] ,
         \stack[5][55] , \stack[5][54] , \stack[5][53] , \stack[5][52] ,
         \stack[5][51] , \stack[5][50] , \stack[5][49] , \stack[5][48] ,
         \stack[5][47] , \stack[5][46] , \stack[5][45] , \stack[5][44] ,
         \stack[5][43] , \stack[5][42] , \stack[5][41] , \stack[5][40] ,
         \stack[5][39] , \stack[5][38] , \stack[5][37] , \stack[5][36] ,
         \stack[5][35] , \stack[5][34] , \stack[5][33] , \stack[5][32] ,
         \stack[5][31] , \stack[5][30] , \stack[5][29] , \stack[5][28] ,
         \stack[5][27] , \stack[5][26] , \stack[5][25] , \stack[5][24] ,
         \stack[5][23] , \stack[5][22] , \stack[5][21] , \stack[5][20] ,
         \stack[5][19] , \stack[5][18] , \stack[5][17] , \stack[5][16] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][63] , \stack[4][62] , \stack[4][61] , \stack[4][60] ,
         \stack[4][59] , \stack[4][58] , \stack[4][57] , \stack[4][56] ,
         \stack[4][55] , \stack[4][54] , \stack[4][53] , \stack[4][52] ,
         \stack[4][51] , \stack[4][50] , \stack[4][49] , \stack[4][48] ,
         \stack[4][47] , \stack[4][46] , \stack[4][45] , \stack[4][44] ,
         \stack[4][43] , \stack[4][42] , \stack[4][41] , \stack[4][40] ,
         \stack[4][39] , \stack[4][38] , \stack[4][37] , \stack[4][36] ,
         \stack[4][35] , \stack[4][34] , \stack[4][33] , \stack[4][32] ,
         \stack[4][31] , \stack[4][30] , \stack[4][29] , \stack[4][28] ,
         \stack[4][27] , \stack[4][26] , \stack[4][25] , \stack[4][24] ,
         \stack[4][23] , \stack[4][22] , \stack[4][21] , \stack[4][20] ,
         \stack[4][19] , \stack[4][18] , \stack[4][17] , \stack[4][16] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][63] , \stack[3][62] , \stack[3][61] , \stack[3][60] ,
         \stack[3][59] , \stack[3][58] , \stack[3][57] , \stack[3][56] ,
         \stack[3][55] , \stack[3][54] , \stack[3][53] , \stack[3][52] ,
         \stack[3][51] , \stack[3][50] , \stack[3][49] , \stack[3][48] ,
         \stack[3][47] , \stack[3][46] , \stack[3][45] , \stack[3][44] ,
         \stack[3][43] , \stack[3][42] , \stack[3][41] , \stack[3][40] ,
         \stack[3][39] , \stack[3][38] , \stack[3][37] , \stack[3][36] ,
         \stack[3][35] , \stack[3][34] , \stack[3][33] , \stack[3][32] ,
         \stack[3][31] , \stack[3][30] , \stack[3][29] , \stack[3][28] ,
         \stack[3][27] , \stack[3][26] , \stack[3][25] , \stack[3][24] ,
         \stack[3][23] , \stack[3][22] , \stack[3][21] , \stack[3][20] ,
         \stack[3][19] , \stack[3][18] , \stack[3][17] , \stack[3][16] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][63] , \stack[2][62] , \stack[2][61] , \stack[2][60] ,
         \stack[2][59] , \stack[2][58] , \stack[2][57] , \stack[2][56] ,
         \stack[2][55] , \stack[2][54] , \stack[2][53] , \stack[2][52] ,
         \stack[2][51] , \stack[2][50] , \stack[2][49] , \stack[2][48] ,
         \stack[2][47] , \stack[2][46] , \stack[2][45] , \stack[2][44] ,
         \stack[2][43] , \stack[2][42] , \stack[2][41] , \stack[2][40] ,
         \stack[2][39] , \stack[2][38] , \stack[2][37] , \stack[2][36] ,
         \stack[2][35] , \stack[2][34] , \stack[2][33] , \stack[2][32] ,
         \stack[2][31] , \stack[2][30] , \stack[2][29] , \stack[2][28] ,
         \stack[2][27] , \stack[2][26] , \stack[2][25] , \stack[2][24] ,
         \stack[2][23] , \stack[2][22] , \stack[2][21] , \stack[2][20] ,
         \stack[2][19] , \stack[2][18] , \stack[2][17] , \stack[2][16] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][63] , \stack[1][62] , \stack[1][61] , \stack[1][60] ,
         \stack[1][59] , \stack[1][58] , \stack[1][57] , \stack[1][56] ,
         \stack[1][55] , \stack[1][54] , \stack[1][53] , \stack[1][52] ,
         \stack[1][51] , \stack[1][50] , \stack[1][49] , \stack[1][48] ,
         \stack[1][47] , \stack[1][46] , \stack[1][45] , \stack[1][44] ,
         \stack[1][43] , \stack[1][42] , \stack[1][41] , \stack[1][40] ,
         \stack[1][39] , \stack[1][38] , \stack[1][37] , \stack[1][36] ,
         \stack[1][35] , \stack[1][34] , \stack[1][33] , \stack[1][32] ,
         \stack[1][31] , \stack[1][30] , \stack[1][29] , \stack[1][28] ,
         \stack[1][27] , \stack[1][26] , \stack[1][25] , \stack[1][24] ,
         \stack[1][23] , \stack[1][22] , \stack[1][21] , \stack[1][20] ,
         \stack[1][19] , \stack[1][18] , \stack[1][17] , \stack[1][16] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \C3/DATA5_0 , \C3/DATA5_1 , \C3/DATA5_2 , \C3/DATA5_3 , \C3/DATA5_4 ,
         \C3/DATA5_5 , \C3/DATA5_6 , \C3/DATA5_7 , \C3/DATA5_8 , \C3/DATA5_9 ,
         \C3/DATA5_10 , \C3/DATA5_11 , \C3/DATA5_12 , \C3/DATA5_13 ,
         \C3/DATA5_14 , \C3/DATA5_15 , \C3/DATA5_16 , \C3/DATA5_17 ,
         \C3/DATA5_18 , \C3/DATA5_19 , \C3/DATA5_20 , \C3/DATA5_21 ,
         \C3/DATA5_22 , \C3/DATA5_23 , \C3/DATA5_24 , \C3/DATA5_25 ,
         \C3/DATA5_26 , \C3/DATA5_27 , \C3/DATA5_28 , \C3/DATA5_29 ,
         \C3/DATA5_30 , \C3/DATA5_31 , \C3/DATA5_32 , \C3/DATA5_33 ,
         \C3/DATA5_34 , \C3/DATA5_35 , \C3/DATA5_36 , \C3/DATA5_37 ,
         \C3/DATA5_38 , \C3/DATA5_39 , \C3/DATA5_40 , \C3/DATA5_41 ,
         \C3/DATA5_42 , \C3/DATA5_43 , \C3/DATA5_44 , \C3/DATA5_45 ,
         \C3/DATA5_46 , \C3/DATA5_47 , \C3/DATA5_48 , \C3/DATA5_49 ,
         \C3/DATA5_50 , \C3/DATA5_51 , \C3/DATA5_52 , \C3/DATA5_53 ,
         \C3/DATA5_54 , \C3/DATA5_55 , \C3/DATA5_56 , \C3/DATA5_57 ,
         \C3/DATA5_58 , \C3/DATA5_59 , \C3/DATA5_60 , \C3/DATA5_61 ,
         \C3/DATA5_62 , \C3/DATA5_63 , n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, \C1/Z_0 ,
         \U1/RSOP_16/C3/Z_63 , \U1/RSOP_16/C3/Z_62 , \U1/RSOP_16/C3/Z_61 ,
         \U1/RSOP_16/C3/Z_60 , \U1/RSOP_16/C3/Z_59 , \U1/RSOP_16/C3/Z_58 ,
         \U1/RSOP_16/C3/Z_57 , \U1/RSOP_16/C3/Z_56 , \U1/RSOP_16/C3/Z_55 ,
         \U1/RSOP_16/C3/Z_54 , \U1/RSOP_16/C3/Z_53 , \U1/RSOP_16/C3/Z_52 ,
         \U1/RSOP_16/C3/Z_51 , \U1/RSOP_16/C3/Z_50 , \U1/RSOP_16/C3/Z_49 ,
         \U1/RSOP_16/C3/Z_48 , \U1/RSOP_16/C3/Z_47 , \U1/RSOP_16/C3/Z_46 ,
         \U1/RSOP_16/C3/Z_45 , \U1/RSOP_16/C3/Z_44 , \U1/RSOP_16/C3/Z_43 ,
         \U1/RSOP_16/C3/Z_42 , \U1/RSOP_16/C3/Z_41 , \U1/RSOP_16/C3/Z_40 ,
         \U1/RSOP_16/C3/Z_39 , \U1/RSOP_16/C3/Z_38 , \U1/RSOP_16/C3/Z_37 ,
         \U1/RSOP_16/C3/Z_36 , \U1/RSOP_16/C3/Z_35 , \U1/RSOP_16/C3/Z_34 ,
         \U1/RSOP_16/C3/Z_33 , \U1/RSOP_16/C3/Z_32 , \U1/RSOP_16/C3/Z_31 ,
         \U1/RSOP_16/C3/Z_30 , \U1/RSOP_16/C3/Z_29 , \U1/RSOP_16/C3/Z_28 ,
         \U1/RSOP_16/C3/Z_27 , \U1/RSOP_16/C3/Z_26 , \U1/RSOP_16/C3/Z_25 ,
         \U1/RSOP_16/C3/Z_24 , \U1/RSOP_16/C3/Z_23 , \U1/RSOP_16/C3/Z_22 ,
         \U1/RSOP_16/C3/Z_21 , \U1/RSOP_16/C3/Z_20 , \U1/RSOP_16/C3/Z_19 ,
         \U1/RSOP_16/C3/Z_18 , \U1/RSOP_16/C3/Z_17 , \U1/RSOP_16/C3/Z_16 ,
         \U1/RSOP_16/C3/Z_15 , \U1/RSOP_16/C3/Z_14 , \U1/RSOP_16/C3/Z_13 ,
         \U1/RSOP_16/C3/Z_12 , \U1/RSOP_16/C3/Z_11 , \U1/RSOP_16/C3/Z_10 ,
         \U1/RSOP_16/C3/Z_9 , \U1/RSOP_16/C3/Z_8 , \U1/RSOP_16/C3/Z_7 ,
         \U1/RSOP_16/C3/Z_6 , \U1/RSOP_16/C3/Z_5 , \U1/RSOP_16/C3/Z_4 ,
         \U1/RSOP_16/C3/Z_3 , \U1/RSOP_16/C3/Z_2 , \U1/RSOP_16/C3/Z_1 ,
         \U1/RSOP_16/C3/Z_0 , \U1/RSOP_16/C2/Z_63 , \U1/RSOP_16/C2/Z_62 ,
         \U1/RSOP_16/C2/Z_61 , \U1/RSOP_16/C2/Z_60 , \U1/RSOP_16/C2/Z_59 ,
         \U1/RSOP_16/C2/Z_58 , \U1/RSOP_16/C2/Z_57 , \U1/RSOP_16/C2/Z_56 ,
         \U1/RSOP_16/C2/Z_55 , \U1/RSOP_16/C2/Z_54 , \U1/RSOP_16/C2/Z_53 ,
         \U1/RSOP_16/C2/Z_52 , \U1/RSOP_16/C2/Z_51 , \U1/RSOP_16/C2/Z_50 ,
         \U1/RSOP_16/C2/Z_49 , \U1/RSOP_16/C2/Z_48 , \U1/RSOP_16/C2/Z_47 ,
         \U1/RSOP_16/C2/Z_46 , \U1/RSOP_16/C2/Z_45 , \U1/RSOP_16/C2/Z_44 ,
         \U1/RSOP_16/C2/Z_43 , \U1/RSOP_16/C2/Z_42 , \U1/RSOP_16/C2/Z_41 ,
         \U1/RSOP_16/C2/Z_40 , \U1/RSOP_16/C2/Z_39 , \U1/RSOP_16/C2/Z_38 ,
         \U1/RSOP_16/C2/Z_37 , \U1/RSOP_16/C2/Z_36 , \U1/RSOP_16/C2/Z_35 ,
         \U1/RSOP_16/C2/Z_34 , \U1/RSOP_16/C2/Z_33 , \U1/RSOP_16/C2/Z_32 ,
         \U1/RSOP_16/C2/Z_31 , \U1/RSOP_16/C2/Z_30 , \U1/RSOP_16/C2/Z_29 ,
         \U1/RSOP_16/C2/Z_28 , \U1/RSOP_16/C2/Z_27 , \U1/RSOP_16/C2/Z_26 ,
         \U1/RSOP_16/C2/Z_25 , \U1/RSOP_16/C2/Z_24 , \U1/RSOP_16/C2/Z_23 ,
         \U1/RSOP_16/C2/Z_22 , \U1/RSOP_16/C2/Z_21 , \U1/RSOP_16/C2/Z_20 ,
         \U1/RSOP_16/C2/Z_19 , \U1/RSOP_16/C2/Z_18 , \U1/RSOP_16/C2/Z_17 ,
         \U1/RSOP_16/C2/Z_16 , \U1/RSOP_16/C2/Z_15 , \U1/RSOP_16/C2/Z_14 ,
         \U1/RSOP_16/C2/Z_13 , \U1/RSOP_16/C2/Z_12 , \U1/RSOP_16/C2/Z_11 ,
         \U1/RSOP_16/C2/Z_10 , \U1/RSOP_16/C2/Z_9 , \U1/RSOP_16/C2/Z_8 ,
         \U1/RSOP_16/C2/Z_7 , \U1/RSOP_16/C2/Z_6 , \U1/RSOP_16/C2/Z_5 ,
         \U1/RSOP_16/C2/Z_4 , \U1/RSOP_16/C2/Z_3 , \U1/RSOP_16/C2/Z_2 ,
         \U1/RSOP_16/C2/Z_1 , \U1/RSOP_16/C2/Z_0 , \DP_OP_25_64_8855/n656 ,
         \DP_OP_25_64_8855/n655 , \DP_OP_25_64_8855/n654 ,
         \DP_OP_25_64_8855/n653 , \DP_OP_25_64_8855/n652 ,
         \DP_OP_25_64_8855/n651 , \DP_OP_25_64_8855/n650 ,
         \DP_OP_25_64_8855/n649 , \DP_OP_25_64_8855/n648 ,
         \DP_OP_25_64_8855/n647 , \DP_OP_25_64_8855/n646 ,
         \DP_OP_25_64_8855/n645 , \DP_OP_25_64_8855/n644 ,
         \DP_OP_25_64_8855/n643 , \DP_OP_25_64_8855/n642 ,
         \DP_OP_25_64_8855/n641 , \DP_OP_25_64_8855/n640 ,
         \DP_OP_25_64_8855/n639 , \DP_OP_25_64_8855/n638 ,
         \DP_OP_25_64_8855/n637 , \DP_OP_25_64_8855/n636 ,
         \DP_OP_25_64_8855/n635 , \DP_OP_25_64_8855/n634 ,
         \DP_OP_25_64_8855/n633 , \DP_OP_25_64_8855/n632 ,
         \DP_OP_25_64_8855/n631 , \DP_OP_25_64_8855/n630 ,
         \DP_OP_25_64_8855/n629 , \DP_OP_25_64_8855/n628 ,
         \DP_OP_25_64_8855/n627 , \DP_OP_25_64_8855/n626 ,
         \DP_OP_25_64_8855/n625 , \DP_OP_25_64_8855/n624 ,
         \DP_OP_25_64_8855/n623 , \DP_OP_25_64_8855/n622 ,
         \DP_OP_25_64_8855/n621 , \DP_OP_25_64_8855/n620 ,
         \DP_OP_25_64_8855/n619 , \DP_OP_25_64_8855/n618 ,
         \DP_OP_25_64_8855/n617 , \DP_OP_25_64_8855/n616 ,
         \DP_OP_25_64_8855/n615 , \DP_OP_25_64_8855/n614 ,
         \DP_OP_25_64_8855/n613 , \DP_OP_25_64_8855/n612 ,
         \DP_OP_25_64_8855/n611 , \DP_OP_25_64_8855/n610 ,
         \DP_OP_25_64_8855/n609 , \DP_OP_25_64_8855/n608 ,
         \DP_OP_25_64_8855/n607 , \DP_OP_25_64_8855/n606 ,
         \DP_OP_25_64_8855/n605 , \DP_OP_25_64_8855/n604 ,
         \DP_OP_25_64_8855/n603 , \DP_OP_25_64_8855/n602 ,
         \DP_OP_25_64_8855/n601 , \DP_OP_25_64_8855/n600 ,
         \DP_OP_25_64_8855/n599 , \DP_OP_25_64_8855/n598 ,
         \DP_OP_25_64_8855/n597 , \DP_OP_25_64_8855/n596 ,
         \DP_OP_25_64_8855/n595 , \DP_OP_25_64_8855/n594 ,
         \DP_OP_25_64_8855/n593 , \DP_OP_25_64_8855/n588 ,
         \DP_OP_25_64_8855/n587 , \DP_OP_25_64_8855/n586 ,
         \DP_OP_25_64_8855/n585 , \DP_OP_25_64_8855/n584 ,
         \DP_OP_25_64_8855/n583 , \DP_OP_25_64_8855/n582 ,
         \DP_OP_25_64_8855/n581 , \DP_OP_25_64_8855/n580 ,
         \DP_OP_25_64_8855/n579 , \DP_OP_25_64_8855/n578 ,
         \DP_OP_25_64_8855/n577 , \DP_OP_25_64_8855/n576 ,
         \DP_OP_25_64_8855/n575 , \DP_OP_25_64_8855/n574 ,
         \DP_OP_25_64_8855/n573 , \DP_OP_25_64_8855/n572 ,
         \DP_OP_25_64_8855/n571 , \DP_OP_25_64_8855/n570 ,
         \DP_OP_25_64_8855/n569 , \DP_OP_25_64_8855/n568 ,
         \DP_OP_25_64_8855/n567 , \DP_OP_25_64_8855/n566 ,
         \DP_OP_25_64_8855/n565 , \DP_OP_25_64_8855/n564 ,
         \DP_OP_25_64_8855/n563 , \DP_OP_25_64_8855/n562 ,
         \DP_OP_25_64_8855/n561 , \DP_OP_25_64_8855/n560 ,
         \DP_OP_25_64_8855/n559 , \DP_OP_25_64_8855/n558 ,
         \DP_OP_25_64_8855/n557 , \DP_OP_25_64_8855/n556 ,
         \DP_OP_25_64_8855/n555 , \DP_OP_25_64_8855/n554 ,
         \DP_OP_25_64_8855/n553 , \DP_OP_25_64_8855/n552 ,
         \DP_OP_25_64_8855/n551 , \DP_OP_25_64_8855/n550 ,
         \DP_OP_25_64_8855/n549 , \DP_OP_25_64_8855/n548 ,
         \DP_OP_25_64_8855/n547 , \DP_OP_25_64_8855/n546 ,
         \DP_OP_25_64_8855/n545 , \DP_OP_25_64_8855/n544 ,
         \DP_OP_25_64_8855/n543 , \DP_OP_25_64_8855/n542 ,
         \DP_OP_25_64_8855/n541 , \DP_OP_25_64_8855/n540 ,
         \DP_OP_25_64_8855/n539 , \DP_OP_25_64_8855/n538 ,
         \DP_OP_25_64_8855/n537 , \DP_OP_25_64_8855/n536 ,
         \DP_OP_25_64_8855/n535 , \DP_OP_25_64_8855/n534 ,
         \DP_OP_25_64_8855/n533 , \DP_OP_25_64_8855/n532 ,
         \DP_OP_25_64_8855/n531 , \DP_OP_25_64_8855/n530 ,
         \DP_OP_25_64_8855/n529 , \DP_OP_25_64_8855/n528 ,
         \DP_OP_25_64_8855/n527 , \DP_OP_25_64_8855/n526 ,
         \DP_OP_25_64_8855/n525 , \DP_OP_25_64_8855/n524 ,
         \DP_OP_25_64_8855/n523 , \DP_OP_25_64_8855/n522 ,
         \DP_OP_25_64_8855/n521 , \DP_OP_25_64_8855/n520 ,
         \DP_OP_25_64_8855/n519 , \DP_OP_25_64_8855/n518 ,
         \DP_OP_25_64_8855/n517 , \DP_OP_25_64_8855/n516 ,
         \DP_OP_25_64_8855/n515 , \DP_OP_25_64_8855/n514 ,
         \DP_OP_25_64_8855/n513 , \DP_OP_25_64_8855/n512 ,
         \DP_OP_25_64_8855/n511 , \DP_OP_25_64_8855/n510 ,
         \DP_OP_25_64_8855/n509 , \DP_OP_25_64_8855/n508 ,
         \DP_OP_25_64_8855/n507 , \DP_OP_25_64_8855/n506 ,
         \DP_OP_25_64_8855/n505 , \DP_OP_25_64_8855/n504 ,
         \DP_OP_25_64_8855/n503 , \DP_OP_25_64_8855/n502 ,
         \DP_OP_25_64_8855/n501 , \DP_OP_25_64_8855/n500 ,
         \DP_OP_25_64_8855/n499 , \DP_OP_25_64_8855/n498 ,
         \DP_OP_25_64_8855/n497 , \DP_OP_25_64_8855/n496 ,
         \DP_OP_25_64_8855/n495 , \DP_OP_25_64_8855/n494 ,
         \DP_OP_25_64_8855/n493 , \DP_OP_25_64_8855/n492 ,
         \DP_OP_25_64_8855/n491 , \DP_OP_25_64_8855/n490 ,
         \DP_OP_25_64_8855/n489 , \DP_OP_25_64_8855/n488 ,
         \DP_OP_25_64_8855/n487 , \DP_OP_25_64_8855/n486 ,
         \DP_OP_25_64_8855/n485 , \DP_OP_25_64_8855/n484 ,
         \DP_OP_25_64_8855/n483 , \DP_OP_25_64_8855/n482 ,
         \DP_OP_25_64_8855/n481 , \DP_OP_25_64_8855/n480 ,
         \DP_OP_25_64_8855/n479 , \DP_OP_25_64_8855/n478 ,
         \DP_OP_25_64_8855/n477 , \DP_OP_25_64_8855/n476 ,
         \DP_OP_25_64_8855/n475 , \DP_OP_25_64_8855/n474 ,
         \DP_OP_25_64_8855/n473 , \DP_OP_25_64_8855/n472 ,
         \DP_OP_25_64_8855/n471 , \DP_OP_25_64_8855/n470 ,
         \DP_OP_25_64_8855/n469 , \DP_OP_25_64_8855/n468 ,
         \DP_OP_25_64_8855/n467 , \DP_OP_25_64_8855/n466 ,
         \DP_OP_25_64_8855/n465 , \DP_OP_25_64_8855/n464 ,
         \DP_OP_25_64_8855/n463 , \DP_OP_25_64_8855/n462 ,
         \DP_OP_25_64_8855/n460 , \DP_OP_25_64_8855/n459 ,
         \DP_OP_25_64_8855/n453 , \DP_OP_25_64_8855/n452 ,
         \DP_OP_25_64_8855/n446 , \DP_OP_25_64_8855/n445 ,
         \DP_OP_25_64_8855/n439 , \DP_OP_25_64_8855/n438 ,
         \DP_OP_25_64_8855/n432 , \DP_OP_25_64_8855/n431 ,
         \DP_OP_25_64_8855/n425 , \DP_OP_25_64_8855/n424 ,
         \DP_OP_25_64_8855/n418 , \DP_OP_25_64_8855/n417 ,
         \DP_OP_25_64_8855/n411 , \DP_OP_25_64_8855/n410 ,
         \DP_OP_25_64_8855/n404 , \DP_OP_25_64_8855/n403 ,
         \DP_OP_25_64_8855/n397 , \DP_OP_25_64_8855/n396 ,
         \DP_OP_25_64_8855/n390 , \DP_OP_25_64_8855/n389 ,
         \DP_OP_25_64_8855/n383 , \DP_OP_25_64_8855/n382 ,
         \DP_OP_25_64_8855/n376 , \DP_OP_25_64_8855/n375 ,
         \DP_OP_25_64_8855/n369 , \DP_OP_25_64_8855/n368 ,
         \DP_OP_25_64_8855/n362 , \DP_OP_25_64_8855/n361 ,
         \DP_OP_25_64_8855/n355 , \DP_OP_25_64_8855/n354 ,
         \DP_OP_25_64_8855/n348 , \DP_OP_25_64_8855/n347 ,
         \DP_OP_25_64_8855/n341 , \DP_OP_25_64_8855/n340 ,
         \DP_OP_25_64_8855/n334 , \DP_OP_25_64_8855/n333 ,
         \DP_OP_25_64_8855/n327 , \DP_OP_25_64_8855/n326 ,
         \DP_OP_25_64_8855/n320 , \DP_OP_25_64_8855/n319 ,
         \DP_OP_25_64_8855/n313 , \DP_OP_25_64_8855/n312 ,
         \DP_OP_25_64_8855/n306 , \DP_OP_25_64_8855/n305 ,
         \DP_OP_25_64_8855/n299 , \DP_OP_25_64_8855/n298 ,
         \DP_OP_25_64_8855/n292 , \DP_OP_25_64_8855/n291 ,
         \DP_OP_25_64_8855/n285 , \DP_OP_25_64_8855/n284 ,
         \DP_OP_25_64_8855/n278 , \DP_OP_25_64_8855/n277 ,
         \DP_OP_25_64_8855/n271 , \DP_OP_25_64_8855/n270 ,
         \DP_OP_25_64_8855/n264 , \DP_OP_25_64_8855/n263 ,
         \DP_OP_25_64_8855/n257 , \DP_OP_25_64_8855/n256 ,
         \DP_OP_25_64_8855/n250 , \DP_OP_25_64_8855/n249 ,
         \DP_OP_25_64_8855/n243 , \DP_OP_25_64_8855/n242 ,
         \DP_OP_25_64_8855/n236 , \DP_OP_25_64_8855/n235 ,
         \DP_OP_25_64_8855/n229 , \DP_OP_25_64_8855/n228 ,
         \DP_OP_25_64_8855/n222 , \DP_OP_25_64_8855/n221 ,
         \DP_OP_25_64_8855/n215 , \DP_OP_25_64_8855/n214 ,
         \DP_OP_25_64_8855/n208 , \DP_OP_25_64_8855/n207 ,
         \DP_OP_25_64_8855/n201 , \DP_OP_25_64_8855/n200 ,
         \DP_OP_25_64_8855/n194 , \DP_OP_25_64_8855/n193 ,
         \DP_OP_25_64_8855/n187 , \DP_OP_25_64_8855/n186 ,
         \DP_OP_25_64_8855/n180 , \DP_OP_25_64_8855/n179 ,
         \DP_OP_25_64_8855/n173 , \DP_OP_25_64_8855/n172 ,
         \DP_OP_25_64_8855/n166 , \DP_OP_25_64_8855/n165 ,
         \DP_OP_25_64_8855/n159 , \DP_OP_25_64_8855/n158 ,
         \DP_OP_25_64_8855/n152 , \DP_OP_25_64_8855/n151 ,
         \DP_OP_25_64_8855/n145 , \DP_OP_25_64_8855/n144 ,
         \DP_OP_25_64_8855/n138 , \DP_OP_25_64_8855/n137 ,
         \DP_OP_25_64_8855/n131 , \DP_OP_25_64_8855/n130 ,
         \DP_OP_25_64_8855/n124 , \DP_OP_25_64_8855/n123 ,
         \DP_OP_25_64_8855/n117 , \DP_OP_25_64_8855/n116 ,
         \DP_OP_25_64_8855/n110 , \DP_OP_25_64_8855/n109 ,
         \DP_OP_25_64_8855/n103 , \DP_OP_25_64_8855/n102 ,
         \DP_OP_25_64_8855/n96 , \DP_OP_25_64_8855/n95 ,
         \DP_OP_25_64_8855/n89 , \DP_OP_25_64_8855/n88 ,
         \DP_OP_25_64_8855/n82 , \DP_OP_25_64_8855/n81 ,
         \DP_OP_25_64_8855/n57 , \DP_OP_25_64_8855/n56 ,
         \DP_OP_25_64_8855/n50 , \DP_OP_25_64_8855/n49 ,
         \DP_OP_25_64_8855/n43 , \DP_OP_25_64_8855/n42 ,
         \DP_OP_25_64_8855/n36 , \DP_OP_25_64_8855/n35 ,
         \DP_OP_25_64_8855/n29 , \DP_OP_25_64_8855/n28 ,
         \DP_OP_25_64_8855/n22 , \DP_OP_25_64_8855/n21 ,
         \DP_OP_25_64_8855/n15 , \DP_OP_25_64_8855/n14 , \DP_OP_25_64_8855/n8 ,
         \DP_OP_25_64_8855/n5 , n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489;

  DFF \stack_reg[0][0]  ( .D(n2632), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \stack_reg[1][0]  ( .D(n2631), .CLK(clk), .RST(rst), .Q(\stack[1][0] )
         );
  DFF \stack_reg[0][1]  ( .D(n2630), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \stack_reg[1][1]  ( .D(n2629), .CLK(clk), .RST(rst), .Q(\stack[1][1] )
         );
  DFF \stack_reg[2][1]  ( .D(n2628), .CLK(clk), .RST(rst), .Q(\stack[2][1] )
         );
  DFF \stack_reg[3][1]  ( .D(n2627), .CLK(clk), .RST(rst), .Q(\stack[3][1] )
         );
  DFF \stack_reg[4][1]  ( .D(n2626), .CLK(clk), .RST(rst), .Q(\stack[4][1] )
         );
  DFF \stack_reg[5][1]  ( .D(n2625), .CLK(clk), .RST(rst), .Q(\stack[5][1] )
         );
  DFF \stack_reg[6][1]  ( .D(n2624), .CLK(clk), .RST(rst), .Q(\stack[6][1] )
         );
  DFF \stack_reg[7][1]  ( .D(n2623), .CLK(clk), .RST(rst), .Q(\stack[7][1] )
         );
  DFF \stack_reg[0][2]  ( .D(n2622), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \stack_reg[1][2]  ( .D(n2621), .CLK(clk), .RST(rst), .Q(\stack[1][2] )
         );
  DFF \stack_reg[2][2]  ( .D(n2620), .CLK(clk), .RST(rst), .Q(\stack[2][2] )
         );
  DFF \stack_reg[3][2]  ( .D(n2619), .CLK(clk), .RST(rst), .Q(\stack[3][2] )
         );
  DFF \stack_reg[4][2]  ( .D(n2618), .CLK(clk), .RST(rst), .Q(\stack[4][2] )
         );
  DFF \stack_reg[5][2]  ( .D(n2617), .CLK(clk), .RST(rst), .Q(\stack[5][2] )
         );
  DFF \stack_reg[6][2]  ( .D(n2616), .CLK(clk), .RST(rst), .Q(\stack[6][2] )
         );
  DFF \stack_reg[7][2]  ( .D(n2615), .CLK(clk), .RST(rst), .Q(\stack[7][2] )
         );
  DFF \stack_reg[0][3]  ( .D(n2614), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \stack_reg[1][3]  ( .D(n2613), .CLK(clk), .RST(rst), .Q(\stack[1][3] )
         );
  DFF \stack_reg[2][3]  ( .D(n2612), .CLK(clk), .RST(rst), .Q(\stack[2][3] )
         );
  DFF \stack_reg[3][3]  ( .D(n2611), .CLK(clk), .RST(rst), .Q(\stack[3][3] )
         );
  DFF \stack_reg[4][3]  ( .D(n2610), .CLK(clk), .RST(rst), .Q(\stack[4][3] )
         );
  DFF \stack_reg[5][3]  ( .D(n2609), .CLK(clk), .RST(rst), .Q(\stack[5][3] )
         );
  DFF \stack_reg[6][3]  ( .D(n2608), .CLK(clk), .RST(rst), .Q(\stack[6][3] )
         );
  DFF \stack_reg[7][3]  ( .D(n2607), .CLK(clk), .RST(rst), .Q(\stack[7][3] )
         );
  DFF \stack_reg[0][4]  ( .D(n2606), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \stack_reg[1][4]  ( .D(n2605), .CLK(clk), .RST(rst), .Q(\stack[1][4] )
         );
  DFF \stack_reg[2][4]  ( .D(n2604), .CLK(clk), .RST(rst), .Q(\stack[2][4] )
         );
  DFF \stack_reg[3][4]  ( .D(n2603), .CLK(clk), .RST(rst), .Q(\stack[3][4] )
         );
  DFF \stack_reg[4][4]  ( .D(n2602), .CLK(clk), .RST(rst), .Q(\stack[4][4] )
         );
  DFF \stack_reg[5][4]  ( .D(n2601), .CLK(clk), .RST(rst), .Q(\stack[5][4] )
         );
  DFF \stack_reg[6][4]  ( .D(n2600), .CLK(clk), .RST(rst), .Q(\stack[6][4] )
         );
  DFF \stack_reg[7][4]  ( .D(n2599), .CLK(clk), .RST(rst), .Q(\stack[7][4] )
         );
  DFF \stack_reg[0][5]  ( .D(n2598), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \stack_reg[1][5]  ( .D(n2597), .CLK(clk), .RST(rst), .Q(\stack[1][5] )
         );
  DFF \stack_reg[2][5]  ( .D(n2596), .CLK(clk), .RST(rst), .Q(\stack[2][5] )
         );
  DFF \stack_reg[3][5]  ( .D(n2595), .CLK(clk), .RST(rst), .Q(\stack[3][5] )
         );
  DFF \stack_reg[4][5]  ( .D(n2594), .CLK(clk), .RST(rst), .Q(\stack[4][5] )
         );
  DFF \stack_reg[5][5]  ( .D(n2593), .CLK(clk), .RST(rst), .Q(\stack[5][5] )
         );
  DFF \stack_reg[6][5]  ( .D(n2592), .CLK(clk), .RST(rst), .Q(\stack[6][5] )
         );
  DFF \stack_reg[7][5]  ( .D(n2591), .CLK(clk), .RST(rst), .Q(\stack[7][5] )
         );
  DFF \stack_reg[0][6]  ( .D(n2590), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \stack_reg[1][6]  ( .D(n2589), .CLK(clk), .RST(rst), .Q(\stack[1][6] )
         );
  DFF \stack_reg[2][6]  ( .D(n2588), .CLK(clk), .RST(rst), .Q(\stack[2][6] )
         );
  DFF \stack_reg[3][6]  ( .D(n2587), .CLK(clk), .RST(rst), .Q(\stack[3][6] )
         );
  DFF \stack_reg[4][6]  ( .D(n2586), .CLK(clk), .RST(rst), .Q(\stack[4][6] )
         );
  DFF \stack_reg[5][6]  ( .D(n2585), .CLK(clk), .RST(rst), .Q(\stack[5][6] )
         );
  DFF \stack_reg[6][6]  ( .D(n2584), .CLK(clk), .RST(rst), .Q(\stack[6][6] )
         );
  DFF \stack_reg[7][6]  ( .D(n2583), .CLK(clk), .RST(rst), .Q(\stack[7][6] )
         );
  DFF \stack_reg[0][7]  ( .D(n2582), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \stack_reg[1][7]  ( .D(n2581), .CLK(clk), .RST(rst), .Q(\stack[1][7] )
         );
  DFF \stack_reg[2][7]  ( .D(n2580), .CLK(clk), .RST(rst), .Q(\stack[2][7] )
         );
  DFF \stack_reg[3][7]  ( .D(n2579), .CLK(clk), .RST(rst), .Q(\stack[3][7] )
         );
  DFF \stack_reg[4][7]  ( .D(n2578), .CLK(clk), .RST(rst), .Q(\stack[4][7] )
         );
  DFF \stack_reg[5][7]  ( .D(n2577), .CLK(clk), .RST(rst), .Q(\stack[5][7] )
         );
  DFF \stack_reg[6][7]  ( .D(n2576), .CLK(clk), .RST(rst), .Q(\stack[6][7] )
         );
  DFF \stack_reg[7][7]  ( .D(n2575), .CLK(clk), .RST(rst), .Q(\stack[7][7] )
         );
  DFF \stack_reg[0][8]  ( .D(n2574), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \stack_reg[1][8]  ( .D(n2573), .CLK(clk), .RST(rst), .Q(\stack[1][8] )
         );
  DFF \stack_reg[2][8]  ( .D(n2572), .CLK(clk), .RST(rst), .Q(\stack[2][8] )
         );
  DFF \stack_reg[3][8]  ( .D(n2571), .CLK(clk), .RST(rst), .Q(\stack[3][8] )
         );
  DFF \stack_reg[4][8]  ( .D(n2570), .CLK(clk), .RST(rst), .Q(\stack[4][8] )
         );
  DFF \stack_reg[5][8]  ( .D(n2569), .CLK(clk), .RST(rst), .Q(\stack[5][8] )
         );
  DFF \stack_reg[6][8]  ( .D(n2568), .CLK(clk), .RST(rst), .Q(\stack[6][8] )
         );
  DFF \stack_reg[7][8]  ( .D(n2567), .CLK(clk), .RST(rst), .Q(\stack[7][8] )
         );
  DFF \stack_reg[0][9]  ( .D(n2566), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \stack_reg[1][9]  ( .D(n2565), .CLK(clk), .RST(rst), .Q(\stack[1][9] )
         );
  DFF \stack_reg[2][9]  ( .D(n2564), .CLK(clk), .RST(rst), .Q(\stack[2][9] )
         );
  DFF \stack_reg[3][9]  ( .D(n2563), .CLK(clk), .RST(rst), .Q(\stack[3][9] )
         );
  DFF \stack_reg[4][9]  ( .D(n2562), .CLK(clk), .RST(rst), .Q(\stack[4][9] )
         );
  DFF \stack_reg[5][9]  ( .D(n2561), .CLK(clk), .RST(rst), .Q(\stack[5][9] )
         );
  DFF \stack_reg[6][9]  ( .D(n2560), .CLK(clk), .RST(rst), .Q(\stack[6][9] )
         );
  DFF \stack_reg[7][9]  ( .D(n2559), .CLK(clk), .RST(rst), .Q(\stack[7][9] )
         );
  DFF \stack_reg[0][10]  ( .D(n2558), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \stack_reg[1][10]  ( .D(n2557), .CLK(clk), .RST(rst), .Q(\stack[1][10] )
         );
  DFF \stack_reg[2][10]  ( .D(n2556), .CLK(clk), .RST(rst), .Q(\stack[2][10] )
         );
  DFF \stack_reg[3][10]  ( .D(n2555), .CLK(clk), .RST(rst), .Q(\stack[3][10] )
         );
  DFF \stack_reg[4][10]  ( .D(n2554), .CLK(clk), .RST(rst), .Q(\stack[4][10] )
         );
  DFF \stack_reg[5][10]  ( .D(n2553), .CLK(clk), .RST(rst), .Q(\stack[5][10] )
         );
  DFF \stack_reg[6][10]  ( .D(n2552), .CLK(clk), .RST(rst), .Q(\stack[6][10] )
         );
  DFF \stack_reg[7][10]  ( .D(n2551), .CLK(clk), .RST(rst), .Q(\stack[7][10] )
         );
  DFF \stack_reg[0][11]  ( .D(n2550), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \stack_reg[1][11]  ( .D(n2549), .CLK(clk), .RST(rst), .Q(\stack[1][11] )
         );
  DFF \stack_reg[2][11]  ( .D(n2548), .CLK(clk), .RST(rst), .Q(\stack[2][11] )
         );
  DFF \stack_reg[3][11]  ( .D(n2547), .CLK(clk), .RST(rst), .Q(\stack[3][11] )
         );
  DFF \stack_reg[4][11]  ( .D(n2546), .CLK(clk), .RST(rst), .Q(\stack[4][11] )
         );
  DFF \stack_reg[5][11]  ( .D(n2545), .CLK(clk), .RST(rst), .Q(\stack[5][11] )
         );
  DFF \stack_reg[6][11]  ( .D(n2544), .CLK(clk), .RST(rst), .Q(\stack[6][11] )
         );
  DFF \stack_reg[7][11]  ( .D(n2543), .CLK(clk), .RST(rst), .Q(\stack[7][11] )
         );
  DFF \stack_reg[0][12]  ( .D(n2542), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \stack_reg[1][12]  ( .D(n2541), .CLK(clk), .RST(rst), .Q(\stack[1][12] )
         );
  DFF \stack_reg[2][12]  ( .D(n2540), .CLK(clk), .RST(rst), .Q(\stack[2][12] )
         );
  DFF \stack_reg[3][12]  ( .D(n2539), .CLK(clk), .RST(rst), .Q(\stack[3][12] )
         );
  DFF \stack_reg[4][12]  ( .D(n2538), .CLK(clk), .RST(rst), .Q(\stack[4][12] )
         );
  DFF \stack_reg[5][12]  ( .D(n2537), .CLK(clk), .RST(rst), .Q(\stack[5][12] )
         );
  DFF \stack_reg[6][12]  ( .D(n2536), .CLK(clk), .RST(rst), .Q(\stack[6][12] )
         );
  DFF \stack_reg[7][12]  ( .D(n2535), .CLK(clk), .RST(rst), .Q(\stack[7][12] )
         );
  DFF \stack_reg[0][13]  ( .D(n2534), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \stack_reg[1][13]  ( .D(n2533), .CLK(clk), .RST(rst), .Q(\stack[1][13] )
         );
  DFF \stack_reg[2][13]  ( .D(n2532), .CLK(clk), .RST(rst), .Q(\stack[2][13] )
         );
  DFF \stack_reg[3][13]  ( .D(n2531), .CLK(clk), .RST(rst), .Q(\stack[3][13] )
         );
  DFF \stack_reg[4][13]  ( .D(n2530), .CLK(clk), .RST(rst), .Q(\stack[4][13] )
         );
  DFF \stack_reg[5][13]  ( .D(n2529), .CLK(clk), .RST(rst), .Q(\stack[5][13] )
         );
  DFF \stack_reg[6][13]  ( .D(n2528), .CLK(clk), .RST(rst), .Q(\stack[6][13] )
         );
  DFF \stack_reg[7][13]  ( .D(n2527), .CLK(clk), .RST(rst), .Q(\stack[7][13] )
         );
  DFF \stack_reg[0][14]  ( .D(n2526), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \stack_reg[1][14]  ( .D(n2525), .CLK(clk), .RST(rst), .Q(\stack[1][14] )
         );
  DFF \stack_reg[2][14]  ( .D(n2524), .CLK(clk), .RST(rst), .Q(\stack[2][14] )
         );
  DFF \stack_reg[3][14]  ( .D(n2523), .CLK(clk), .RST(rst), .Q(\stack[3][14] )
         );
  DFF \stack_reg[4][14]  ( .D(n2522), .CLK(clk), .RST(rst), .Q(\stack[4][14] )
         );
  DFF \stack_reg[5][14]  ( .D(n2521), .CLK(clk), .RST(rst), .Q(\stack[5][14] )
         );
  DFF \stack_reg[6][14]  ( .D(n2520), .CLK(clk), .RST(rst), .Q(\stack[6][14] )
         );
  DFF \stack_reg[7][14]  ( .D(n2519), .CLK(clk), .RST(rst), .Q(\stack[7][14] )
         );
  DFF \stack_reg[0][15]  ( .D(n2518), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \stack_reg[1][15]  ( .D(n2517), .CLK(clk), .RST(rst), .Q(\stack[1][15] )
         );
  DFF \stack_reg[2][15]  ( .D(n2516), .CLK(clk), .RST(rst), .Q(\stack[2][15] )
         );
  DFF \stack_reg[3][15]  ( .D(n2515), .CLK(clk), .RST(rst), .Q(\stack[3][15] )
         );
  DFF \stack_reg[4][15]  ( .D(n2514), .CLK(clk), .RST(rst), .Q(\stack[4][15] )
         );
  DFF \stack_reg[5][15]  ( .D(n2513), .CLK(clk), .RST(rst), .Q(\stack[5][15] )
         );
  DFF \stack_reg[6][15]  ( .D(n2512), .CLK(clk), .RST(rst), .Q(\stack[6][15] )
         );
  DFF \stack_reg[7][15]  ( .D(n2511), .CLK(clk), .RST(rst), .Q(\stack[7][15] )
         );
  DFF \stack_reg[0][16]  ( .D(n2510), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \stack_reg[1][16]  ( .D(n2509), .CLK(clk), .RST(rst), .Q(\stack[1][16] )
         );
  DFF \stack_reg[2][16]  ( .D(n2508), .CLK(clk), .RST(rst), .Q(\stack[2][16] )
         );
  DFF \stack_reg[3][16]  ( .D(n2507), .CLK(clk), .RST(rst), .Q(\stack[3][16] )
         );
  DFF \stack_reg[4][16]  ( .D(n2506), .CLK(clk), .RST(rst), .Q(\stack[4][16] )
         );
  DFF \stack_reg[5][16]  ( .D(n2505), .CLK(clk), .RST(rst), .Q(\stack[5][16] )
         );
  DFF \stack_reg[6][16]  ( .D(n2504), .CLK(clk), .RST(rst), .Q(\stack[6][16] )
         );
  DFF \stack_reg[7][16]  ( .D(n2503), .CLK(clk), .RST(rst), .Q(\stack[7][16] )
         );
  DFF \stack_reg[0][17]  ( .D(n2502), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \stack_reg[1][17]  ( .D(n2501), .CLK(clk), .RST(rst), .Q(\stack[1][17] )
         );
  DFF \stack_reg[2][17]  ( .D(n2500), .CLK(clk), .RST(rst), .Q(\stack[2][17] )
         );
  DFF \stack_reg[3][17]  ( .D(n2499), .CLK(clk), .RST(rst), .Q(\stack[3][17] )
         );
  DFF \stack_reg[4][17]  ( .D(n2498), .CLK(clk), .RST(rst), .Q(\stack[4][17] )
         );
  DFF \stack_reg[5][17]  ( .D(n2497), .CLK(clk), .RST(rst), .Q(\stack[5][17] )
         );
  DFF \stack_reg[6][17]  ( .D(n2496), .CLK(clk), .RST(rst), .Q(\stack[6][17] )
         );
  DFF \stack_reg[7][17]  ( .D(n2495), .CLK(clk), .RST(rst), .Q(\stack[7][17] )
         );
  DFF \stack_reg[0][18]  ( .D(n2494), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \stack_reg[1][18]  ( .D(n2493), .CLK(clk), .RST(rst), .Q(\stack[1][18] )
         );
  DFF \stack_reg[2][18]  ( .D(n2492), .CLK(clk), .RST(rst), .Q(\stack[2][18] )
         );
  DFF \stack_reg[3][18]  ( .D(n2491), .CLK(clk), .RST(rst), .Q(\stack[3][18] )
         );
  DFF \stack_reg[4][18]  ( .D(n2490), .CLK(clk), .RST(rst), .Q(\stack[4][18] )
         );
  DFF \stack_reg[5][18]  ( .D(n2489), .CLK(clk), .RST(rst), .Q(\stack[5][18] )
         );
  DFF \stack_reg[6][18]  ( .D(n2488), .CLK(clk), .RST(rst), .Q(\stack[6][18] )
         );
  DFF \stack_reg[7][18]  ( .D(n2487), .CLK(clk), .RST(rst), .Q(\stack[7][18] )
         );
  DFF \stack_reg[0][19]  ( .D(n2486), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \stack_reg[1][19]  ( .D(n2485), .CLK(clk), .RST(rst), .Q(\stack[1][19] )
         );
  DFF \stack_reg[2][19]  ( .D(n2484), .CLK(clk), .RST(rst), .Q(\stack[2][19] )
         );
  DFF \stack_reg[3][19]  ( .D(n2483), .CLK(clk), .RST(rst), .Q(\stack[3][19] )
         );
  DFF \stack_reg[4][19]  ( .D(n2482), .CLK(clk), .RST(rst), .Q(\stack[4][19] )
         );
  DFF \stack_reg[5][19]  ( .D(n2481), .CLK(clk), .RST(rst), .Q(\stack[5][19] )
         );
  DFF \stack_reg[6][19]  ( .D(n2480), .CLK(clk), .RST(rst), .Q(\stack[6][19] )
         );
  DFF \stack_reg[7][19]  ( .D(n2479), .CLK(clk), .RST(rst), .Q(\stack[7][19] )
         );
  DFF \stack_reg[0][20]  ( .D(n2478), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \stack_reg[1][20]  ( .D(n2477), .CLK(clk), .RST(rst), .Q(\stack[1][20] )
         );
  DFF \stack_reg[2][20]  ( .D(n2476), .CLK(clk), .RST(rst), .Q(\stack[2][20] )
         );
  DFF \stack_reg[3][20]  ( .D(n2475), .CLK(clk), .RST(rst), .Q(\stack[3][20] )
         );
  DFF \stack_reg[4][20]  ( .D(n2474), .CLK(clk), .RST(rst), .Q(\stack[4][20] )
         );
  DFF \stack_reg[5][20]  ( .D(n2473), .CLK(clk), .RST(rst), .Q(\stack[5][20] )
         );
  DFF \stack_reg[6][20]  ( .D(n2472), .CLK(clk), .RST(rst), .Q(\stack[6][20] )
         );
  DFF \stack_reg[7][20]  ( .D(n2471), .CLK(clk), .RST(rst), .Q(\stack[7][20] )
         );
  DFF \stack_reg[0][21]  ( .D(n2470), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \stack_reg[1][21]  ( .D(n2469), .CLK(clk), .RST(rst), .Q(\stack[1][21] )
         );
  DFF \stack_reg[2][21]  ( .D(n2468), .CLK(clk), .RST(rst), .Q(\stack[2][21] )
         );
  DFF \stack_reg[3][21]  ( .D(n2467), .CLK(clk), .RST(rst), .Q(\stack[3][21] )
         );
  DFF \stack_reg[4][21]  ( .D(n2466), .CLK(clk), .RST(rst), .Q(\stack[4][21] )
         );
  DFF \stack_reg[5][21]  ( .D(n2465), .CLK(clk), .RST(rst), .Q(\stack[5][21] )
         );
  DFF \stack_reg[6][21]  ( .D(n2464), .CLK(clk), .RST(rst), .Q(\stack[6][21] )
         );
  DFF \stack_reg[7][21]  ( .D(n2463), .CLK(clk), .RST(rst), .Q(\stack[7][21] )
         );
  DFF \stack_reg[0][22]  ( .D(n2462), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \stack_reg[1][22]  ( .D(n2461), .CLK(clk), .RST(rst), .Q(\stack[1][22] )
         );
  DFF \stack_reg[2][22]  ( .D(n2460), .CLK(clk), .RST(rst), .Q(\stack[2][22] )
         );
  DFF \stack_reg[3][22]  ( .D(n2459), .CLK(clk), .RST(rst), .Q(\stack[3][22] )
         );
  DFF \stack_reg[4][22]  ( .D(n2458), .CLK(clk), .RST(rst), .Q(\stack[4][22] )
         );
  DFF \stack_reg[5][22]  ( .D(n2457), .CLK(clk), .RST(rst), .Q(\stack[5][22] )
         );
  DFF \stack_reg[6][22]  ( .D(n2456), .CLK(clk), .RST(rst), .Q(\stack[6][22] )
         );
  DFF \stack_reg[7][22]  ( .D(n2455), .CLK(clk), .RST(rst), .Q(\stack[7][22] )
         );
  DFF \stack_reg[0][23]  ( .D(n2454), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \stack_reg[1][23]  ( .D(n2453), .CLK(clk), .RST(rst), .Q(\stack[1][23] )
         );
  DFF \stack_reg[2][23]  ( .D(n2452), .CLK(clk), .RST(rst), .Q(\stack[2][23] )
         );
  DFF \stack_reg[3][23]  ( .D(n2451), .CLK(clk), .RST(rst), .Q(\stack[3][23] )
         );
  DFF \stack_reg[4][23]  ( .D(n2450), .CLK(clk), .RST(rst), .Q(\stack[4][23] )
         );
  DFF \stack_reg[5][23]  ( .D(n2449), .CLK(clk), .RST(rst), .Q(\stack[5][23] )
         );
  DFF \stack_reg[6][23]  ( .D(n2448), .CLK(clk), .RST(rst), .Q(\stack[6][23] )
         );
  DFF \stack_reg[7][23]  ( .D(n2447), .CLK(clk), .RST(rst), .Q(\stack[7][23] )
         );
  DFF \stack_reg[0][24]  ( .D(n2446), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \stack_reg[1][24]  ( .D(n2445), .CLK(clk), .RST(rst), .Q(\stack[1][24] )
         );
  DFF \stack_reg[2][24]  ( .D(n2444), .CLK(clk), .RST(rst), .Q(\stack[2][24] )
         );
  DFF \stack_reg[3][24]  ( .D(n2443), .CLK(clk), .RST(rst), .Q(\stack[3][24] )
         );
  DFF \stack_reg[4][24]  ( .D(n2442), .CLK(clk), .RST(rst), .Q(\stack[4][24] )
         );
  DFF \stack_reg[5][24]  ( .D(n2441), .CLK(clk), .RST(rst), .Q(\stack[5][24] )
         );
  DFF \stack_reg[6][24]  ( .D(n2440), .CLK(clk), .RST(rst), .Q(\stack[6][24] )
         );
  DFF \stack_reg[7][24]  ( .D(n2439), .CLK(clk), .RST(rst), .Q(\stack[7][24] )
         );
  DFF \stack_reg[0][25]  ( .D(n2438), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \stack_reg[1][25]  ( .D(n2437), .CLK(clk), .RST(rst), .Q(\stack[1][25] )
         );
  DFF \stack_reg[2][25]  ( .D(n2436), .CLK(clk), .RST(rst), .Q(\stack[2][25] )
         );
  DFF \stack_reg[3][25]  ( .D(n2435), .CLK(clk), .RST(rst), .Q(\stack[3][25] )
         );
  DFF \stack_reg[4][25]  ( .D(n2434), .CLK(clk), .RST(rst), .Q(\stack[4][25] )
         );
  DFF \stack_reg[5][25]  ( .D(n2433), .CLK(clk), .RST(rst), .Q(\stack[5][25] )
         );
  DFF \stack_reg[6][25]  ( .D(n2432), .CLK(clk), .RST(rst), .Q(\stack[6][25] )
         );
  DFF \stack_reg[7][25]  ( .D(n2431), .CLK(clk), .RST(rst), .Q(\stack[7][25] )
         );
  DFF \stack_reg[0][26]  ( .D(n2430), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \stack_reg[1][26]  ( .D(n2429), .CLK(clk), .RST(rst), .Q(\stack[1][26] )
         );
  DFF \stack_reg[2][26]  ( .D(n2428), .CLK(clk), .RST(rst), .Q(\stack[2][26] )
         );
  DFF \stack_reg[3][26]  ( .D(n2427), .CLK(clk), .RST(rst), .Q(\stack[3][26] )
         );
  DFF \stack_reg[4][26]  ( .D(n2426), .CLK(clk), .RST(rst), .Q(\stack[4][26] )
         );
  DFF \stack_reg[5][26]  ( .D(n2425), .CLK(clk), .RST(rst), .Q(\stack[5][26] )
         );
  DFF \stack_reg[6][26]  ( .D(n2424), .CLK(clk), .RST(rst), .Q(\stack[6][26] )
         );
  DFF \stack_reg[7][26]  ( .D(n2423), .CLK(clk), .RST(rst), .Q(\stack[7][26] )
         );
  DFF \stack_reg[0][27]  ( .D(n2422), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \stack_reg[1][27]  ( .D(n2421), .CLK(clk), .RST(rst), .Q(\stack[1][27] )
         );
  DFF \stack_reg[2][27]  ( .D(n2420), .CLK(clk), .RST(rst), .Q(\stack[2][27] )
         );
  DFF \stack_reg[3][27]  ( .D(n2419), .CLK(clk), .RST(rst), .Q(\stack[3][27] )
         );
  DFF \stack_reg[4][27]  ( .D(n2418), .CLK(clk), .RST(rst), .Q(\stack[4][27] )
         );
  DFF \stack_reg[5][27]  ( .D(n2417), .CLK(clk), .RST(rst), .Q(\stack[5][27] )
         );
  DFF \stack_reg[6][27]  ( .D(n2416), .CLK(clk), .RST(rst), .Q(\stack[6][27] )
         );
  DFF \stack_reg[7][27]  ( .D(n2415), .CLK(clk), .RST(rst), .Q(\stack[7][27] )
         );
  DFF \stack_reg[0][28]  ( .D(n2414), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \stack_reg[1][28]  ( .D(n2413), .CLK(clk), .RST(rst), .Q(\stack[1][28] )
         );
  DFF \stack_reg[2][28]  ( .D(n2412), .CLK(clk), .RST(rst), .Q(\stack[2][28] )
         );
  DFF \stack_reg[3][28]  ( .D(n2411), .CLK(clk), .RST(rst), .Q(\stack[3][28] )
         );
  DFF \stack_reg[4][28]  ( .D(n2410), .CLK(clk), .RST(rst), .Q(\stack[4][28] )
         );
  DFF \stack_reg[5][28]  ( .D(n2409), .CLK(clk), .RST(rst), .Q(\stack[5][28] )
         );
  DFF \stack_reg[6][28]  ( .D(n2408), .CLK(clk), .RST(rst), .Q(\stack[6][28] )
         );
  DFF \stack_reg[7][28]  ( .D(n2407), .CLK(clk), .RST(rst), .Q(\stack[7][28] )
         );
  DFF \stack_reg[0][29]  ( .D(n2406), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \stack_reg[1][29]  ( .D(n2405), .CLK(clk), .RST(rst), .Q(\stack[1][29] )
         );
  DFF \stack_reg[2][29]  ( .D(n2404), .CLK(clk), .RST(rst), .Q(\stack[2][29] )
         );
  DFF \stack_reg[3][29]  ( .D(n2403), .CLK(clk), .RST(rst), .Q(\stack[3][29] )
         );
  DFF \stack_reg[4][29]  ( .D(n2402), .CLK(clk), .RST(rst), .Q(\stack[4][29] )
         );
  DFF \stack_reg[5][29]  ( .D(n2401), .CLK(clk), .RST(rst), .Q(\stack[5][29] )
         );
  DFF \stack_reg[6][29]  ( .D(n2400), .CLK(clk), .RST(rst), .Q(\stack[6][29] )
         );
  DFF \stack_reg[7][29]  ( .D(n2399), .CLK(clk), .RST(rst), .Q(\stack[7][29] )
         );
  DFF \stack_reg[0][30]  ( .D(n2398), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \stack_reg[1][30]  ( .D(n2397), .CLK(clk), .RST(rst), .Q(\stack[1][30] )
         );
  DFF \stack_reg[2][30]  ( .D(n2396), .CLK(clk), .RST(rst), .Q(\stack[2][30] )
         );
  DFF \stack_reg[3][30]  ( .D(n2395), .CLK(clk), .RST(rst), .Q(\stack[3][30] )
         );
  DFF \stack_reg[4][30]  ( .D(n2394), .CLK(clk), .RST(rst), .Q(\stack[4][30] )
         );
  DFF \stack_reg[5][30]  ( .D(n2393), .CLK(clk), .RST(rst), .Q(\stack[5][30] )
         );
  DFF \stack_reg[6][30]  ( .D(n2392), .CLK(clk), .RST(rst), .Q(\stack[6][30] )
         );
  DFF \stack_reg[7][30]  ( .D(n2391), .CLK(clk), .RST(rst), .Q(\stack[7][30] )
         );
  DFF \stack_reg[0][31]  ( .D(n2390), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \stack_reg[1][31]  ( .D(n2389), .CLK(clk), .RST(rst), .Q(\stack[1][31] )
         );
  DFF \stack_reg[2][31]  ( .D(n2388), .CLK(clk), .RST(rst), .Q(\stack[2][31] )
         );
  DFF \stack_reg[3][31]  ( .D(n2387), .CLK(clk), .RST(rst), .Q(\stack[3][31] )
         );
  DFF \stack_reg[4][31]  ( .D(n2386), .CLK(clk), .RST(rst), .Q(\stack[4][31] )
         );
  DFF \stack_reg[5][31]  ( .D(n2385), .CLK(clk), .RST(rst), .Q(\stack[5][31] )
         );
  DFF \stack_reg[6][31]  ( .D(n2384), .CLK(clk), .RST(rst), .Q(\stack[6][31] )
         );
  DFF \stack_reg[7][31]  ( .D(n2383), .CLK(clk), .RST(rst), .Q(\stack[7][31] )
         );
  DFF \stack_reg[0][32]  ( .D(n2382), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \stack_reg[1][32]  ( .D(n2381), .CLK(clk), .RST(rst), .Q(\stack[1][32] )
         );
  DFF \stack_reg[2][32]  ( .D(n2380), .CLK(clk), .RST(rst), .Q(\stack[2][32] )
         );
  DFF \stack_reg[3][32]  ( .D(n2379), .CLK(clk), .RST(rst), .Q(\stack[3][32] )
         );
  DFF \stack_reg[4][32]  ( .D(n2378), .CLK(clk), .RST(rst), .Q(\stack[4][32] )
         );
  DFF \stack_reg[5][32]  ( .D(n2377), .CLK(clk), .RST(rst), .Q(\stack[5][32] )
         );
  DFF \stack_reg[6][32]  ( .D(n2376), .CLK(clk), .RST(rst), .Q(\stack[6][32] )
         );
  DFF \stack_reg[7][32]  ( .D(n2375), .CLK(clk), .RST(rst), .Q(\stack[7][32] )
         );
  DFF \stack_reg[0][33]  ( .D(n2374), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \stack_reg[1][33]  ( .D(n2373), .CLK(clk), .RST(rst), .Q(\stack[1][33] )
         );
  DFF \stack_reg[2][33]  ( .D(n2372), .CLK(clk), .RST(rst), .Q(\stack[2][33] )
         );
  DFF \stack_reg[3][33]  ( .D(n2371), .CLK(clk), .RST(rst), .Q(\stack[3][33] )
         );
  DFF \stack_reg[4][33]  ( .D(n2370), .CLK(clk), .RST(rst), .Q(\stack[4][33] )
         );
  DFF \stack_reg[5][33]  ( .D(n2369), .CLK(clk), .RST(rst), .Q(\stack[5][33] )
         );
  DFF \stack_reg[6][33]  ( .D(n2368), .CLK(clk), .RST(rst), .Q(\stack[6][33] )
         );
  DFF \stack_reg[7][33]  ( .D(n2367), .CLK(clk), .RST(rst), .Q(\stack[7][33] )
         );
  DFF \stack_reg[0][34]  ( .D(n2366), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \stack_reg[1][34]  ( .D(n2365), .CLK(clk), .RST(rst), .Q(\stack[1][34] )
         );
  DFF \stack_reg[2][34]  ( .D(n2364), .CLK(clk), .RST(rst), .Q(\stack[2][34] )
         );
  DFF \stack_reg[3][34]  ( .D(n2363), .CLK(clk), .RST(rst), .Q(\stack[3][34] )
         );
  DFF \stack_reg[4][34]  ( .D(n2362), .CLK(clk), .RST(rst), .Q(\stack[4][34] )
         );
  DFF \stack_reg[5][34]  ( .D(n2361), .CLK(clk), .RST(rst), .Q(\stack[5][34] )
         );
  DFF \stack_reg[6][34]  ( .D(n2360), .CLK(clk), .RST(rst), .Q(\stack[6][34] )
         );
  DFF \stack_reg[7][34]  ( .D(n2359), .CLK(clk), .RST(rst), .Q(\stack[7][34] )
         );
  DFF \stack_reg[0][35]  ( .D(n2358), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \stack_reg[1][35]  ( .D(n2357), .CLK(clk), .RST(rst), .Q(\stack[1][35] )
         );
  DFF \stack_reg[2][35]  ( .D(n2356), .CLK(clk), .RST(rst), .Q(\stack[2][35] )
         );
  DFF \stack_reg[3][35]  ( .D(n2355), .CLK(clk), .RST(rst), .Q(\stack[3][35] )
         );
  DFF \stack_reg[4][35]  ( .D(n2354), .CLK(clk), .RST(rst), .Q(\stack[4][35] )
         );
  DFF \stack_reg[5][35]  ( .D(n2353), .CLK(clk), .RST(rst), .Q(\stack[5][35] )
         );
  DFF \stack_reg[6][35]  ( .D(n2352), .CLK(clk), .RST(rst), .Q(\stack[6][35] )
         );
  DFF \stack_reg[7][35]  ( .D(n2351), .CLK(clk), .RST(rst), .Q(\stack[7][35] )
         );
  DFF \stack_reg[0][36]  ( .D(n2350), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \stack_reg[1][36]  ( .D(n2349), .CLK(clk), .RST(rst), .Q(\stack[1][36] )
         );
  DFF \stack_reg[2][36]  ( .D(n2348), .CLK(clk), .RST(rst), .Q(\stack[2][36] )
         );
  DFF \stack_reg[3][36]  ( .D(n2347), .CLK(clk), .RST(rst), .Q(\stack[3][36] )
         );
  DFF \stack_reg[4][36]  ( .D(n2346), .CLK(clk), .RST(rst), .Q(\stack[4][36] )
         );
  DFF \stack_reg[5][36]  ( .D(n2345), .CLK(clk), .RST(rst), .Q(\stack[5][36] )
         );
  DFF \stack_reg[6][36]  ( .D(n2344), .CLK(clk), .RST(rst), .Q(\stack[6][36] )
         );
  DFF \stack_reg[7][36]  ( .D(n2343), .CLK(clk), .RST(rst), .Q(\stack[7][36] )
         );
  DFF \stack_reg[0][37]  ( .D(n2342), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \stack_reg[1][37]  ( .D(n2341), .CLK(clk), .RST(rst), .Q(\stack[1][37] )
         );
  DFF \stack_reg[2][37]  ( .D(n2340), .CLK(clk), .RST(rst), .Q(\stack[2][37] )
         );
  DFF \stack_reg[3][37]  ( .D(n2339), .CLK(clk), .RST(rst), .Q(\stack[3][37] )
         );
  DFF \stack_reg[4][37]  ( .D(n2338), .CLK(clk), .RST(rst), .Q(\stack[4][37] )
         );
  DFF \stack_reg[5][37]  ( .D(n2337), .CLK(clk), .RST(rst), .Q(\stack[5][37] )
         );
  DFF \stack_reg[6][37]  ( .D(n2336), .CLK(clk), .RST(rst), .Q(\stack[6][37] )
         );
  DFF \stack_reg[7][37]  ( .D(n2335), .CLK(clk), .RST(rst), .Q(\stack[7][37] )
         );
  DFF \stack_reg[0][38]  ( .D(n2334), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \stack_reg[1][38]  ( .D(n2333), .CLK(clk), .RST(rst), .Q(\stack[1][38] )
         );
  DFF \stack_reg[2][38]  ( .D(n2332), .CLK(clk), .RST(rst), .Q(\stack[2][38] )
         );
  DFF \stack_reg[3][38]  ( .D(n2331), .CLK(clk), .RST(rst), .Q(\stack[3][38] )
         );
  DFF \stack_reg[4][38]  ( .D(n2330), .CLK(clk), .RST(rst), .Q(\stack[4][38] )
         );
  DFF \stack_reg[5][38]  ( .D(n2329), .CLK(clk), .RST(rst), .Q(\stack[5][38] )
         );
  DFF \stack_reg[6][38]  ( .D(n2328), .CLK(clk), .RST(rst), .Q(\stack[6][38] )
         );
  DFF \stack_reg[7][38]  ( .D(n2327), .CLK(clk), .RST(rst), .Q(\stack[7][38] )
         );
  DFF \stack_reg[0][39]  ( .D(n2326), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \stack_reg[1][39]  ( .D(n2325), .CLK(clk), .RST(rst), .Q(\stack[1][39] )
         );
  DFF \stack_reg[2][39]  ( .D(n2324), .CLK(clk), .RST(rst), .Q(\stack[2][39] )
         );
  DFF \stack_reg[3][39]  ( .D(n2323), .CLK(clk), .RST(rst), .Q(\stack[3][39] )
         );
  DFF \stack_reg[4][39]  ( .D(n2322), .CLK(clk), .RST(rst), .Q(\stack[4][39] )
         );
  DFF \stack_reg[5][39]  ( .D(n2321), .CLK(clk), .RST(rst), .Q(\stack[5][39] )
         );
  DFF \stack_reg[6][39]  ( .D(n2320), .CLK(clk), .RST(rst), .Q(\stack[6][39] )
         );
  DFF \stack_reg[7][39]  ( .D(n2319), .CLK(clk), .RST(rst), .Q(\stack[7][39] )
         );
  DFF \stack_reg[0][40]  ( .D(n2318), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \stack_reg[1][40]  ( .D(n2317), .CLK(clk), .RST(rst), .Q(\stack[1][40] )
         );
  DFF \stack_reg[2][40]  ( .D(n2316), .CLK(clk), .RST(rst), .Q(\stack[2][40] )
         );
  DFF \stack_reg[3][40]  ( .D(n2315), .CLK(clk), .RST(rst), .Q(\stack[3][40] )
         );
  DFF \stack_reg[4][40]  ( .D(n2314), .CLK(clk), .RST(rst), .Q(\stack[4][40] )
         );
  DFF \stack_reg[5][40]  ( .D(n2313), .CLK(clk), .RST(rst), .Q(\stack[5][40] )
         );
  DFF \stack_reg[6][40]  ( .D(n2312), .CLK(clk), .RST(rst), .Q(\stack[6][40] )
         );
  DFF \stack_reg[7][40]  ( .D(n2311), .CLK(clk), .RST(rst), .Q(\stack[7][40] )
         );
  DFF \stack_reg[0][41]  ( .D(n2310), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \stack_reg[1][41]  ( .D(n2309), .CLK(clk), .RST(rst), .Q(\stack[1][41] )
         );
  DFF \stack_reg[2][41]  ( .D(n2308), .CLK(clk), .RST(rst), .Q(\stack[2][41] )
         );
  DFF \stack_reg[3][41]  ( .D(n2307), .CLK(clk), .RST(rst), .Q(\stack[3][41] )
         );
  DFF \stack_reg[4][41]  ( .D(n2306), .CLK(clk), .RST(rst), .Q(\stack[4][41] )
         );
  DFF \stack_reg[5][41]  ( .D(n2305), .CLK(clk), .RST(rst), .Q(\stack[5][41] )
         );
  DFF \stack_reg[6][41]  ( .D(n2304), .CLK(clk), .RST(rst), .Q(\stack[6][41] )
         );
  DFF \stack_reg[7][41]  ( .D(n2303), .CLK(clk), .RST(rst), .Q(\stack[7][41] )
         );
  DFF \stack_reg[0][42]  ( .D(n2302), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \stack_reg[1][42]  ( .D(n2301), .CLK(clk), .RST(rst), .Q(\stack[1][42] )
         );
  DFF \stack_reg[2][42]  ( .D(n2300), .CLK(clk), .RST(rst), .Q(\stack[2][42] )
         );
  DFF \stack_reg[3][42]  ( .D(n2299), .CLK(clk), .RST(rst), .Q(\stack[3][42] )
         );
  DFF \stack_reg[4][42]  ( .D(n2298), .CLK(clk), .RST(rst), .Q(\stack[4][42] )
         );
  DFF \stack_reg[5][42]  ( .D(n2297), .CLK(clk), .RST(rst), .Q(\stack[5][42] )
         );
  DFF \stack_reg[6][42]  ( .D(n2296), .CLK(clk), .RST(rst), .Q(\stack[6][42] )
         );
  DFF \stack_reg[7][42]  ( .D(n2295), .CLK(clk), .RST(rst), .Q(\stack[7][42] )
         );
  DFF \stack_reg[0][43]  ( .D(n2294), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \stack_reg[1][43]  ( .D(n2293), .CLK(clk), .RST(rst), .Q(\stack[1][43] )
         );
  DFF \stack_reg[2][43]  ( .D(n2292), .CLK(clk), .RST(rst), .Q(\stack[2][43] )
         );
  DFF \stack_reg[3][43]  ( .D(n2291), .CLK(clk), .RST(rst), .Q(\stack[3][43] )
         );
  DFF \stack_reg[4][43]  ( .D(n2290), .CLK(clk), .RST(rst), .Q(\stack[4][43] )
         );
  DFF \stack_reg[5][43]  ( .D(n2289), .CLK(clk), .RST(rst), .Q(\stack[5][43] )
         );
  DFF \stack_reg[6][43]  ( .D(n2288), .CLK(clk), .RST(rst), .Q(\stack[6][43] )
         );
  DFF \stack_reg[7][43]  ( .D(n2287), .CLK(clk), .RST(rst), .Q(\stack[7][43] )
         );
  DFF \stack_reg[0][44]  ( .D(n2286), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \stack_reg[1][44]  ( .D(n2285), .CLK(clk), .RST(rst), .Q(\stack[1][44] )
         );
  DFF \stack_reg[2][44]  ( .D(n2284), .CLK(clk), .RST(rst), .Q(\stack[2][44] )
         );
  DFF \stack_reg[3][44]  ( .D(n2283), .CLK(clk), .RST(rst), .Q(\stack[3][44] )
         );
  DFF \stack_reg[4][44]  ( .D(n2282), .CLK(clk), .RST(rst), .Q(\stack[4][44] )
         );
  DFF \stack_reg[5][44]  ( .D(n2281), .CLK(clk), .RST(rst), .Q(\stack[5][44] )
         );
  DFF \stack_reg[6][44]  ( .D(n2280), .CLK(clk), .RST(rst), .Q(\stack[6][44] )
         );
  DFF \stack_reg[7][44]  ( .D(n2279), .CLK(clk), .RST(rst), .Q(\stack[7][44] )
         );
  DFF \stack_reg[0][45]  ( .D(n2278), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \stack_reg[1][45]  ( .D(n2277), .CLK(clk), .RST(rst), .Q(\stack[1][45] )
         );
  DFF \stack_reg[2][45]  ( .D(n2276), .CLK(clk), .RST(rst), .Q(\stack[2][45] )
         );
  DFF \stack_reg[3][45]  ( .D(n2275), .CLK(clk), .RST(rst), .Q(\stack[3][45] )
         );
  DFF \stack_reg[4][45]  ( .D(n2274), .CLK(clk), .RST(rst), .Q(\stack[4][45] )
         );
  DFF \stack_reg[5][45]  ( .D(n2273), .CLK(clk), .RST(rst), .Q(\stack[5][45] )
         );
  DFF \stack_reg[6][45]  ( .D(n2272), .CLK(clk), .RST(rst), .Q(\stack[6][45] )
         );
  DFF \stack_reg[7][45]  ( .D(n2271), .CLK(clk), .RST(rst), .Q(\stack[7][45] )
         );
  DFF \stack_reg[0][46]  ( .D(n2270), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \stack_reg[1][46]  ( .D(n2269), .CLK(clk), .RST(rst), .Q(\stack[1][46] )
         );
  DFF \stack_reg[2][46]  ( .D(n2268), .CLK(clk), .RST(rst), .Q(\stack[2][46] )
         );
  DFF \stack_reg[3][46]  ( .D(n2267), .CLK(clk), .RST(rst), .Q(\stack[3][46] )
         );
  DFF \stack_reg[4][46]  ( .D(n2266), .CLK(clk), .RST(rst), .Q(\stack[4][46] )
         );
  DFF \stack_reg[5][46]  ( .D(n2265), .CLK(clk), .RST(rst), .Q(\stack[5][46] )
         );
  DFF \stack_reg[6][46]  ( .D(n2264), .CLK(clk), .RST(rst), .Q(\stack[6][46] )
         );
  DFF \stack_reg[7][46]  ( .D(n2263), .CLK(clk), .RST(rst), .Q(\stack[7][46] )
         );
  DFF \stack_reg[0][47]  ( .D(n2262), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \stack_reg[1][47]  ( .D(n2261), .CLK(clk), .RST(rst), .Q(\stack[1][47] )
         );
  DFF \stack_reg[2][47]  ( .D(n2260), .CLK(clk), .RST(rst), .Q(\stack[2][47] )
         );
  DFF \stack_reg[3][47]  ( .D(n2259), .CLK(clk), .RST(rst), .Q(\stack[3][47] )
         );
  DFF \stack_reg[4][47]  ( .D(n2258), .CLK(clk), .RST(rst), .Q(\stack[4][47] )
         );
  DFF \stack_reg[5][47]  ( .D(n2257), .CLK(clk), .RST(rst), .Q(\stack[5][47] )
         );
  DFF \stack_reg[6][47]  ( .D(n2256), .CLK(clk), .RST(rst), .Q(\stack[6][47] )
         );
  DFF \stack_reg[7][47]  ( .D(n2255), .CLK(clk), .RST(rst), .Q(\stack[7][47] )
         );
  DFF \stack_reg[0][48]  ( .D(n2254), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \stack_reg[1][48]  ( .D(n2253), .CLK(clk), .RST(rst), .Q(\stack[1][48] )
         );
  DFF \stack_reg[2][48]  ( .D(n2252), .CLK(clk), .RST(rst), .Q(\stack[2][48] )
         );
  DFF \stack_reg[3][48]  ( .D(n2251), .CLK(clk), .RST(rst), .Q(\stack[3][48] )
         );
  DFF \stack_reg[4][48]  ( .D(n2250), .CLK(clk), .RST(rst), .Q(\stack[4][48] )
         );
  DFF \stack_reg[5][48]  ( .D(n2249), .CLK(clk), .RST(rst), .Q(\stack[5][48] )
         );
  DFF \stack_reg[6][48]  ( .D(n2248), .CLK(clk), .RST(rst), .Q(\stack[6][48] )
         );
  DFF \stack_reg[7][48]  ( .D(n2247), .CLK(clk), .RST(rst), .Q(\stack[7][48] )
         );
  DFF \stack_reg[0][49]  ( .D(n2246), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \stack_reg[1][49]  ( .D(n2245), .CLK(clk), .RST(rst), .Q(\stack[1][49] )
         );
  DFF \stack_reg[2][49]  ( .D(n2244), .CLK(clk), .RST(rst), .Q(\stack[2][49] )
         );
  DFF \stack_reg[3][49]  ( .D(n2243), .CLK(clk), .RST(rst), .Q(\stack[3][49] )
         );
  DFF \stack_reg[4][49]  ( .D(n2242), .CLK(clk), .RST(rst), .Q(\stack[4][49] )
         );
  DFF \stack_reg[5][49]  ( .D(n2241), .CLK(clk), .RST(rst), .Q(\stack[5][49] )
         );
  DFF \stack_reg[6][49]  ( .D(n2240), .CLK(clk), .RST(rst), .Q(\stack[6][49] )
         );
  DFF \stack_reg[7][49]  ( .D(n2239), .CLK(clk), .RST(rst), .Q(\stack[7][49] )
         );
  DFF \stack_reg[0][50]  ( .D(n2238), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \stack_reg[1][50]  ( .D(n2237), .CLK(clk), .RST(rst), .Q(\stack[1][50] )
         );
  DFF \stack_reg[2][50]  ( .D(n2236), .CLK(clk), .RST(rst), .Q(\stack[2][50] )
         );
  DFF \stack_reg[3][50]  ( .D(n2235), .CLK(clk), .RST(rst), .Q(\stack[3][50] )
         );
  DFF \stack_reg[4][50]  ( .D(n2234), .CLK(clk), .RST(rst), .Q(\stack[4][50] )
         );
  DFF \stack_reg[5][50]  ( .D(n2233), .CLK(clk), .RST(rst), .Q(\stack[5][50] )
         );
  DFF \stack_reg[6][50]  ( .D(n2232), .CLK(clk), .RST(rst), .Q(\stack[6][50] )
         );
  DFF \stack_reg[7][50]  ( .D(n2231), .CLK(clk), .RST(rst), .Q(\stack[7][50] )
         );
  DFF \stack_reg[0][51]  ( .D(n2230), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \stack_reg[1][51]  ( .D(n2229), .CLK(clk), .RST(rst), .Q(\stack[1][51] )
         );
  DFF \stack_reg[2][51]  ( .D(n2228), .CLK(clk), .RST(rst), .Q(\stack[2][51] )
         );
  DFF \stack_reg[3][51]  ( .D(n2227), .CLK(clk), .RST(rst), .Q(\stack[3][51] )
         );
  DFF \stack_reg[4][51]  ( .D(n2226), .CLK(clk), .RST(rst), .Q(\stack[4][51] )
         );
  DFF \stack_reg[5][51]  ( .D(n2225), .CLK(clk), .RST(rst), .Q(\stack[5][51] )
         );
  DFF \stack_reg[6][51]  ( .D(n2224), .CLK(clk), .RST(rst), .Q(\stack[6][51] )
         );
  DFF \stack_reg[7][51]  ( .D(n2223), .CLK(clk), .RST(rst), .Q(\stack[7][51] )
         );
  DFF \stack_reg[0][52]  ( .D(n2222), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \stack_reg[1][52]  ( .D(n2221), .CLK(clk), .RST(rst), .Q(\stack[1][52] )
         );
  DFF \stack_reg[2][52]  ( .D(n2220), .CLK(clk), .RST(rst), .Q(\stack[2][52] )
         );
  DFF \stack_reg[3][52]  ( .D(n2219), .CLK(clk), .RST(rst), .Q(\stack[3][52] )
         );
  DFF \stack_reg[4][52]  ( .D(n2218), .CLK(clk), .RST(rst), .Q(\stack[4][52] )
         );
  DFF \stack_reg[5][52]  ( .D(n2217), .CLK(clk), .RST(rst), .Q(\stack[5][52] )
         );
  DFF \stack_reg[6][52]  ( .D(n2216), .CLK(clk), .RST(rst), .Q(\stack[6][52] )
         );
  DFF \stack_reg[7][52]  ( .D(n2215), .CLK(clk), .RST(rst), .Q(\stack[7][52] )
         );
  DFF \stack_reg[0][53]  ( .D(n2214), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \stack_reg[1][53]  ( .D(n2213), .CLK(clk), .RST(rst), .Q(\stack[1][53] )
         );
  DFF \stack_reg[2][53]  ( .D(n2212), .CLK(clk), .RST(rst), .Q(\stack[2][53] )
         );
  DFF \stack_reg[3][53]  ( .D(n2211), .CLK(clk), .RST(rst), .Q(\stack[3][53] )
         );
  DFF \stack_reg[4][53]  ( .D(n2210), .CLK(clk), .RST(rst), .Q(\stack[4][53] )
         );
  DFF \stack_reg[5][53]  ( .D(n2209), .CLK(clk), .RST(rst), .Q(\stack[5][53] )
         );
  DFF \stack_reg[6][53]  ( .D(n2208), .CLK(clk), .RST(rst), .Q(\stack[6][53] )
         );
  DFF \stack_reg[7][53]  ( .D(n2207), .CLK(clk), .RST(rst), .Q(\stack[7][53] )
         );
  DFF \stack_reg[0][54]  ( .D(n2206), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \stack_reg[1][54]  ( .D(n2205), .CLK(clk), .RST(rst), .Q(\stack[1][54] )
         );
  DFF \stack_reg[2][54]  ( .D(n2204), .CLK(clk), .RST(rst), .Q(\stack[2][54] )
         );
  DFF \stack_reg[3][54]  ( .D(n2203), .CLK(clk), .RST(rst), .Q(\stack[3][54] )
         );
  DFF \stack_reg[4][54]  ( .D(n2202), .CLK(clk), .RST(rst), .Q(\stack[4][54] )
         );
  DFF \stack_reg[5][54]  ( .D(n2201), .CLK(clk), .RST(rst), .Q(\stack[5][54] )
         );
  DFF \stack_reg[6][54]  ( .D(n2200), .CLK(clk), .RST(rst), .Q(\stack[6][54] )
         );
  DFF \stack_reg[7][54]  ( .D(n2199), .CLK(clk), .RST(rst), .Q(\stack[7][54] )
         );
  DFF \stack_reg[0][55]  ( .D(n2198), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \stack_reg[1][55]  ( .D(n2197), .CLK(clk), .RST(rst), .Q(\stack[1][55] )
         );
  DFF \stack_reg[2][55]  ( .D(n2196), .CLK(clk), .RST(rst), .Q(\stack[2][55] )
         );
  DFF \stack_reg[3][55]  ( .D(n2195), .CLK(clk), .RST(rst), .Q(\stack[3][55] )
         );
  DFF \stack_reg[4][55]  ( .D(n2194), .CLK(clk), .RST(rst), .Q(\stack[4][55] )
         );
  DFF \stack_reg[5][55]  ( .D(n2193), .CLK(clk), .RST(rst), .Q(\stack[5][55] )
         );
  DFF \stack_reg[6][55]  ( .D(n2192), .CLK(clk), .RST(rst), .Q(\stack[6][55] )
         );
  DFF \stack_reg[7][55]  ( .D(n2191), .CLK(clk), .RST(rst), .Q(\stack[7][55] )
         );
  DFF \stack_reg[0][56]  ( .D(n2190), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \stack_reg[1][56]  ( .D(n2189), .CLK(clk), .RST(rst), .Q(\stack[1][56] )
         );
  DFF \stack_reg[2][56]  ( .D(n2188), .CLK(clk), .RST(rst), .Q(\stack[2][56] )
         );
  DFF \stack_reg[3][56]  ( .D(n2187), .CLK(clk), .RST(rst), .Q(\stack[3][56] )
         );
  DFF \stack_reg[4][56]  ( .D(n2186), .CLK(clk), .RST(rst), .Q(\stack[4][56] )
         );
  DFF \stack_reg[5][56]  ( .D(n2185), .CLK(clk), .RST(rst), .Q(\stack[5][56] )
         );
  DFF \stack_reg[6][56]  ( .D(n2184), .CLK(clk), .RST(rst), .Q(\stack[6][56] )
         );
  DFF \stack_reg[7][56]  ( .D(n2183), .CLK(clk), .RST(rst), .Q(\stack[7][56] )
         );
  DFF \stack_reg[0][57]  ( .D(n2182), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \stack_reg[1][57]  ( .D(n2181), .CLK(clk), .RST(rst), .Q(\stack[1][57] )
         );
  DFF \stack_reg[2][57]  ( .D(n2180), .CLK(clk), .RST(rst), .Q(\stack[2][57] )
         );
  DFF \stack_reg[3][57]  ( .D(n2179), .CLK(clk), .RST(rst), .Q(\stack[3][57] )
         );
  DFF \stack_reg[4][57]  ( .D(n2178), .CLK(clk), .RST(rst), .Q(\stack[4][57] )
         );
  DFF \stack_reg[5][57]  ( .D(n2177), .CLK(clk), .RST(rst), .Q(\stack[5][57] )
         );
  DFF \stack_reg[6][57]  ( .D(n2176), .CLK(clk), .RST(rst), .Q(\stack[6][57] )
         );
  DFF \stack_reg[7][57]  ( .D(n2175), .CLK(clk), .RST(rst), .Q(\stack[7][57] )
         );
  DFF \stack_reg[0][58]  ( .D(n2174), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \stack_reg[1][58]  ( .D(n2173), .CLK(clk), .RST(rst), .Q(\stack[1][58] )
         );
  DFF \stack_reg[2][58]  ( .D(n2172), .CLK(clk), .RST(rst), .Q(\stack[2][58] )
         );
  DFF \stack_reg[3][58]  ( .D(n2171), .CLK(clk), .RST(rst), .Q(\stack[3][58] )
         );
  DFF \stack_reg[4][58]  ( .D(n2170), .CLK(clk), .RST(rst), .Q(\stack[4][58] )
         );
  DFF \stack_reg[5][58]  ( .D(n2169), .CLK(clk), .RST(rst), .Q(\stack[5][58] )
         );
  DFF \stack_reg[6][58]  ( .D(n2168), .CLK(clk), .RST(rst), .Q(\stack[6][58] )
         );
  DFF \stack_reg[7][58]  ( .D(n2167), .CLK(clk), .RST(rst), .Q(\stack[7][58] )
         );
  DFF \stack_reg[0][59]  ( .D(n2166), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \stack_reg[1][59]  ( .D(n2165), .CLK(clk), .RST(rst), .Q(\stack[1][59] )
         );
  DFF \stack_reg[2][59]  ( .D(n2164), .CLK(clk), .RST(rst), .Q(\stack[2][59] )
         );
  DFF \stack_reg[3][59]  ( .D(n2163), .CLK(clk), .RST(rst), .Q(\stack[3][59] )
         );
  DFF \stack_reg[4][59]  ( .D(n2162), .CLK(clk), .RST(rst), .Q(\stack[4][59] )
         );
  DFF \stack_reg[5][59]  ( .D(n2161), .CLK(clk), .RST(rst), .Q(\stack[5][59] )
         );
  DFF \stack_reg[6][59]  ( .D(n2160), .CLK(clk), .RST(rst), .Q(\stack[6][59] )
         );
  DFF \stack_reg[7][59]  ( .D(n2159), .CLK(clk), .RST(rst), .Q(\stack[7][59] )
         );
  DFF \stack_reg[0][60]  ( .D(n2158), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \stack_reg[1][60]  ( .D(n2157), .CLK(clk), .RST(rst), .Q(\stack[1][60] )
         );
  DFF \stack_reg[2][60]  ( .D(n2156), .CLK(clk), .RST(rst), .Q(\stack[2][60] )
         );
  DFF \stack_reg[3][60]  ( .D(n2155), .CLK(clk), .RST(rst), .Q(\stack[3][60] )
         );
  DFF \stack_reg[4][60]  ( .D(n2154), .CLK(clk), .RST(rst), .Q(\stack[4][60] )
         );
  DFF \stack_reg[5][60]  ( .D(n2153), .CLK(clk), .RST(rst), .Q(\stack[5][60] )
         );
  DFF \stack_reg[6][60]  ( .D(n2152), .CLK(clk), .RST(rst), .Q(\stack[6][60] )
         );
  DFF \stack_reg[7][60]  ( .D(n2151), .CLK(clk), .RST(rst), .Q(\stack[7][60] )
         );
  DFF \stack_reg[0][61]  ( .D(n2150), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \stack_reg[1][61]  ( .D(n2149), .CLK(clk), .RST(rst), .Q(\stack[1][61] )
         );
  DFF \stack_reg[2][61]  ( .D(n2148), .CLK(clk), .RST(rst), .Q(\stack[2][61] )
         );
  DFF \stack_reg[3][61]  ( .D(n2147), .CLK(clk), .RST(rst), .Q(\stack[3][61] )
         );
  DFF \stack_reg[4][61]  ( .D(n2146), .CLK(clk), .RST(rst), .Q(\stack[4][61] )
         );
  DFF \stack_reg[5][61]  ( .D(n2145), .CLK(clk), .RST(rst), .Q(\stack[5][61] )
         );
  DFF \stack_reg[6][61]  ( .D(n2144), .CLK(clk), .RST(rst), .Q(\stack[6][61] )
         );
  DFF \stack_reg[7][61]  ( .D(n2143), .CLK(clk), .RST(rst), .Q(\stack[7][61] )
         );
  DFF \stack_reg[0][62]  ( .D(n2142), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \stack_reg[1][62]  ( .D(n2141), .CLK(clk), .RST(rst), .Q(\stack[1][62] )
         );
  DFF \stack_reg[2][62]  ( .D(n2140), .CLK(clk), .RST(rst), .Q(\stack[2][62] )
         );
  DFF \stack_reg[3][62]  ( .D(n2139), .CLK(clk), .RST(rst), .Q(\stack[3][62] )
         );
  DFF \stack_reg[4][62]  ( .D(n2138), .CLK(clk), .RST(rst), .Q(\stack[4][62] )
         );
  DFF \stack_reg[5][62]  ( .D(n2137), .CLK(clk), .RST(rst), .Q(\stack[5][62] )
         );
  DFF \stack_reg[6][62]  ( .D(n2136), .CLK(clk), .RST(rst), .Q(\stack[6][62] )
         );
  DFF \stack_reg[7][62]  ( .D(n2135), .CLK(clk), .RST(rst), .Q(\stack[7][62] )
         );
  DFF \stack_reg[0][63]  ( .D(n2134), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \stack_reg[1][63]  ( .D(n2133), .CLK(clk), .RST(rst), .Q(\stack[1][63] )
         );
  DFF \stack_reg[2][63]  ( .D(n2132), .CLK(clk), .RST(rst), .Q(\stack[2][63] )
         );
  DFF \stack_reg[3][63]  ( .D(n2131), .CLK(clk), .RST(rst), .Q(\stack[3][63] )
         );
  DFF \stack_reg[4][63]  ( .D(n2130), .CLK(clk), .RST(rst), .Q(\stack[4][63] )
         );
  DFF \stack_reg[5][63]  ( .D(n2129), .CLK(clk), .RST(rst), .Q(\stack[5][63] )
         );
  DFF \stack_reg[6][63]  ( .D(n2128), .CLK(clk), .RST(rst), .Q(\stack[6][63] )
         );
  DFF \stack_reg[7][63]  ( .D(n2127), .CLK(clk), .RST(rst), .Q(\stack[7][63] )
         );
  DFF \stack_reg[2][0]  ( .D(n2126), .CLK(clk), .RST(rst), .Q(\stack[2][0] )
         );
  DFF \stack_reg[3][0]  ( .D(n2125), .CLK(clk), .RST(rst), .Q(\stack[3][0] )
         );
  DFF \stack_reg[4][0]  ( .D(n2124), .CLK(clk), .RST(rst), .Q(\stack[4][0] )
         );
  DFF \stack_reg[5][0]  ( .D(n2123), .CLK(clk), .RST(rst), .Q(\stack[5][0] )
         );
  DFF \stack_reg[6][0]  ( .D(n2122), .CLK(clk), .RST(rst), .Q(\stack[6][0] )
         );
  DFF \stack_reg[7][0]  ( .D(n2121), .CLK(clk), .RST(rst), .Q(\stack[7][0] )
         );
  XOR \DP_OP_25_64_8855/U383  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_0 ), .Z(
        \DP_OP_25_64_8855/n656 ) );
  XOR \DP_OP_25_64_8855/U382  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_1 ), .Z(
        \DP_OP_25_64_8855/n655 ) );
  XOR \DP_OP_25_64_8855/U381  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_2 ), .Z(
        \DP_OP_25_64_8855/n654 ) );
  XOR \DP_OP_25_64_8855/U380  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_3 ), .Z(
        \DP_OP_25_64_8855/n653 ) );
  XOR \DP_OP_25_64_8855/U379  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_4 ), .Z(
        \DP_OP_25_64_8855/n652 ) );
  XOR \DP_OP_25_64_8855/U378  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_5 ), .Z(
        \DP_OP_25_64_8855/n651 ) );
  XOR \DP_OP_25_64_8855/U377  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_6 ), .Z(
        \DP_OP_25_64_8855/n650 ) );
  XOR \DP_OP_25_64_8855/U376  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_7 ), .Z(
        \DP_OP_25_64_8855/n649 ) );
  XOR \DP_OP_25_64_8855/U375  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_8 ), .Z(
        \DP_OP_25_64_8855/n648 ) );
  XOR \DP_OP_25_64_8855/U374  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_9 ), .Z(
        \DP_OP_25_64_8855/n647 ) );
  XOR \DP_OP_25_64_8855/U373  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_10 ), .Z(
        \DP_OP_25_64_8855/n646 ) );
  XOR \DP_OP_25_64_8855/U372  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_11 ), .Z(
        \DP_OP_25_64_8855/n645 ) );
  XOR \DP_OP_25_64_8855/U371  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_12 ), .Z(
        \DP_OP_25_64_8855/n644 ) );
  XOR \DP_OP_25_64_8855/U370  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_13 ), .Z(
        \DP_OP_25_64_8855/n643 ) );
  XOR \DP_OP_25_64_8855/U369  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_14 ), .Z(
        \DP_OP_25_64_8855/n642 ) );
  XOR \DP_OP_25_64_8855/U368  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_15 ), .Z(
        \DP_OP_25_64_8855/n641 ) );
  XOR \DP_OP_25_64_8855/U367  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_16 ), .Z(
        \DP_OP_25_64_8855/n640 ) );
  XOR \DP_OP_25_64_8855/U366  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_17 ), .Z(
        \DP_OP_25_64_8855/n639 ) );
  XOR \DP_OP_25_64_8855/U365  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_18 ), .Z(
        \DP_OP_25_64_8855/n638 ) );
  XOR \DP_OP_25_64_8855/U364  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_19 ), .Z(
        \DP_OP_25_64_8855/n637 ) );
  XOR \DP_OP_25_64_8855/U363  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_20 ), .Z(
        \DP_OP_25_64_8855/n636 ) );
  XOR \DP_OP_25_64_8855/U309  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_21 ), .Z(
        \DP_OP_25_64_8855/n635 ) );
  XOR \DP_OP_25_64_8855/U308  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_22 ), .Z(
        \DP_OP_25_64_8855/n634 ) );
  XOR \DP_OP_25_64_8855/U307  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_23 ), .Z(
        \DP_OP_25_64_8855/n633 ) );
  XOR \DP_OP_25_64_8855/U306  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_24 ), .Z(
        \DP_OP_25_64_8855/n632 ) );
  XOR \DP_OP_25_64_8855/U305  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_25 ), .Z(
        \DP_OP_25_64_8855/n631 ) );
  XOR \DP_OP_25_64_8855/U304  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_26 ), .Z(
        \DP_OP_25_64_8855/n630 ) );
  XOR \DP_OP_25_64_8855/U303  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_27 ), .Z(
        \DP_OP_25_64_8855/n629 ) );
  XOR \DP_OP_25_64_8855/U302  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_28 ), .Z(
        \DP_OP_25_64_8855/n628 ) );
  XOR \DP_OP_25_64_8855/U301  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_29 ), .Z(
        \DP_OP_25_64_8855/n627 ) );
  XOR \DP_OP_25_64_8855/U300  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_30 ), .Z(
        \DP_OP_25_64_8855/n626 ) );
  XOR \DP_OP_25_64_8855/U299  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_31 ), .Z(
        \DP_OP_25_64_8855/n625 ) );
  XOR \DP_OP_25_64_8855/U298  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_32 ), .Z(
        \DP_OP_25_64_8855/n624 ) );
  XOR \DP_OP_25_64_8855/U297  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_33 ), .Z(
        \DP_OP_25_64_8855/n623 ) );
  XOR \DP_OP_25_64_8855/U296  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_34 ), .Z(
        \DP_OP_25_64_8855/n622 ) );
  XOR \DP_OP_25_64_8855/U295  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_35 ), .Z(
        \DP_OP_25_64_8855/n621 ) );
  XOR \DP_OP_25_64_8855/U294  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_36 ), .Z(
        \DP_OP_25_64_8855/n620 ) );
  XOR \DP_OP_25_64_8855/U293  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_37 ), .Z(
        \DP_OP_25_64_8855/n619 ) );
  XOR \DP_OP_25_64_8855/U292  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_38 ), .Z(
        \DP_OP_25_64_8855/n618 ) );
  XOR \DP_OP_25_64_8855/U291  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_39 ), .Z(
        \DP_OP_25_64_8855/n617 ) );
  XOR \DP_OP_25_64_8855/U290  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_40 ), .Z(
        \DP_OP_25_64_8855/n616 ) );
  XOR \DP_OP_25_64_8855/U289  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_41 ), .Z(
        \DP_OP_25_64_8855/n615 ) );
  XOR \DP_OP_25_64_8855/U288  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_42 ), .Z(
        \DP_OP_25_64_8855/n614 ) );
  XOR \DP_OP_25_64_8855/U287  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_43 ), .Z(
        \DP_OP_25_64_8855/n613 ) );
  XOR \DP_OP_25_64_8855/U286  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_44 ), .Z(
        \DP_OP_25_64_8855/n612 ) );
  XOR \DP_OP_25_64_8855/U285  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_45 ), .Z(
        \DP_OP_25_64_8855/n611 ) );
  XOR \DP_OP_25_64_8855/U284  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_46 ), .Z(
        \DP_OP_25_64_8855/n610 ) );
  XOR \DP_OP_25_64_8855/U283  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_47 ), .Z(
        \DP_OP_25_64_8855/n609 ) );
  XOR \DP_OP_25_64_8855/U282  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_48 ), .Z(
        \DP_OP_25_64_8855/n608 ) );
  XOR \DP_OP_25_64_8855/U281  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_49 ), .Z(
        \DP_OP_25_64_8855/n607 ) );
  XOR \DP_OP_25_64_8855/U280  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_50 ), .Z(
        \DP_OP_25_64_8855/n606 ) );
  XOR \DP_OP_25_64_8855/U279  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_51 ), .Z(
        \DP_OP_25_64_8855/n605 ) );
  XOR \DP_OP_25_64_8855/U278  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_52 ), .Z(
        \DP_OP_25_64_8855/n604 ) );
  XOR \DP_OP_25_64_8855/U277  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_53 ), .Z(
        \DP_OP_25_64_8855/n603 ) );
  XOR \DP_OP_25_64_8855/U276  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_54 ), .Z(
        \DP_OP_25_64_8855/n602 ) );
  XOR \DP_OP_25_64_8855/U275  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_55 ), .Z(
        \DP_OP_25_64_8855/n601 ) );
  XOR \DP_OP_25_64_8855/U274  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_56 ), .Z(
        \DP_OP_25_64_8855/n600 ) );
  XOR \DP_OP_25_64_8855/U273  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_57 ), .Z(
        \DP_OP_25_64_8855/n599 ) );
  XOR \DP_OP_25_64_8855/U272  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_58 ), .Z(
        \DP_OP_25_64_8855/n598 ) );
  XOR \DP_OP_25_64_8855/U271  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_59 ), .Z(
        \DP_OP_25_64_8855/n597 ) );
  XOR \DP_OP_25_64_8855/U270  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_60 ), .Z(
        \DP_OP_25_64_8855/n596 ) );
  XOR \DP_OP_25_64_8855/U269  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_61 ), .Z(
        \DP_OP_25_64_8855/n595 ) );
  XOR \DP_OP_25_64_8855/U268  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_62 ), .Z(
        \DP_OP_25_64_8855/n594 ) );
  XOR \DP_OP_25_64_8855/U267  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_63 ), .Z(
        \DP_OP_25_64_8855/n593 ) );
  XOR \DP_OP_25_64_8855/U264  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_8855/n525 ) );
  XOR \DP_OP_25_64_8855/U263  ( .A(\DP_OP_25_64_8855/n525 ), .B(
        \DP_OP_25_64_8855/n656 ), .Z(\C3/DATA5_0 ) );
  XOR \DP_OP_25_64_8855/U209  ( .A(\DP_OP_25_64_8855/n655 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_8855/n524 ) );
  XOR \DP_OP_25_64_8855/U208  ( .A(\DP_OP_25_64_8855/n588 ), .B(
        \DP_OP_25_64_8855/n524 ), .Z(\C3/DATA5_1 ) );
  XOR \DP_OP_25_64_8855/U207  ( .A(\DP_OP_25_64_8855/n654 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_8855/n523 ) );
  XOR \DP_OP_25_64_8855/U206  ( .A(\DP_OP_25_64_8855/n587 ), .B(
        \DP_OP_25_64_8855/n523 ), .Z(\C3/DATA5_2 ) );
  XOR \DP_OP_25_64_8855/U205  ( .A(\DP_OP_25_64_8855/n653 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_8855/n522 ) );
  XOR \DP_OP_25_64_8855/U204  ( .A(\DP_OP_25_64_8855/n586 ), .B(
        \DP_OP_25_64_8855/n522 ), .Z(\C3/DATA5_3 ) );
  XOR \DP_OP_25_64_8855/U203  ( .A(\DP_OP_25_64_8855/n652 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_8855/n521 ) );
  XOR \DP_OP_25_64_8855/U202  ( .A(\DP_OP_25_64_8855/n585 ), .B(
        \DP_OP_25_64_8855/n521 ), .Z(\C3/DATA5_4 ) );
  XOR \DP_OP_25_64_8855/U201  ( .A(\DP_OP_25_64_8855/n651 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_8855/n520 ) );
  XOR \DP_OP_25_64_8855/U200  ( .A(\DP_OP_25_64_8855/n584 ), .B(
        \DP_OP_25_64_8855/n520 ), .Z(\C3/DATA5_5 ) );
  XOR \DP_OP_25_64_8855/U199  ( .A(\DP_OP_25_64_8855/n650 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_8855/n519 ) );
  XOR \DP_OP_25_64_8855/U198  ( .A(\DP_OP_25_64_8855/n583 ), .B(
        \DP_OP_25_64_8855/n519 ), .Z(\C3/DATA5_6 ) );
  XOR \DP_OP_25_64_8855/U197  ( .A(\DP_OP_25_64_8855/n649 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_8855/n518 ) );
  XOR \DP_OP_25_64_8855/U196  ( .A(\DP_OP_25_64_8855/n582 ), .B(
        \DP_OP_25_64_8855/n518 ), .Z(\C3/DATA5_7 ) );
  XOR \DP_OP_25_64_8855/U195  ( .A(\DP_OP_25_64_8855/n648 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_8855/n517 ) );
  XOR \DP_OP_25_64_8855/U194  ( .A(\DP_OP_25_64_8855/n581 ), .B(
        \DP_OP_25_64_8855/n517 ), .Z(\C3/DATA5_8 ) );
  XOR \DP_OP_25_64_8855/U193  ( .A(\DP_OP_25_64_8855/n647 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_8855/n516 ) );
  XOR \DP_OP_25_64_8855/U192  ( .A(\DP_OP_25_64_8855/n580 ), .B(
        \DP_OP_25_64_8855/n516 ), .Z(\C3/DATA5_9 ) );
  XOR \DP_OP_25_64_8855/U191  ( .A(\DP_OP_25_64_8855/n646 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_8855/n515 ) );
  XOR \DP_OP_25_64_8855/U190  ( .A(\DP_OP_25_64_8855/n579 ), .B(
        \DP_OP_25_64_8855/n515 ), .Z(\C3/DATA5_10 ) );
  XOR \DP_OP_25_64_8855/U189  ( .A(\DP_OP_25_64_8855/n645 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_8855/n514 ) );
  XOR \DP_OP_25_64_8855/U188  ( .A(\DP_OP_25_64_8855/n578 ), .B(
        \DP_OP_25_64_8855/n514 ), .Z(\C3/DATA5_11 ) );
  XOR \DP_OP_25_64_8855/U187  ( .A(\DP_OP_25_64_8855/n644 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_8855/n513 ) );
  XOR \DP_OP_25_64_8855/U186  ( .A(\DP_OP_25_64_8855/n577 ), .B(
        \DP_OP_25_64_8855/n513 ), .Z(\C3/DATA5_12 ) );
  XOR \DP_OP_25_64_8855/U185  ( .A(\DP_OP_25_64_8855/n643 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_8855/n512 ) );
  XOR \DP_OP_25_64_8855/U184  ( .A(\DP_OP_25_64_8855/n576 ), .B(
        \DP_OP_25_64_8855/n512 ), .Z(\C3/DATA5_13 ) );
  XOR \DP_OP_25_64_8855/U183  ( .A(\DP_OP_25_64_8855/n642 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_8855/n511 ) );
  XOR \DP_OP_25_64_8855/U182  ( .A(\DP_OP_25_64_8855/n575 ), .B(
        \DP_OP_25_64_8855/n511 ), .Z(\C3/DATA5_14 ) );
  XOR \DP_OP_25_64_8855/U181  ( .A(\DP_OP_25_64_8855/n641 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_8855/n510 ) );
  XOR \DP_OP_25_64_8855/U180  ( .A(\DP_OP_25_64_8855/n574 ), .B(
        \DP_OP_25_64_8855/n510 ), .Z(\C3/DATA5_15 ) );
  XOR \DP_OP_25_64_8855/U179  ( .A(\DP_OP_25_64_8855/n640 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_8855/n509 ) );
  XOR \DP_OP_25_64_8855/U178  ( .A(\DP_OP_25_64_8855/n573 ), .B(
        \DP_OP_25_64_8855/n509 ), .Z(\C3/DATA5_16 ) );
  XOR \DP_OP_25_64_8855/U177  ( .A(\DP_OP_25_64_8855/n639 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_8855/n508 ) );
  XOR \DP_OP_25_64_8855/U176  ( .A(\DP_OP_25_64_8855/n572 ), .B(
        \DP_OP_25_64_8855/n508 ), .Z(\C3/DATA5_17 ) );
  XOR \DP_OP_25_64_8855/U175  ( .A(\DP_OP_25_64_8855/n638 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_8855/n507 ) );
  XOR \DP_OP_25_64_8855/U174  ( .A(\DP_OP_25_64_8855/n571 ), .B(
        \DP_OP_25_64_8855/n507 ), .Z(\C3/DATA5_18 ) );
  XOR \DP_OP_25_64_8855/U173  ( .A(\DP_OP_25_64_8855/n637 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_8855/n506 ) );
  XOR \DP_OP_25_64_8855/U172  ( .A(\DP_OP_25_64_8855/n570 ), .B(
        \DP_OP_25_64_8855/n506 ), .Z(\C3/DATA5_19 ) );
  XOR \DP_OP_25_64_8855/U171  ( .A(\DP_OP_25_64_8855/n636 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_8855/n505 ) );
  XOR \DP_OP_25_64_8855/U170  ( .A(\DP_OP_25_64_8855/n569 ), .B(
        \DP_OP_25_64_8855/n505 ), .Z(\C3/DATA5_20 ) );
  XOR \DP_OP_25_64_8855/U169  ( .A(\DP_OP_25_64_8855/n635 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_8855/n504 ) );
  XOR \DP_OP_25_64_8855/U168  ( .A(\DP_OP_25_64_8855/n568 ), .B(
        \DP_OP_25_64_8855/n504 ), .Z(\C3/DATA5_21 ) );
  XOR \DP_OP_25_64_8855/U167  ( .A(\DP_OP_25_64_8855/n634 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_8855/n503 ) );
  XOR \DP_OP_25_64_8855/U166  ( .A(\DP_OP_25_64_8855/n567 ), .B(
        \DP_OP_25_64_8855/n503 ), .Z(\C3/DATA5_22 ) );
  XOR \DP_OP_25_64_8855/U165  ( .A(\DP_OP_25_64_8855/n633 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_8855/n502 ) );
  XOR \DP_OP_25_64_8855/U164  ( .A(\DP_OP_25_64_8855/n566 ), .B(
        \DP_OP_25_64_8855/n502 ), .Z(\C3/DATA5_23 ) );
  XOR \DP_OP_25_64_8855/U163  ( .A(\DP_OP_25_64_8855/n632 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_8855/n501 ) );
  XOR \DP_OP_25_64_8855/U109  ( .A(\DP_OP_25_64_8855/n565 ), .B(
        \DP_OP_25_64_8855/n501 ), .Z(\C3/DATA5_24 ) );
  XOR \DP_OP_25_64_8855/U108  ( .A(\DP_OP_25_64_8855/n631 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_8855/n500 ) );
  XOR \DP_OP_25_64_8855/U107  ( .A(\DP_OP_25_64_8855/n564 ), .B(
        \DP_OP_25_64_8855/n500 ), .Z(\C3/DATA5_25 ) );
  XOR \DP_OP_25_64_8855/U106  ( .A(\DP_OP_25_64_8855/n630 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_8855/n499 ) );
  XOR \DP_OP_25_64_8855/U105  ( .A(\DP_OP_25_64_8855/n563 ), .B(
        \DP_OP_25_64_8855/n499 ), .Z(\C3/DATA5_26 ) );
  XOR \DP_OP_25_64_8855/U104  ( .A(\DP_OP_25_64_8855/n629 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_8855/n498 ) );
  XOR \DP_OP_25_64_8855/U103  ( .A(\DP_OP_25_64_8855/n562 ), .B(
        \DP_OP_25_64_8855/n498 ), .Z(\C3/DATA5_27 ) );
  XOR \DP_OP_25_64_8855/U102  ( .A(\DP_OP_25_64_8855/n628 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_8855/n497 ) );
  XOR \DP_OP_25_64_8855/U101  ( .A(\DP_OP_25_64_8855/n561 ), .B(
        \DP_OP_25_64_8855/n497 ), .Z(\C3/DATA5_28 ) );
  XOR \DP_OP_25_64_8855/U100  ( .A(\DP_OP_25_64_8855/n627 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_8855/n496 ) );
  XOR \DP_OP_25_64_8855/U99  ( .A(\DP_OP_25_64_8855/n560 ), .B(
        \DP_OP_25_64_8855/n496 ), .Z(\C3/DATA5_29 ) );
  XOR \DP_OP_25_64_8855/U98  ( .A(\DP_OP_25_64_8855/n626 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_8855/n495 ) );
  XOR \DP_OP_25_64_8855/U97  ( .A(\DP_OP_25_64_8855/n559 ), .B(
        \DP_OP_25_64_8855/n495 ), .Z(\C3/DATA5_30 ) );
  XOR \DP_OP_25_64_8855/U96  ( .A(\DP_OP_25_64_8855/n625 ), .B(
        \U1/RSOP_16/C2/Z_31 ), .Z(\DP_OP_25_64_8855/n494 ) );
  XOR \DP_OP_25_64_8855/U95  ( .A(\DP_OP_25_64_8855/n558 ), .B(
        \DP_OP_25_64_8855/n494 ), .Z(\C3/DATA5_31 ) );
  XOR \DP_OP_25_64_8855/U94  ( .A(\DP_OP_25_64_8855/n624 ), .B(
        \U1/RSOP_16/C2/Z_32 ), .Z(\DP_OP_25_64_8855/n493 ) );
  XOR \DP_OP_25_64_8855/U93  ( .A(\DP_OP_25_64_8855/n557 ), .B(
        \DP_OP_25_64_8855/n493 ), .Z(\C3/DATA5_32 ) );
  XOR \DP_OP_25_64_8855/U92  ( .A(\DP_OP_25_64_8855/n623 ), .B(
        \U1/RSOP_16/C2/Z_33 ), .Z(\DP_OP_25_64_8855/n492 ) );
  XOR \DP_OP_25_64_8855/U91  ( .A(\DP_OP_25_64_8855/n556 ), .B(
        \DP_OP_25_64_8855/n492 ), .Z(\C3/DATA5_33 ) );
  XOR \DP_OP_25_64_8855/U90  ( .A(\DP_OP_25_64_8855/n622 ), .B(
        \U1/RSOP_16/C2/Z_34 ), .Z(\DP_OP_25_64_8855/n491 ) );
  XOR \DP_OP_25_64_8855/U89  ( .A(\DP_OP_25_64_8855/n555 ), .B(
        \DP_OP_25_64_8855/n491 ), .Z(\C3/DATA5_34 ) );
  XOR \DP_OP_25_64_8855/U88  ( .A(\DP_OP_25_64_8855/n621 ), .B(
        \U1/RSOP_16/C2/Z_35 ), .Z(\DP_OP_25_64_8855/n490 ) );
  XOR \DP_OP_25_64_8855/U87  ( .A(\DP_OP_25_64_8855/n554 ), .B(
        \DP_OP_25_64_8855/n490 ), .Z(\C3/DATA5_35 ) );
  XOR \DP_OP_25_64_8855/U86  ( .A(\DP_OP_25_64_8855/n620 ), .B(
        \U1/RSOP_16/C2/Z_36 ), .Z(\DP_OP_25_64_8855/n489 ) );
  XOR \DP_OP_25_64_8855/U85  ( .A(\DP_OP_25_64_8855/n553 ), .B(
        \DP_OP_25_64_8855/n489 ), .Z(\C3/DATA5_36 ) );
  XOR \DP_OP_25_64_8855/U84  ( .A(\DP_OP_25_64_8855/n619 ), .B(
        \U1/RSOP_16/C2/Z_37 ), .Z(\DP_OP_25_64_8855/n488 ) );
  XOR \DP_OP_25_64_8855/U83  ( .A(\DP_OP_25_64_8855/n552 ), .B(
        \DP_OP_25_64_8855/n488 ), .Z(\C3/DATA5_37 ) );
  XOR \DP_OP_25_64_8855/U82  ( .A(\DP_OP_25_64_8855/n618 ), .B(
        \U1/RSOP_16/C2/Z_38 ), .Z(\DP_OP_25_64_8855/n487 ) );
  XOR \DP_OP_25_64_8855/U81  ( .A(\DP_OP_25_64_8855/n551 ), .B(
        \DP_OP_25_64_8855/n487 ), .Z(\C3/DATA5_38 ) );
  XOR \DP_OP_25_64_8855/U80  ( .A(\DP_OP_25_64_8855/n617 ), .B(
        \U1/RSOP_16/C2/Z_39 ), .Z(\DP_OP_25_64_8855/n486 ) );
  XOR \DP_OP_25_64_8855/U79  ( .A(\DP_OP_25_64_8855/n550 ), .B(
        \DP_OP_25_64_8855/n486 ), .Z(\C3/DATA5_39 ) );
  XOR \DP_OP_25_64_8855/U78  ( .A(\DP_OP_25_64_8855/n616 ), .B(
        \U1/RSOP_16/C2/Z_40 ), .Z(\DP_OP_25_64_8855/n485 ) );
  XOR \DP_OP_25_64_8855/U77  ( .A(\DP_OP_25_64_8855/n549 ), .B(
        \DP_OP_25_64_8855/n485 ), .Z(\C3/DATA5_40 ) );
  XOR \DP_OP_25_64_8855/U76  ( .A(\DP_OP_25_64_8855/n615 ), .B(
        \U1/RSOP_16/C2/Z_41 ), .Z(\DP_OP_25_64_8855/n484 ) );
  XOR \DP_OP_25_64_8855/U75  ( .A(\DP_OP_25_64_8855/n548 ), .B(
        \DP_OP_25_64_8855/n484 ), .Z(\C3/DATA5_41 ) );
  XOR \DP_OP_25_64_8855/U74  ( .A(\DP_OP_25_64_8855/n614 ), .B(
        \U1/RSOP_16/C2/Z_42 ), .Z(\DP_OP_25_64_8855/n483 ) );
  XOR \DP_OP_25_64_8855/U73  ( .A(\DP_OP_25_64_8855/n547 ), .B(
        \DP_OP_25_64_8855/n483 ), .Z(\C3/DATA5_42 ) );
  XOR \DP_OP_25_64_8855/U72  ( .A(\DP_OP_25_64_8855/n613 ), .B(
        \U1/RSOP_16/C2/Z_43 ), .Z(\DP_OP_25_64_8855/n482 ) );
  XOR \DP_OP_25_64_8855/U71  ( .A(\DP_OP_25_64_8855/n546 ), .B(
        \DP_OP_25_64_8855/n482 ), .Z(\C3/DATA5_43 ) );
  XOR \DP_OP_25_64_8855/U70  ( .A(\DP_OP_25_64_8855/n612 ), .B(
        \U1/RSOP_16/C2/Z_44 ), .Z(\DP_OP_25_64_8855/n481 ) );
  XOR \DP_OP_25_64_8855/U69  ( .A(\DP_OP_25_64_8855/n545 ), .B(
        \DP_OP_25_64_8855/n481 ), .Z(\C3/DATA5_44 ) );
  XOR \DP_OP_25_64_8855/U68  ( .A(\DP_OP_25_64_8855/n611 ), .B(
        \U1/RSOP_16/C2/Z_45 ), .Z(\DP_OP_25_64_8855/n480 ) );
  XOR \DP_OP_25_64_8855/U67  ( .A(\DP_OP_25_64_8855/n544 ), .B(
        \DP_OP_25_64_8855/n480 ), .Z(\C3/DATA5_45 ) );
  XOR \DP_OP_25_64_8855/U66  ( .A(\DP_OP_25_64_8855/n610 ), .B(
        \U1/RSOP_16/C2/Z_46 ), .Z(\DP_OP_25_64_8855/n479 ) );
  XOR \DP_OP_25_64_8855/U65  ( .A(\DP_OP_25_64_8855/n543 ), .B(
        \DP_OP_25_64_8855/n479 ), .Z(\C3/DATA5_46 ) );
  XOR \DP_OP_25_64_8855/U64  ( .A(\DP_OP_25_64_8855/n609 ), .B(
        \U1/RSOP_16/C2/Z_47 ), .Z(\DP_OP_25_64_8855/n478 ) );
  XOR \DP_OP_25_64_8855/U63  ( .A(\DP_OP_25_64_8855/n542 ), .B(
        \DP_OP_25_64_8855/n478 ), .Z(\C3/DATA5_47 ) );
  XOR \DP_OP_25_64_8855/U62  ( .A(\DP_OP_25_64_8855/n608 ), .B(
        \U1/RSOP_16/C2/Z_48 ), .Z(\DP_OP_25_64_8855/n477 ) );
  XOR \DP_OP_25_64_8855/U61  ( .A(\DP_OP_25_64_8855/n541 ), .B(
        \DP_OP_25_64_8855/n477 ), .Z(\C3/DATA5_48 ) );
  XOR \DP_OP_25_64_8855/U60  ( .A(\DP_OP_25_64_8855/n607 ), .B(
        \U1/RSOP_16/C2/Z_49 ), .Z(\DP_OP_25_64_8855/n476 ) );
  XOR \DP_OP_25_64_8855/U59  ( .A(\DP_OP_25_64_8855/n540 ), .B(
        \DP_OP_25_64_8855/n476 ), .Z(\C3/DATA5_49 ) );
  XOR \DP_OP_25_64_8855/U58  ( .A(\DP_OP_25_64_8855/n606 ), .B(
        \U1/RSOP_16/C2/Z_50 ), .Z(\DP_OP_25_64_8855/n475 ) );
  XOR \DP_OP_25_64_8855/U57  ( .A(\DP_OP_25_64_8855/n539 ), .B(
        \DP_OP_25_64_8855/n475 ), .Z(\C3/DATA5_50 ) );
  XOR \DP_OP_25_64_8855/U56  ( .A(\DP_OP_25_64_8855/n605 ), .B(
        \U1/RSOP_16/C2/Z_51 ), .Z(\DP_OP_25_64_8855/n474 ) );
  XOR \DP_OP_25_64_8855/U55  ( .A(\DP_OP_25_64_8855/n538 ), .B(
        \DP_OP_25_64_8855/n474 ), .Z(\C3/DATA5_51 ) );
  XOR \DP_OP_25_64_8855/U54  ( .A(\DP_OP_25_64_8855/n604 ), .B(
        \U1/RSOP_16/C2/Z_52 ), .Z(\DP_OP_25_64_8855/n473 ) );
  XOR \DP_OP_25_64_8855/U53  ( .A(\DP_OP_25_64_8855/n537 ), .B(
        \DP_OP_25_64_8855/n473 ), .Z(\C3/DATA5_52 ) );
  XOR \DP_OP_25_64_8855/U52  ( .A(\DP_OP_25_64_8855/n603 ), .B(
        \U1/RSOP_16/C2/Z_53 ), .Z(\DP_OP_25_64_8855/n472 ) );
  XOR \DP_OP_25_64_8855/U51  ( .A(\DP_OP_25_64_8855/n536 ), .B(
        \DP_OP_25_64_8855/n472 ), .Z(\C3/DATA5_53 ) );
  XOR \DP_OP_25_64_8855/U50  ( .A(\DP_OP_25_64_8855/n602 ), .B(
        \U1/RSOP_16/C2/Z_54 ), .Z(\DP_OP_25_64_8855/n471 ) );
  XOR \DP_OP_25_64_8855/U49  ( .A(\DP_OP_25_64_8855/n535 ), .B(
        \DP_OP_25_64_8855/n471 ), .Z(\C3/DATA5_54 ) );
  XOR \DP_OP_25_64_8855/U48  ( .A(\DP_OP_25_64_8855/n601 ), .B(
        \U1/RSOP_16/C2/Z_55 ), .Z(\DP_OP_25_64_8855/n470 ) );
  XOR \DP_OP_25_64_8855/U47  ( .A(\DP_OP_25_64_8855/n534 ), .B(
        \DP_OP_25_64_8855/n470 ), .Z(\C3/DATA5_55 ) );
  XOR \DP_OP_25_64_8855/U46  ( .A(\DP_OP_25_64_8855/n600 ), .B(
        \U1/RSOP_16/C2/Z_56 ), .Z(\DP_OP_25_64_8855/n469 ) );
  XOR \DP_OP_25_64_8855/U45  ( .A(\DP_OP_25_64_8855/n533 ), .B(
        \DP_OP_25_64_8855/n469 ), .Z(\C3/DATA5_56 ) );
  XOR \DP_OP_25_64_8855/U44  ( .A(\DP_OP_25_64_8855/n599 ), .B(
        \U1/RSOP_16/C2/Z_57 ), .Z(\DP_OP_25_64_8855/n468 ) );
  XOR \DP_OP_25_64_8855/U43  ( .A(\DP_OP_25_64_8855/n532 ), .B(
        \DP_OP_25_64_8855/n468 ), .Z(\C3/DATA5_57 ) );
  XOR \DP_OP_25_64_8855/U42  ( .A(\DP_OP_25_64_8855/n598 ), .B(
        \U1/RSOP_16/C2/Z_58 ), .Z(\DP_OP_25_64_8855/n467 ) );
  XOR \DP_OP_25_64_8855/U41  ( .A(\DP_OP_25_64_8855/n531 ), .B(
        \DP_OP_25_64_8855/n467 ), .Z(\C3/DATA5_58 ) );
  XOR \DP_OP_25_64_8855/U40  ( .A(\DP_OP_25_64_8855/n597 ), .B(
        \U1/RSOP_16/C2/Z_59 ), .Z(\DP_OP_25_64_8855/n466 ) );
  XOR \DP_OP_25_64_8855/U30  ( .A(\DP_OP_25_64_8855/n530 ), .B(
        \DP_OP_25_64_8855/n466 ), .Z(\C3/DATA5_59 ) );
  XOR \DP_OP_25_64_8855/U20  ( .A(\DP_OP_25_64_8855/n596 ), .B(
        \U1/RSOP_16/C2/Z_60 ), .Z(\DP_OP_25_64_8855/n465 ) );
  XOR \DP_OP_25_64_8855/U10  ( .A(\DP_OP_25_64_8855/n529 ), .B(
        \DP_OP_25_64_8855/n465 ), .Z(\C3/DATA5_60 ) );
  XOR \DP_OP_25_64_8855/U9  ( .A(\DP_OP_25_64_8855/n595 ), .B(
        \U1/RSOP_16/C2/Z_61 ), .Z(\DP_OP_25_64_8855/n464 ) );
  XOR \DP_OP_25_64_8855/U8  ( .A(\DP_OP_25_64_8855/n528 ), .B(
        \DP_OP_25_64_8855/n464 ), .Z(\C3/DATA5_61 ) );
  XOR \DP_OP_25_64_8855/U7  ( .A(\DP_OP_25_64_8855/n594 ), .B(
        \U1/RSOP_16/C2/Z_62 ), .Z(\DP_OP_25_64_8855/n463 ) );
  XOR \DP_OP_25_64_8855/U6  ( .A(\DP_OP_25_64_8855/n527 ), .B(
        \DP_OP_25_64_8855/n463 ), .Z(\C3/DATA5_62 ) );
  XOR \DP_OP_25_64_8855/U5  ( .A(\DP_OP_25_64_8855/n593 ), .B(
        \U1/RSOP_16/C2/Z_63 ), .Z(\DP_OP_25_64_8855/n462 ) );
  XOR \DP_OP_25_64_8855/U4  ( .A(\DP_OP_25_64_8855/n526 ), .B(
        \DP_OP_25_64_8855/n462 ), .Z(\C3/DATA5_63 ) );
  NAND \DP_OP_25_64_8855/U162  ( .A(\DP_OP_25_64_8855/n594 ), .B(
        \U1/RSOP_16/C2/Z_62 ), .Z(\DP_OP_25_64_8855/n5 ) );
  NAND \DP_OP_25_64_8855/U262  ( .A(\DP_OP_25_64_8855/n527 ), .B(
        \DP_OP_25_64_8855/n463 ), .Z(\DP_OP_25_64_8855/n8 ) );
  NAND \DP_OP_25_64_8855/U362  ( .A(\DP_OP_25_64_8855/n5 ), .B(
        \DP_OP_25_64_8855/n8 ), .Z(\DP_OP_25_64_8855/n526 ) );
  NAND \DP_OP_25_64_8855/U161  ( .A(\DP_OP_25_64_8855/n595 ), .B(
        \U1/RSOP_16/C2/Z_61 ), .Z(\DP_OP_25_64_8855/n14 ) );
  NAND \DP_OP_25_64_8855/U261  ( .A(\DP_OP_25_64_8855/n528 ), .B(
        \DP_OP_25_64_8855/n464 ), .Z(\DP_OP_25_64_8855/n15 ) );
  NAND \DP_OP_25_64_8855/U361  ( .A(\DP_OP_25_64_8855/n14 ), .B(
        \DP_OP_25_64_8855/n15 ), .Z(\DP_OP_25_64_8855/n527 ) );
  NAND \DP_OP_25_64_8855/U160  ( .A(\DP_OP_25_64_8855/n596 ), .B(
        \U1/RSOP_16/C2/Z_60 ), .Z(\DP_OP_25_64_8855/n21 ) );
  NAND \DP_OP_25_64_8855/U260  ( .A(\DP_OP_25_64_8855/n529 ), .B(
        \DP_OP_25_64_8855/n465 ), .Z(\DP_OP_25_64_8855/n22 ) );
  NAND \DP_OP_25_64_8855/U360  ( .A(\DP_OP_25_64_8855/n21 ), .B(
        \DP_OP_25_64_8855/n22 ), .Z(\DP_OP_25_64_8855/n528 ) );
  NAND \DP_OP_25_64_8855/U159  ( .A(\DP_OP_25_64_8855/n597 ), .B(
        \U1/RSOP_16/C2/Z_59 ), .Z(\DP_OP_25_64_8855/n28 ) );
  NAND \DP_OP_25_64_8855/U259  ( .A(\DP_OP_25_64_8855/n530 ), .B(
        \DP_OP_25_64_8855/n466 ), .Z(\DP_OP_25_64_8855/n29 ) );
  NAND \DP_OP_25_64_8855/U359  ( .A(\DP_OP_25_64_8855/n28 ), .B(
        \DP_OP_25_64_8855/n29 ), .Z(\DP_OP_25_64_8855/n529 ) );
  NAND \DP_OP_25_64_8855/U158  ( .A(\DP_OP_25_64_8855/n598 ), .B(
        \U1/RSOP_16/C2/Z_58 ), .Z(\DP_OP_25_64_8855/n35 ) );
  NAND \DP_OP_25_64_8855/U258  ( .A(\DP_OP_25_64_8855/n531 ), .B(
        \DP_OP_25_64_8855/n467 ), .Z(\DP_OP_25_64_8855/n36 ) );
  NAND \DP_OP_25_64_8855/U358  ( .A(\DP_OP_25_64_8855/n35 ), .B(
        \DP_OP_25_64_8855/n36 ), .Z(\DP_OP_25_64_8855/n530 ) );
  NAND \DP_OP_25_64_8855/U157  ( .A(\DP_OP_25_64_8855/n599 ), .B(
        \U1/RSOP_16/C2/Z_57 ), .Z(\DP_OP_25_64_8855/n42 ) );
  NAND \DP_OP_25_64_8855/U257  ( .A(\DP_OP_25_64_8855/n532 ), .B(
        \DP_OP_25_64_8855/n468 ), .Z(\DP_OP_25_64_8855/n43 ) );
  NAND \DP_OP_25_64_8855/U357  ( .A(\DP_OP_25_64_8855/n42 ), .B(
        \DP_OP_25_64_8855/n43 ), .Z(\DP_OP_25_64_8855/n531 ) );
  NAND \DP_OP_25_64_8855/U156  ( .A(\DP_OP_25_64_8855/n600 ), .B(
        \U1/RSOP_16/C2/Z_56 ), .Z(\DP_OP_25_64_8855/n49 ) );
  NAND \DP_OP_25_64_8855/U256  ( .A(\DP_OP_25_64_8855/n533 ), .B(
        \DP_OP_25_64_8855/n469 ), .Z(\DP_OP_25_64_8855/n50 ) );
  NAND \DP_OP_25_64_8855/U356  ( .A(\DP_OP_25_64_8855/n49 ), .B(
        \DP_OP_25_64_8855/n50 ), .Z(\DP_OP_25_64_8855/n532 ) );
  NAND \DP_OP_25_64_8855/U155  ( .A(\DP_OP_25_64_8855/n601 ), .B(
        \U1/RSOP_16/C2/Z_55 ), .Z(\DP_OP_25_64_8855/n56 ) );
  NAND \DP_OP_25_64_8855/U255  ( .A(\DP_OP_25_64_8855/n534 ), .B(
        \DP_OP_25_64_8855/n470 ), .Z(\DP_OP_25_64_8855/n57 ) );
  NAND \DP_OP_25_64_8855/U355  ( .A(\DP_OP_25_64_8855/n56 ), .B(
        \DP_OP_25_64_8855/n57 ), .Z(\DP_OP_25_64_8855/n533 ) );
  NAND \DP_OP_25_64_8855/U154  ( .A(\DP_OP_25_64_8855/n602 ), .B(
        \U1/RSOP_16/C2/Z_54 ), .Z(\DP_OP_25_64_8855/n81 ) );
  NAND \DP_OP_25_64_8855/U254  ( .A(\DP_OP_25_64_8855/n535 ), .B(
        \DP_OP_25_64_8855/n471 ), .Z(\DP_OP_25_64_8855/n82 ) );
  NAND \DP_OP_25_64_8855/U354  ( .A(\DP_OP_25_64_8855/n81 ), .B(
        \DP_OP_25_64_8855/n82 ), .Z(\DP_OP_25_64_8855/n534 ) );
  NAND \DP_OP_25_64_8855/U153  ( .A(\DP_OP_25_64_8855/n603 ), .B(
        \U1/RSOP_16/C2/Z_53 ), .Z(\DP_OP_25_64_8855/n88 ) );
  NAND \DP_OP_25_64_8855/U253  ( .A(\DP_OP_25_64_8855/n536 ), .B(
        \DP_OP_25_64_8855/n472 ), .Z(\DP_OP_25_64_8855/n89 ) );
  NAND \DP_OP_25_64_8855/U353  ( .A(\DP_OP_25_64_8855/n88 ), .B(
        \DP_OP_25_64_8855/n89 ), .Z(\DP_OP_25_64_8855/n535 ) );
  NAND \DP_OP_25_64_8855/U152  ( .A(\DP_OP_25_64_8855/n604 ), .B(
        \U1/RSOP_16/C2/Z_52 ), .Z(\DP_OP_25_64_8855/n95 ) );
  NAND \DP_OP_25_64_8855/U252  ( .A(\DP_OP_25_64_8855/n537 ), .B(
        \DP_OP_25_64_8855/n473 ), .Z(\DP_OP_25_64_8855/n96 ) );
  NAND \DP_OP_25_64_8855/U352  ( .A(\DP_OP_25_64_8855/n95 ), .B(
        \DP_OP_25_64_8855/n96 ), .Z(\DP_OP_25_64_8855/n536 ) );
  NAND \DP_OP_25_64_8855/U151  ( .A(\DP_OP_25_64_8855/n605 ), .B(
        \U1/RSOP_16/C2/Z_51 ), .Z(\DP_OP_25_64_8855/n102 ) );
  NAND \DP_OP_25_64_8855/U251  ( .A(\DP_OP_25_64_8855/n538 ), .B(
        \DP_OP_25_64_8855/n474 ), .Z(\DP_OP_25_64_8855/n103 ) );
  NAND \DP_OP_25_64_8855/U351  ( .A(\DP_OP_25_64_8855/n102 ), .B(
        \DP_OP_25_64_8855/n103 ), .Z(\DP_OP_25_64_8855/n537 ) );
  NAND \DP_OP_25_64_8855/U150  ( .A(\DP_OP_25_64_8855/n606 ), .B(
        \U1/RSOP_16/C2/Z_50 ), .Z(\DP_OP_25_64_8855/n109 ) );
  NAND \DP_OP_25_64_8855/U250  ( .A(\DP_OP_25_64_8855/n539 ), .B(
        \DP_OP_25_64_8855/n475 ), .Z(\DP_OP_25_64_8855/n110 ) );
  NAND \DP_OP_25_64_8855/U350  ( .A(\DP_OP_25_64_8855/n109 ), .B(
        \DP_OP_25_64_8855/n110 ), .Z(\DP_OP_25_64_8855/n538 ) );
  NAND \DP_OP_25_64_8855/U149  ( .A(\DP_OP_25_64_8855/n607 ), .B(
        \U1/RSOP_16/C2/Z_49 ), .Z(\DP_OP_25_64_8855/n116 ) );
  NAND \DP_OP_25_64_8855/U249  ( .A(\DP_OP_25_64_8855/n540 ), .B(
        \DP_OP_25_64_8855/n476 ), .Z(\DP_OP_25_64_8855/n117 ) );
  NAND \DP_OP_25_64_8855/U349  ( .A(\DP_OP_25_64_8855/n116 ), .B(
        \DP_OP_25_64_8855/n117 ), .Z(\DP_OP_25_64_8855/n539 ) );
  NAND \DP_OP_25_64_8855/U148  ( .A(\DP_OP_25_64_8855/n608 ), .B(
        \U1/RSOP_16/C2/Z_48 ), .Z(\DP_OP_25_64_8855/n123 ) );
  NAND \DP_OP_25_64_8855/U248  ( .A(\DP_OP_25_64_8855/n541 ), .B(
        \DP_OP_25_64_8855/n477 ), .Z(\DP_OP_25_64_8855/n124 ) );
  NAND \DP_OP_25_64_8855/U348  ( .A(\DP_OP_25_64_8855/n123 ), .B(
        \DP_OP_25_64_8855/n124 ), .Z(\DP_OP_25_64_8855/n540 ) );
  NAND \DP_OP_25_64_8855/U147  ( .A(\DP_OP_25_64_8855/n609 ), .B(
        \U1/RSOP_16/C2/Z_47 ), .Z(\DP_OP_25_64_8855/n130 ) );
  NAND \DP_OP_25_64_8855/U247  ( .A(\DP_OP_25_64_8855/n542 ), .B(
        \DP_OP_25_64_8855/n478 ), .Z(\DP_OP_25_64_8855/n131 ) );
  NAND \DP_OP_25_64_8855/U347  ( .A(\DP_OP_25_64_8855/n130 ), .B(
        \DP_OP_25_64_8855/n131 ), .Z(\DP_OP_25_64_8855/n541 ) );
  NAND \DP_OP_25_64_8855/U146  ( .A(\DP_OP_25_64_8855/n610 ), .B(
        \U1/RSOP_16/C2/Z_46 ), .Z(\DP_OP_25_64_8855/n137 ) );
  NAND \DP_OP_25_64_8855/U246  ( .A(\DP_OP_25_64_8855/n543 ), .B(
        \DP_OP_25_64_8855/n479 ), .Z(\DP_OP_25_64_8855/n138 ) );
  NAND \DP_OP_25_64_8855/U346  ( .A(\DP_OP_25_64_8855/n137 ), .B(
        \DP_OP_25_64_8855/n138 ), .Z(\DP_OP_25_64_8855/n542 ) );
  NAND \DP_OP_25_64_8855/U145  ( .A(\DP_OP_25_64_8855/n611 ), .B(
        \U1/RSOP_16/C2/Z_45 ), .Z(\DP_OP_25_64_8855/n144 ) );
  NAND \DP_OP_25_64_8855/U245  ( .A(\DP_OP_25_64_8855/n544 ), .B(
        \DP_OP_25_64_8855/n480 ), .Z(\DP_OP_25_64_8855/n145 ) );
  NAND \DP_OP_25_64_8855/U345  ( .A(\DP_OP_25_64_8855/n144 ), .B(
        \DP_OP_25_64_8855/n145 ), .Z(\DP_OP_25_64_8855/n543 ) );
  NAND \DP_OP_25_64_8855/U144  ( .A(\DP_OP_25_64_8855/n612 ), .B(
        \U1/RSOP_16/C2/Z_44 ), .Z(\DP_OP_25_64_8855/n151 ) );
  NAND \DP_OP_25_64_8855/U244  ( .A(\DP_OP_25_64_8855/n545 ), .B(
        \DP_OP_25_64_8855/n481 ), .Z(\DP_OP_25_64_8855/n152 ) );
  NAND \DP_OP_25_64_8855/U344  ( .A(\DP_OP_25_64_8855/n151 ), .B(
        \DP_OP_25_64_8855/n152 ), .Z(\DP_OP_25_64_8855/n544 ) );
  NAND \DP_OP_25_64_8855/U143  ( .A(\DP_OP_25_64_8855/n613 ), .B(
        \U1/RSOP_16/C2/Z_43 ), .Z(\DP_OP_25_64_8855/n158 ) );
  NAND \DP_OP_25_64_8855/U243  ( .A(\DP_OP_25_64_8855/n546 ), .B(
        \DP_OP_25_64_8855/n482 ), .Z(\DP_OP_25_64_8855/n159 ) );
  NAND \DP_OP_25_64_8855/U343  ( .A(\DP_OP_25_64_8855/n158 ), .B(
        \DP_OP_25_64_8855/n159 ), .Z(\DP_OP_25_64_8855/n545 ) );
  NAND \DP_OP_25_64_8855/U142  ( .A(\DP_OP_25_64_8855/n614 ), .B(
        \U1/RSOP_16/C2/Z_42 ), .Z(\DP_OP_25_64_8855/n165 ) );
  NAND \DP_OP_25_64_8855/U242  ( .A(\DP_OP_25_64_8855/n547 ), .B(
        \DP_OP_25_64_8855/n483 ), .Z(\DP_OP_25_64_8855/n166 ) );
  NAND \DP_OP_25_64_8855/U342  ( .A(\DP_OP_25_64_8855/n165 ), .B(
        \DP_OP_25_64_8855/n166 ), .Z(\DP_OP_25_64_8855/n546 ) );
  NAND \DP_OP_25_64_8855/U141  ( .A(\DP_OP_25_64_8855/n615 ), .B(
        \U1/RSOP_16/C2/Z_41 ), .Z(\DP_OP_25_64_8855/n172 ) );
  NAND \DP_OP_25_64_8855/U241  ( .A(\DP_OP_25_64_8855/n548 ), .B(
        \DP_OP_25_64_8855/n484 ), .Z(\DP_OP_25_64_8855/n173 ) );
  NAND \DP_OP_25_64_8855/U341  ( .A(\DP_OP_25_64_8855/n172 ), .B(
        \DP_OP_25_64_8855/n173 ), .Z(\DP_OP_25_64_8855/n547 ) );
  NAND \DP_OP_25_64_8855/U140  ( .A(\DP_OP_25_64_8855/n616 ), .B(
        \U1/RSOP_16/C2/Z_40 ), .Z(\DP_OP_25_64_8855/n179 ) );
  NAND \DP_OP_25_64_8855/U240  ( .A(\DP_OP_25_64_8855/n549 ), .B(
        \DP_OP_25_64_8855/n485 ), .Z(\DP_OP_25_64_8855/n180 ) );
  NAND \DP_OP_25_64_8855/U340  ( .A(\DP_OP_25_64_8855/n179 ), .B(
        \DP_OP_25_64_8855/n180 ), .Z(\DP_OP_25_64_8855/n548 ) );
  NAND \DP_OP_25_64_8855/U139  ( .A(\DP_OP_25_64_8855/n617 ), .B(
        \U1/RSOP_16/C2/Z_39 ), .Z(\DP_OP_25_64_8855/n186 ) );
  NAND \DP_OP_25_64_8855/U239  ( .A(\DP_OP_25_64_8855/n550 ), .B(
        \DP_OP_25_64_8855/n486 ), .Z(\DP_OP_25_64_8855/n187 ) );
  NAND \DP_OP_25_64_8855/U339  ( .A(\DP_OP_25_64_8855/n186 ), .B(
        \DP_OP_25_64_8855/n187 ), .Z(\DP_OP_25_64_8855/n549 ) );
  NAND \DP_OP_25_64_8855/U138  ( .A(\DP_OP_25_64_8855/n618 ), .B(
        \U1/RSOP_16/C2/Z_38 ), .Z(\DP_OP_25_64_8855/n193 ) );
  NAND \DP_OP_25_64_8855/U238  ( .A(\DP_OP_25_64_8855/n551 ), .B(
        \DP_OP_25_64_8855/n487 ), .Z(\DP_OP_25_64_8855/n194 ) );
  NAND \DP_OP_25_64_8855/U338  ( .A(\DP_OP_25_64_8855/n193 ), .B(
        \DP_OP_25_64_8855/n194 ), .Z(\DP_OP_25_64_8855/n550 ) );
  NAND \DP_OP_25_64_8855/U137  ( .A(\DP_OP_25_64_8855/n619 ), .B(
        \U1/RSOP_16/C2/Z_37 ), .Z(\DP_OP_25_64_8855/n200 ) );
  NAND \DP_OP_25_64_8855/U237  ( .A(\DP_OP_25_64_8855/n552 ), .B(
        \DP_OP_25_64_8855/n488 ), .Z(\DP_OP_25_64_8855/n201 ) );
  NAND \DP_OP_25_64_8855/U337  ( .A(\DP_OP_25_64_8855/n200 ), .B(
        \DP_OP_25_64_8855/n201 ), .Z(\DP_OP_25_64_8855/n551 ) );
  NAND \DP_OP_25_64_8855/U136  ( .A(\DP_OP_25_64_8855/n620 ), .B(
        \U1/RSOP_16/C2/Z_36 ), .Z(\DP_OP_25_64_8855/n207 ) );
  NAND \DP_OP_25_64_8855/U236  ( .A(\DP_OP_25_64_8855/n553 ), .B(
        \DP_OP_25_64_8855/n489 ), .Z(\DP_OP_25_64_8855/n208 ) );
  NAND \DP_OP_25_64_8855/U336  ( .A(\DP_OP_25_64_8855/n207 ), .B(
        \DP_OP_25_64_8855/n208 ), .Z(\DP_OP_25_64_8855/n552 ) );
  NAND \DP_OP_25_64_8855/U135  ( .A(\DP_OP_25_64_8855/n621 ), .B(
        \U1/RSOP_16/C2/Z_35 ), .Z(\DP_OP_25_64_8855/n214 ) );
  NAND \DP_OP_25_64_8855/U235  ( .A(\DP_OP_25_64_8855/n554 ), .B(
        \DP_OP_25_64_8855/n490 ), .Z(\DP_OP_25_64_8855/n215 ) );
  NAND \DP_OP_25_64_8855/U335  ( .A(\DP_OP_25_64_8855/n214 ), .B(
        \DP_OP_25_64_8855/n215 ), .Z(\DP_OP_25_64_8855/n553 ) );
  NAND \DP_OP_25_64_8855/U134  ( .A(\DP_OP_25_64_8855/n622 ), .B(
        \U1/RSOP_16/C2/Z_34 ), .Z(\DP_OP_25_64_8855/n221 ) );
  NAND \DP_OP_25_64_8855/U234  ( .A(\DP_OP_25_64_8855/n555 ), .B(
        \DP_OP_25_64_8855/n491 ), .Z(\DP_OP_25_64_8855/n222 ) );
  NAND \DP_OP_25_64_8855/U334  ( .A(\DP_OP_25_64_8855/n221 ), .B(
        \DP_OP_25_64_8855/n222 ), .Z(\DP_OP_25_64_8855/n554 ) );
  NAND \DP_OP_25_64_8855/U133  ( .A(\DP_OP_25_64_8855/n623 ), .B(
        \U1/RSOP_16/C2/Z_33 ), .Z(\DP_OP_25_64_8855/n228 ) );
  NAND \DP_OP_25_64_8855/U233  ( .A(\DP_OP_25_64_8855/n556 ), .B(
        \DP_OP_25_64_8855/n492 ), .Z(\DP_OP_25_64_8855/n229 ) );
  NAND \DP_OP_25_64_8855/U333  ( .A(\DP_OP_25_64_8855/n228 ), .B(
        \DP_OP_25_64_8855/n229 ), .Z(\DP_OP_25_64_8855/n555 ) );
  NAND \DP_OP_25_64_8855/U132  ( .A(\DP_OP_25_64_8855/n624 ), .B(
        \U1/RSOP_16/C2/Z_32 ), .Z(\DP_OP_25_64_8855/n235 ) );
  NAND \DP_OP_25_64_8855/U232  ( .A(\DP_OP_25_64_8855/n557 ), .B(
        \DP_OP_25_64_8855/n493 ), .Z(\DP_OP_25_64_8855/n236 ) );
  NAND \DP_OP_25_64_8855/U332  ( .A(\DP_OP_25_64_8855/n235 ), .B(
        \DP_OP_25_64_8855/n236 ), .Z(\DP_OP_25_64_8855/n556 ) );
  NAND \DP_OP_25_64_8855/U131  ( .A(\DP_OP_25_64_8855/n625 ), .B(
        \U1/RSOP_16/C2/Z_31 ), .Z(\DP_OP_25_64_8855/n242 ) );
  NAND \DP_OP_25_64_8855/U231  ( .A(\DP_OP_25_64_8855/n558 ), .B(
        \DP_OP_25_64_8855/n494 ), .Z(\DP_OP_25_64_8855/n243 ) );
  NAND \DP_OP_25_64_8855/U331  ( .A(\DP_OP_25_64_8855/n242 ), .B(
        \DP_OP_25_64_8855/n243 ), .Z(\DP_OP_25_64_8855/n557 ) );
  NAND \DP_OP_25_64_8855/U130  ( .A(\DP_OP_25_64_8855/n626 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_8855/n249 ) );
  NAND \DP_OP_25_64_8855/U230  ( .A(\DP_OP_25_64_8855/n559 ), .B(
        \DP_OP_25_64_8855/n495 ), .Z(\DP_OP_25_64_8855/n250 ) );
  NAND \DP_OP_25_64_8855/U330  ( .A(\DP_OP_25_64_8855/n249 ), .B(
        \DP_OP_25_64_8855/n250 ), .Z(\DP_OP_25_64_8855/n558 ) );
  NAND \DP_OP_25_64_8855/U129  ( .A(\DP_OP_25_64_8855/n627 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_8855/n256 ) );
  NAND \DP_OP_25_64_8855/U229  ( .A(\DP_OP_25_64_8855/n560 ), .B(
        \DP_OP_25_64_8855/n496 ), .Z(\DP_OP_25_64_8855/n257 ) );
  NAND \DP_OP_25_64_8855/U329  ( .A(\DP_OP_25_64_8855/n256 ), .B(
        \DP_OP_25_64_8855/n257 ), .Z(\DP_OP_25_64_8855/n559 ) );
  NAND \DP_OP_25_64_8855/U128  ( .A(\DP_OP_25_64_8855/n628 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_8855/n263 ) );
  NAND \DP_OP_25_64_8855/U228  ( .A(\DP_OP_25_64_8855/n561 ), .B(
        \DP_OP_25_64_8855/n497 ), .Z(\DP_OP_25_64_8855/n264 ) );
  NAND \DP_OP_25_64_8855/U328  ( .A(\DP_OP_25_64_8855/n263 ), .B(
        \DP_OP_25_64_8855/n264 ), .Z(\DP_OP_25_64_8855/n560 ) );
  NAND \DP_OP_25_64_8855/U127  ( .A(\DP_OP_25_64_8855/n629 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_8855/n270 ) );
  NAND \DP_OP_25_64_8855/U227  ( .A(\DP_OP_25_64_8855/n562 ), .B(
        \DP_OP_25_64_8855/n498 ), .Z(\DP_OP_25_64_8855/n271 ) );
  NAND \DP_OP_25_64_8855/U327  ( .A(\DP_OP_25_64_8855/n270 ), .B(
        \DP_OP_25_64_8855/n271 ), .Z(\DP_OP_25_64_8855/n561 ) );
  NAND \DP_OP_25_64_8855/U126  ( .A(\DP_OP_25_64_8855/n630 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_8855/n277 ) );
  NAND \DP_OP_25_64_8855/U226  ( .A(\DP_OP_25_64_8855/n563 ), .B(
        \DP_OP_25_64_8855/n499 ), .Z(\DP_OP_25_64_8855/n278 ) );
  NAND \DP_OP_25_64_8855/U326  ( .A(\DP_OP_25_64_8855/n277 ), .B(
        \DP_OP_25_64_8855/n278 ), .Z(\DP_OP_25_64_8855/n562 ) );
  NAND \DP_OP_25_64_8855/U125  ( .A(\DP_OP_25_64_8855/n631 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_8855/n284 ) );
  NAND \DP_OP_25_64_8855/U225  ( .A(\DP_OP_25_64_8855/n564 ), .B(
        \DP_OP_25_64_8855/n500 ), .Z(\DP_OP_25_64_8855/n285 ) );
  NAND \DP_OP_25_64_8855/U325  ( .A(\DP_OP_25_64_8855/n284 ), .B(
        \DP_OP_25_64_8855/n285 ), .Z(\DP_OP_25_64_8855/n563 ) );
  NAND \DP_OP_25_64_8855/U124  ( .A(\DP_OP_25_64_8855/n632 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_8855/n291 ) );
  NAND \DP_OP_25_64_8855/U224  ( .A(\DP_OP_25_64_8855/n565 ), .B(
        \DP_OP_25_64_8855/n501 ), .Z(\DP_OP_25_64_8855/n292 ) );
  NAND \DP_OP_25_64_8855/U324  ( .A(\DP_OP_25_64_8855/n291 ), .B(
        \DP_OP_25_64_8855/n292 ), .Z(\DP_OP_25_64_8855/n564 ) );
  NAND \DP_OP_25_64_8855/U123  ( .A(\DP_OP_25_64_8855/n633 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_8855/n298 ) );
  NAND \DP_OP_25_64_8855/U223  ( .A(\DP_OP_25_64_8855/n566 ), .B(
        \DP_OP_25_64_8855/n502 ), .Z(\DP_OP_25_64_8855/n299 ) );
  NAND \DP_OP_25_64_8855/U323  ( .A(\DP_OP_25_64_8855/n298 ), .B(
        \DP_OP_25_64_8855/n299 ), .Z(\DP_OP_25_64_8855/n565 ) );
  NAND \DP_OP_25_64_8855/U122  ( .A(\DP_OP_25_64_8855/n634 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_8855/n305 ) );
  NAND \DP_OP_25_64_8855/U222  ( .A(\DP_OP_25_64_8855/n567 ), .B(
        \DP_OP_25_64_8855/n503 ), .Z(\DP_OP_25_64_8855/n306 ) );
  NAND \DP_OP_25_64_8855/U322  ( .A(\DP_OP_25_64_8855/n305 ), .B(
        \DP_OP_25_64_8855/n306 ), .Z(\DP_OP_25_64_8855/n566 ) );
  NAND \DP_OP_25_64_8855/U121  ( .A(\DP_OP_25_64_8855/n635 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_8855/n312 ) );
  NAND \DP_OP_25_64_8855/U221  ( .A(\DP_OP_25_64_8855/n568 ), .B(
        \DP_OP_25_64_8855/n504 ), .Z(\DP_OP_25_64_8855/n313 ) );
  NAND \DP_OP_25_64_8855/U321  ( .A(\DP_OP_25_64_8855/n312 ), .B(
        \DP_OP_25_64_8855/n313 ), .Z(\DP_OP_25_64_8855/n567 ) );
  NAND \DP_OP_25_64_8855/U120  ( .A(\DP_OP_25_64_8855/n636 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_8855/n319 ) );
  NAND \DP_OP_25_64_8855/U220  ( .A(\DP_OP_25_64_8855/n569 ), .B(
        \DP_OP_25_64_8855/n505 ), .Z(\DP_OP_25_64_8855/n320 ) );
  NAND \DP_OP_25_64_8855/U320  ( .A(\DP_OP_25_64_8855/n319 ), .B(
        \DP_OP_25_64_8855/n320 ), .Z(\DP_OP_25_64_8855/n568 ) );
  NAND \DP_OP_25_64_8855/U119  ( .A(\DP_OP_25_64_8855/n637 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_8855/n326 ) );
  NAND \DP_OP_25_64_8855/U219  ( .A(\DP_OP_25_64_8855/n570 ), .B(
        \DP_OP_25_64_8855/n506 ), .Z(\DP_OP_25_64_8855/n327 ) );
  NAND \DP_OP_25_64_8855/U319  ( .A(\DP_OP_25_64_8855/n326 ), .B(
        \DP_OP_25_64_8855/n327 ), .Z(\DP_OP_25_64_8855/n569 ) );
  NAND \DP_OP_25_64_8855/U118  ( .A(\DP_OP_25_64_8855/n638 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_8855/n333 ) );
  NAND \DP_OP_25_64_8855/U218  ( .A(\DP_OP_25_64_8855/n571 ), .B(
        \DP_OP_25_64_8855/n507 ), .Z(\DP_OP_25_64_8855/n334 ) );
  NAND \DP_OP_25_64_8855/U318  ( .A(\DP_OP_25_64_8855/n333 ), .B(
        \DP_OP_25_64_8855/n334 ), .Z(\DP_OP_25_64_8855/n570 ) );
  NAND \DP_OP_25_64_8855/U117  ( .A(\DP_OP_25_64_8855/n639 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_8855/n340 ) );
  NAND \DP_OP_25_64_8855/U217  ( .A(\DP_OP_25_64_8855/n572 ), .B(
        \DP_OP_25_64_8855/n508 ), .Z(\DP_OP_25_64_8855/n341 ) );
  NAND \DP_OP_25_64_8855/U317  ( .A(\DP_OP_25_64_8855/n340 ), .B(
        \DP_OP_25_64_8855/n341 ), .Z(\DP_OP_25_64_8855/n571 ) );
  NAND \DP_OP_25_64_8855/U116  ( .A(\DP_OP_25_64_8855/n640 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_8855/n347 ) );
  NAND \DP_OP_25_64_8855/U216  ( .A(\DP_OP_25_64_8855/n573 ), .B(
        \DP_OP_25_64_8855/n509 ), .Z(\DP_OP_25_64_8855/n348 ) );
  NAND \DP_OP_25_64_8855/U316  ( .A(\DP_OP_25_64_8855/n347 ), .B(
        \DP_OP_25_64_8855/n348 ), .Z(\DP_OP_25_64_8855/n572 ) );
  NAND \DP_OP_25_64_8855/U115  ( .A(\DP_OP_25_64_8855/n641 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_8855/n354 ) );
  NAND \DP_OP_25_64_8855/U215  ( .A(\DP_OP_25_64_8855/n574 ), .B(
        \DP_OP_25_64_8855/n510 ), .Z(\DP_OP_25_64_8855/n355 ) );
  NAND \DP_OP_25_64_8855/U315  ( .A(\DP_OP_25_64_8855/n354 ), .B(
        \DP_OP_25_64_8855/n355 ), .Z(\DP_OP_25_64_8855/n573 ) );
  NAND \DP_OP_25_64_8855/U114  ( .A(\DP_OP_25_64_8855/n642 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_8855/n361 ) );
  NAND \DP_OP_25_64_8855/U214  ( .A(\DP_OP_25_64_8855/n575 ), .B(
        \DP_OP_25_64_8855/n511 ), .Z(\DP_OP_25_64_8855/n362 ) );
  NAND \DP_OP_25_64_8855/U314  ( .A(\DP_OP_25_64_8855/n361 ), .B(
        \DP_OP_25_64_8855/n362 ), .Z(\DP_OP_25_64_8855/n574 ) );
  NAND \DP_OP_25_64_8855/U113  ( .A(\DP_OP_25_64_8855/n643 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_8855/n368 ) );
  NAND \DP_OP_25_64_8855/U213  ( .A(\DP_OP_25_64_8855/n576 ), .B(
        \DP_OP_25_64_8855/n512 ), .Z(\DP_OP_25_64_8855/n369 ) );
  NAND \DP_OP_25_64_8855/U313  ( .A(\DP_OP_25_64_8855/n368 ), .B(
        \DP_OP_25_64_8855/n369 ), .Z(\DP_OP_25_64_8855/n575 ) );
  NAND \DP_OP_25_64_8855/U112  ( .A(\DP_OP_25_64_8855/n644 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_8855/n375 ) );
  NAND \DP_OP_25_64_8855/U212  ( .A(\DP_OP_25_64_8855/n577 ), .B(
        \DP_OP_25_64_8855/n513 ), .Z(\DP_OP_25_64_8855/n376 ) );
  NAND \DP_OP_25_64_8855/U312  ( .A(\DP_OP_25_64_8855/n375 ), .B(
        \DP_OP_25_64_8855/n376 ), .Z(\DP_OP_25_64_8855/n576 ) );
  NAND \DP_OP_25_64_8855/U111  ( .A(\DP_OP_25_64_8855/n645 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_8855/n382 ) );
  NAND \DP_OP_25_64_8855/U211  ( .A(\DP_OP_25_64_8855/n578 ), .B(
        \DP_OP_25_64_8855/n514 ), .Z(\DP_OP_25_64_8855/n383 ) );
  NAND \DP_OP_25_64_8855/U311  ( .A(\DP_OP_25_64_8855/n382 ), .B(
        \DP_OP_25_64_8855/n383 ), .Z(\DP_OP_25_64_8855/n577 ) );
  NAND \DP_OP_25_64_8855/U110  ( .A(\DP_OP_25_64_8855/n646 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_8855/n389 ) );
  NAND \DP_OP_25_64_8855/U210  ( .A(\DP_OP_25_64_8855/n579 ), .B(
        \DP_OP_25_64_8855/n515 ), .Z(\DP_OP_25_64_8855/n390 ) );
  NAND \DP_OP_25_64_8855/U310  ( .A(\DP_OP_25_64_8855/n389 ), .B(
        \DP_OP_25_64_8855/n390 ), .Z(\DP_OP_25_64_8855/n578 ) );
  NAND \DP_OP_25_64_8855/U19  ( .A(\DP_OP_25_64_8855/n647 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_8855/n396 ) );
  NAND \DP_OP_25_64_8855/U29  ( .A(\DP_OP_25_64_8855/n580 ), .B(
        \DP_OP_25_64_8855/n516 ), .Z(\DP_OP_25_64_8855/n397 ) );
  NAND \DP_OP_25_64_8855/U39  ( .A(\DP_OP_25_64_8855/n396 ), .B(
        \DP_OP_25_64_8855/n397 ), .Z(\DP_OP_25_64_8855/n579 ) );
  NAND \DP_OP_25_64_8855/U18  ( .A(\DP_OP_25_64_8855/n648 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_8855/n403 ) );
  NAND \DP_OP_25_64_8855/U28  ( .A(\DP_OP_25_64_8855/n581 ), .B(
        \DP_OP_25_64_8855/n517 ), .Z(\DP_OP_25_64_8855/n404 ) );
  NAND \DP_OP_25_64_8855/U38  ( .A(\DP_OP_25_64_8855/n403 ), .B(
        \DP_OP_25_64_8855/n404 ), .Z(\DP_OP_25_64_8855/n580 ) );
  NAND \DP_OP_25_64_8855/U17  ( .A(\DP_OP_25_64_8855/n649 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_8855/n410 ) );
  NAND \DP_OP_25_64_8855/U27  ( .A(\DP_OP_25_64_8855/n582 ), .B(
        \DP_OP_25_64_8855/n518 ), .Z(\DP_OP_25_64_8855/n411 ) );
  NAND \DP_OP_25_64_8855/U37  ( .A(\DP_OP_25_64_8855/n410 ), .B(
        \DP_OP_25_64_8855/n411 ), .Z(\DP_OP_25_64_8855/n581 ) );
  NAND \DP_OP_25_64_8855/U16  ( .A(\DP_OP_25_64_8855/n650 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_8855/n417 ) );
  NAND \DP_OP_25_64_8855/U26  ( .A(\DP_OP_25_64_8855/n583 ), .B(
        \DP_OP_25_64_8855/n519 ), .Z(\DP_OP_25_64_8855/n418 ) );
  NAND \DP_OP_25_64_8855/U36  ( .A(\DP_OP_25_64_8855/n417 ), .B(
        \DP_OP_25_64_8855/n418 ), .Z(\DP_OP_25_64_8855/n582 ) );
  NAND \DP_OP_25_64_8855/U15  ( .A(\DP_OP_25_64_8855/n651 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_8855/n424 ) );
  NAND \DP_OP_25_64_8855/U25  ( .A(\DP_OP_25_64_8855/n584 ), .B(
        \DP_OP_25_64_8855/n520 ), .Z(\DP_OP_25_64_8855/n425 ) );
  NAND \DP_OP_25_64_8855/U35  ( .A(\DP_OP_25_64_8855/n424 ), .B(
        \DP_OP_25_64_8855/n425 ), .Z(\DP_OP_25_64_8855/n583 ) );
  NAND \DP_OP_25_64_8855/U14  ( .A(\DP_OP_25_64_8855/n652 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_8855/n431 ) );
  NAND \DP_OP_25_64_8855/U24  ( .A(\DP_OP_25_64_8855/n585 ), .B(
        \DP_OP_25_64_8855/n521 ), .Z(\DP_OP_25_64_8855/n432 ) );
  NAND \DP_OP_25_64_8855/U34  ( .A(\DP_OP_25_64_8855/n431 ), .B(
        \DP_OP_25_64_8855/n432 ), .Z(\DP_OP_25_64_8855/n584 ) );
  NAND \DP_OP_25_64_8855/U13  ( .A(\DP_OP_25_64_8855/n653 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_8855/n438 ) );
  NAND \DP_OP_25_64_8855/U23  ( .A(\DP_OP_25_64_8855/n586 ), .B(
        \DP_OP_25_64_8855/n522 ), .Z(\DP_OP_25_64_8855/n439 ) );
  NAND \DP_OP_25_64_8855/U33  ( .A(\DP_OP_25_64_8855/n438 ), .B(
        \DP_OP_25_64_8855/n439 ), .Z(\DP_OP_25_64_8855/n585 ) );
  NAND \DP_OP_25_64_8855/U12  ( .A(\DP_OP_25_64_8855/n654 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_8855/n445 ) );
  NAND \DP_OP_25_64_8855/U22  ( .A(\DP_OP_25_64_8855/n587 ), .B(
        \DP_OP_25_64_8855/n523 ), .Z(\DP_OP_25_64_8855/n446 ) );
  NAND \DP_OP_25_64_8855/U32  ( .A(\DP_OP_25_64_8855/n445 ), .B(
        \DP_OP_25_64_8855/n446 ), .Z(\DP_OP_25_64_8855/n586 ) );
  NAND \DP_OP_25_64_8855/U11  ( .A(\DP_OP_25_64_8855/n655 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_8855/n452 ) );
  NAND \DP_OP_25_64_8855/U21  ( .A(\DP_OP_25_64_8855/n588 ), .B(
        \DP_OP_25_64_8855/n524 ), .Z(\DP_OP_25_64_8855/n453 ) );
  NAND \DP_OP_25_64_8855/U31  ( .A(\DP_OP_25_64_8855/n452 ), .B(
        \DP_OP_25_64_8855/n453 ), .Z(\DP_OP_25_64_8855/n587 ) );
  NAND \DP_OP_25_64_8855/U1  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_8855/n459 ) );
  NAND \DP_OP_25_64_8855/U2  ( .A(\DP_OP_25_64_8855/n525 ), .B(
        \DP_OP_25_64_8855/n656 ), .Z(\DP_OP_25_64_8855/n460 ) );
  NAND \DP_OP_25_64_8855/U3  ( .A(\DP_OP_25_64_8855/n459 ), .B(
        \DP_OP_25_64_8855/n460 ), .Z(\DP_OP_25_64_8855/n588 ) );
  XNOR U2968 ( .A(n11882), .B(n11881), .Z(n11853) );
  XOR U2969 ( .A(n3763), .B(n3764), .Z(n3738) );
  XNOR U2970 ( .A(n13222), .B(n13221), .Z(n13193) );
  XOR U2971 ( .A(n3694), .B(n3695), .Z(n3670) );
  XNOR U2972 ( .A(n10354), .B(n10353), .Z(n10325) );
  XNOR U2973 ( .A(n11261), .B(n11260), .Z(n11232) );
  XNOR U2974 ( .A(n13904), .B(n13903), .Z(n13875) );
  XOR U2975 ( .A(n3623), .B(n3624), .Z(n3599) );
  XNOR U2976 ( .A(n7754), .B(n7753), .Z(n7745) );
  XNOR U2977 ( .A(n7572), .B(n7571), .Z(n7486) );
  XNOR U2978 ( .A(n7965), .B(n7964), .Z(n8002) );
  XNOR U2979 ( .A(n8461), .B(n8460), .Z(n8487) );
  XNOR U2980 ( .A(n8760), .B(n8759), .Z(n8678) );
  XOR U2981 ( .A(n9274), .B(n9273), .Z(n9227) );
  XNOR U2982 ( .A(n9541), .B(n9540), .Z(n9512) );
  XNOR U2983 ( .A(n9799), .B(n9798), .Z(n9770) );
  XNOR U2984 ( .A(n9192), .B(n9191), .Z(n9186) );
  XNOR U2985 ( .A(n9052), .B(n9051), .Z(n8898) );
  XNOR U2986 ( .A(n9471), .B(n9470), .Z(n9465) );
  XNOR U2987 ( .A(n10073), .B(n10072), .Z(n10044) );
  XNOR U2988 ( .A(n9595), .B(n9594), .Z(n9418) );
  XOR U2989 ( .A(n9722), .B(n9723), .Z(n9715) );
  XOR U2990 ( .A(n10378), .B(n10377), .Z(n10307) );
  XNOR U2991 ( .A(n10657), .B(n10656), .Z(n10628) );
  XNOR U2992 ( .A(n10951), .B(n10950), .Z(n10922) );
  XNOR U2993 ( .A(n10002), .B(n10003), .Z(n10124) );
  XNOR U2994 ( .A(n10162), .B(n10161), .Z(n9961) );
  XNOR U2995 ( .A(n10911), .B(n10910), .Z(n10902) );
  XNOR U2996 ( .A(n11561), .B(n11560), .Z(n11532) );
  XNOR U2997 ( .A(n11509), .B(n11508), .Z(n11500) );
  XNOR U2998 ( .A(n12212), .B(n12211), .Z(n12183) );
  XNOR U2999 ( .A(n4994), .B(n4993), .Z(n4911) );
  XNOR U3000 ( .A(n12172), .B(n12171), .Z(n12163) );
  XNOR U3001 ( .A(n12540), .B(n12539), .Z(n12511) );
  XOR U3002 ( .A(n5197), .B(n5198), .Z(n5297) );
  XNOR U3003 ( .A(n12148), .B(n12147), .Z(n12139) );
  XNOR U3004 ( .A(n12876), .B(n12875), .Z(n12847) );
  XNOR U3005 ( .A(n13182), .B(n13181), .Z(n13173) );
  XNOR U3006 ( .A(n13552), .B(n13551), .Z(n13523) );
  XNOR U3007 ( .A(n13276), .B(n13275), .Z(n13122) );
  XNOR U3008 ( .A(n13588), .B(n13587), .Z(n13592) );
  XNOR U3009 ( .A(n14259), .B(n14258), .Z(n14263) );
  XNOR U3010 ( .A(n14711), .B(n14710), .Z(n14707) );
  XOR U3011 ( .A(n4722), .B(n4723), .Z(n4628) );
  XOR U3012 ( .A(n3567), .B(n3568), .Z(n3543) );
  XNOR U3013 ( .A(n14525), .B(n14524), .Z(n14743) );
  XNOR U3014 ( .A(n14188), .B(n14187), .Z(n14179) );
  XNOR U3015 ( .A(n14514), .B(n14515), .Z(n14513) );
  XOR U3016 ( .A(n5652), .B(n5653), .Z(n5801) );
  XOR U3017 ( .A(n5005), .B(n5006), .Z(n4887) );
  XOR U3018 ( .A(n5486), .B(n5487), .Z(n5478) );
  XOR U3019 ( .A(n5310), .B(n5311), .Z(n5171) );
  XNOR U3020 ( .A(n5326), .B(n5327), .Z(n5470) );
  XNOR U3021 ( .A(n6265), .B(n6266), .Z(n6259) );
  XNOR U3022 ( .A(n6453), .B(n6454), .Z(n6447) );
  XOR U3023 ( .A(n6632), .B(n6633), .Z(n6696) );
  XNOR U3024 ( .A(n6247), .B(n6248), .Z(n6241) );
  XNOR U3025 ( .A(n6838), .B(n6839), .Z(n6898) );
  XNOR U3026 ( .A(n6856), .B(n6857), .Z(n6850) );
  XOR U3027 ( .A(n7054), .B(n7055), .Z(n7046) );
  XNOR U3028 ( .A(n7337), .B(n7336), .Z(n7266) );
  XNOR U3029 ( .A(n7791), .B(n7790), .Z(n7700) );
  XOR U3030 ( .A(n7970), .B(n7971), .Z(n7996) );
  XNOR U3031 ( .A(n5085), .B(n5086), .Z(n5079) );
  XOR U3032 ( .A(n7928), .B(n7929), .Z(n8027) );
  XNOR U3033 ( .A(n7952), .B(n7953), .Z(n8010) );
  XNOR U3034 ( .A(n4946), .B(n4947), .Z(n4940) );
  XOR U3035 ( .A(n8192), .B(n8193), .Z(n8184) );
  XOR U3036 ( .A(n8495), .B(n8496), .Z(n8452) );
  XNOR U3037 ( .A(n8508), .B(n8507), .Z(n8437) );
  XOR U3038 ( .A(n9021), .B(n9022), .Z(n8955) );
  XOR U3039 ( .A(n8138), .B(n8139), .Z(n8286) );
  XNOR U3040 ( .A(n8047), .B(n8046), .Z(n7905) );
  XOR U3041 ( .A(n7681), .B(n7682), .Z(n7673) );
  XNOR U3042 ( .A(n7456), .B(n7457), .Z(n7589) );
  XNOR U3043 ( .A(n8395), .B(n8396), .Z(n8537) );
  XNOR U3044 ( .A(n9285), .B(n9286), .Z(n9215) );
  XNOR U3045 ( .A(n9234), .B(n9233), .Z(n9273) );
  XNOR U3046 ( .A(n8940), .B(n8939), .Z(n8934) );
  XOR U3047 ( .A(n5522), .B(n5523), .Z(n5599) );
  XOR U3048 ( .A(n5221), .B(n5222), .Z(n5213) );
  XOR U3049 ( .A(n8641), .B(n8642), .Z(n8633) );
  XOR U3050 ( .A(n9203), .B(n9204), .Z(n9195) );
  XNOR U3051 ( .A(n5435), .B(n5434), .Z(n5363) );
  XNOR U3052 ( .A(n4537), .B(n4538), .Z(n4531) );
  XNOR U3053 ( .A(n9316), .B(n9315), .Z(n9150) );
  XNOR U3054 ( .A(n9453), .B(n9452), .Z(n9447) );
  XOR U3055 ( .A(n9828), .B(n9829), .Z(n9738) );
  XNOR U3056 ( .A(n9765), .B(n9764), .Z(n9756) );
  XNOR U3057 ( .A(n9816), .B(n9817), .Z(n9746) );
  XNOR U3058 ( .A(n9805), .B(n9804), .Z(n9809) );
  XNOR U3059 ( .A(n10079), .B(n10078), .Z(n10083) );
  XNOR U3060 ( .A(n4928), .B(n4929), .Z(n4922) );
  XNOR U3061 ( .A(n9835), .B(n9834), .Z(n9729) );
  XNOR U3062 ( .A(n10360), .B(n10359), .Z(n10364) );
  XOR U3063 ( .A(n9996), .B(n9997), .Z(n10130) );
  XOR U3064 ( .A(n10008), .B(n10009), .Z(n10119) );
  XNOR U3065 ( .A(n10314), .B(n10313), .Z(n10377) );
  XNOR U3066 ( .A(n10663), .B(n10662), .Z(n10667) );
  XNOR U3067 ( .A(n4301), .B(n4302), .Z(n4295) );
  XNOR U3068 ( .A(n9871), .B(n9870), .Z(n9681) );
  XOR U3069 ( .A(n10271), .B(n10272), .Z(n10406) );
  XOR U3070 ( .A(n10586), .B(n10587), .Z(n10684) );
  XNOR U3071 ( .A(n10957), .B(n10956), .Z(n10961) );
  XOR U3072 ( .A(n3909), .B(n3910), .Z(n3925) );
  XNOR U3073 ( .A(n10899), .B(n10898), .Z(n10890) );
  XNOR U3074 ( .A(n10974), .B(n10975), .Z(n10880) );
  XNOR U3075 ( .A(n11285), .B(n11284), .Z(n11206) );
  XNOR U3076 ( .A(n11267), .B(n11266), .Z(n11271) );
  XNOR U3077 ( .A(n11567), .B(n11566), .Z(n11571) );
  XOR U3078 ( .A(n4650), .B(n4651), .Z(n4643) );
  XNOR U3079 ( .A(n11888), .B(n11887), .Z(n11892) );
  XNOR U3080 ( .A(n10444), .B(n10443), .Z(n10230) );
  XNOR U3081 ( .A(n4845), .B(n4844), .Z(n4773) );
  XNOR U3082 ( .A(n4519), .B(n4520), .Z(n4579) );
  XOR U3083 ( .A(n11496), .B(n11497), .Z(n11594) );
  XNOR U3084 ( .A(n11585), .B(n11584), .Z(n11589) );
  XNOR U3085 ( .A(n11912), .B(n11911), .Z(n11916) );
  XOR U3086 ( .A(n10527), .B(n10528), .Z(n10745) );
  XOR U3087 ( .A(n4401), .B(n4402), .Z(n4396) );
  XOR U3088 ( .A(n4233), .B(n4234), .Z(n4185) );
  XNOR U3089 ( .A(n12218), .B(n12217), .Z(n12222) );
  XNOR U3090 ( .A(n12546), .B(n12545), .Z(n12550) );
  XOR U3091 ( .A(n12135), .B(n12136), .Z(n12245) );
  XNOR U3092 ( .A(n12564), .B(n12563), .Z(n12568) );
  XNOR U3093 ( .A(n12882), .B(n12881), .Z(n12886) );
  XNOR U3094 ( .A(n12836), .B(n12835), .Z(n12827) );
  XNOR U3095 ( .A(n5140), .B(n5139), .Z(n5044) );
  XOR U3096 ( .A(n4126), .B(n4127), .Z(n4079) );
  XNOR U3097 ( .A(n12451), .B(n12452), .Z(n12593) );
  XNOR U3098 ( .A(n13228), .B(n13227), .Z(n13232) );
  XNOR U3099 ( .A(n17180), .B(n4029), .Z(n3982) );
  XOR U3100 ( .A(n12781), .B(n12782), .Z(n12773) );
  XNOR U3101 ( .A(n12912), .B(n12911), .Z(n12916) );
  XNOR U3102 ( .A(n13258), .B(n13257), .Z(n13156) );
  XNOR U3103 ( .A(n13576), .B(n13575), .Z(n13580) );
  XNOR U3104 ( .A(n13558), .B(n13557), .Z(n13562) );
  XNOR U3105 ( .A(n13910), .B(n13909), .Z(n13914) );
  XNOR U3106 ( .A(n5191), .B(n5192), .Z(n5302) );
  XOR U3107 ( .A(n4180), .B(n4181), .Z(n4243) );
  XNOR U3108 ( .A(n13928), .B(n13927), .Z(n13932) );
  XNOR U3109 ( .A(n14253), .B(n14252), .Z(n14223) );
  XOR U3110 ( .A(n4585), .B(n4586), .Z(n4502) );
  XOR U3111 ( .A(n3933), .B(n3934), .Z(n3886) );
  XNOR U3112 ( .A(n13482), .B(n13481), .Z(n13473) );
  XNOR U3113 ( .A(n13955), .B(n13956), .Z(n13958) );
  XNOR U3114 ( .A(n13940), .B(n13939), .Z(n13944) );
  XNOR U3115 ( .A(n14212), .B(n14211), .Z(n14203) );
  XOR U3116 ( .A(n5037), .B(n5038), .Z(n5149) );
  XOR U3117 ( .A(n3853), .B(n3854), .Z(n3806) );
  XNOR U3118 ( .A(n13618), .B(n13617), .Z(n13452) );
  XNOR U3119 ( .A(n14289), .B(n14288), .Z(n14293) );
  XNOR U3120 ( .A(n14687), .B(n14686), .Z(n14536) );
  XOR U3121 ( .A(n5492), .B(n5493), .Z(n5629) );
  XOR U3122 ( .A(n13809), .B(n13810), .Z(n13980) );
  XOR U3123 ( .A(n14175), .B(n14176), .Z(n14322) );
  XNOR U3124 ( .A(n14759), .B(n14758), .Z(n14785) );
  XNOR U3125 ( .A(n14795), .B(n14794), .Z(n14508) );
  XOR U3126 ( .A(n4856), .B(n4857), .Z(n4749) );
  XOR U3127 ( .A(n3769), .B(n3770), .Z(n3721) );
  XOR U3128 ( .A(n3508), .B(n3509), .Z(n3484) );
  XOR U3129 ( .A(n5332), .B(n5333), .Z(n5324) );
  XOR U3130 ( .A(n4271), .B(n4272), .Z(n4359) );
  XOR U3131 ( .A(n4168), .B(n4169), .Z(n4163) );
  XOR U3132 ( .A(n3700), .B(n3701), .Z(n3654) );
  XNOR U3133 ( .A(n17338), .B(n3465), .Z(n3441) );
  XOR U3134 ( .A(n5025), .B(n5026), .Z(n5020) );
  XOR U3135 ( .A(n3629), .B(n3630), .Z(n3582) );
  XOR U3136 ( .A(n3417), .B(n3418), .Z(n3394) );
  XOR U3137 ( .A(n14065), .B(n14066), .Z(n13719) );
  XOR U3138 ( .A(n13359), .B(n13360), .Z(n13025) );
  XOR U3139 ( .A(n12677), .B(n12678), .Z(n12355) );
  XOR U3140 ( .A(n12019), .B(n12020), .Z(n11710) );
  XOR U3141 ( .A(n11386), .B(n11387), .Z(n11088) );
  XOR U3142 ( .A(n10776), .B(n10777), .Z(n10491) );
  XOR U3143 ( .A(n10191), .B(n10192), .Z(n9918) );
  XOR U3144 ( .A(n9630), .B(n9631), .Z(n9369) );
  XOR U3145 ( .A(n9093), .B(n9094), .Z(n8843) );
  XOR U3146 ( .A(n8579), .B(n8580), .Z(n8341) );
  XOR U3147 ( .A(n8088), .B(n8089), .Z(n7862) );
  XOR U3148 ( .A(n7625), .B(n7626), .Z(n7408) );
  XOR U3149 ( .A(n7179), .B(n7180), .Z(n6976) );
  XOR U3150 ( .A(n6758), .B(n6759), .Z(n6567) );
  XOR U3151 ( .A(n6361), .B(n6362), .Z(n6181) );
  XOR U3152 ( .A(n5646), .B(n5647), .Z(n5806) );
  XNOR U3153 ( .A(n5480), .B(n5481), .Z(n5636) );
  XOR U3154 ( .A(n4490), .B(n4489), .Z(n4601) );
  XOR U3155 ( .A(n3573), .B(n3574), .Z(n3526) );
  XOR U3156 ( .A(n3379), .B(n3380), .Z(n3356) );
  XOR U3157 ( .A(n5167), .B(n5168), .Z(n5161) );
  XOR U3158 ( .A(n4479), .B(n4480), .Z(n4365) );
  XOR U3159 ( .A(n3429), .B(n3430), .Z(n3421) );
  IV U3160 ( .A(n17471), .Z(n2967) );
  IV U3161 ( .A(\stack[1][0] ), .Z(n2968) );
  IV U3162 ( .A(\stack[1][1] ), .Z(n2969) );
  IV U3163 ( .A(\stack[1][2] ), .Z(n2970) );
  IV U3164 ( .A(\stack[1][4] ), .Z(n2971) );
  IV U3165 ( .A(\stack[1][11] ), .Z(n2972) );
  IV U3166 ( .A(\stack[1][12] ), .Z(n2973) );
  IV U3167 ( .A(\stack[1][13] ), .Z(n2974) );
  IV U3168 ( .A(\stack[1][14] ), .Z(n2975) );
  IV U3169 ( .A(\stack[1][15] ), .Z(n2976) );
  IV U3170 ( .A(\stack[1][16] ), .Z(n2977) );
  IV U3171 ( .A(\stack[1][21] ), .Z(n2978) );
  IV U3172 ( .A(\stack[1][22] ), .Z(n2979) );
  IV U3173 ( .A(\stack[1][23] ), .Z(n2980) );
  IV U3174 ( .A(\stack[1][24] ), .Z(n2981) );
  IV U3175 ( .A(\stack[1][25] ), .Z(n2982) );
  IV U3176 ( .A(\stack[1][26] ), .Z(n2983) );
  IV U3177 ( .A(\stack[1][27] ), .Z(n2984) );
  IV U3178 ( .A(\stack[1][28] ), .Z(n2985) );
  IV U3179 ( .A(\stack[1][29] ), .Z(n2986) );
  IV U3180 ( .A(\stack[1][30] ), .Z(n2987) );
  IV U3181 ( .A(\stack[1][31] ), .Z(n2988) );
  IV U3182 ( .A(\stack[1][32] ), .Z(n2989) );
  IV U3183 ( .A(\stack[1][33] ), .Z(n2990) );
  IV U3184 ( .A(\stack[1][34] ), .Z(n2991) );
  IV U3185 ( .A(\stack[1][35] ), .Z(n2992) );
  IV U3186 ( .A(\stack[1][36] ), .Z(n2993) );
  IV U3187 ( .A(o[0]), .Z(n2994) );
  IV U3188 ( .A(o[1]), .Z(n2995) );
  IV U3189 ( .A(o[2]), .Z(n2996) );
  IV U3190 ( .A(o[3]), .Z(n2997) );
  IV U3191 ( .A(o[4]), .Z(n2998) );
  IV U3192 ( .A(o[5]), .Z(n2999) );
  IV U3193 ( .A(o[6]), .Z(n3000) );
  IV U3194 ( .A(o[7]), .Z(n3001) );
  IV U3195 ( .A(o[8]), .Z(n3002) );
  IV U3196 ( .A(o[9]), .Z(n3003) );
  IV U3197 ( .A(o[10]), .Z(n3004) );
  IV U3198 ( .A(o[11]), .Z(n3005) );
  IV U3199 ( .A(o[12]), .Z(n3006) );
  IV U3200 ( .A(o[13]), .Z(n3007) );
  IV U3201 ( .A(o[14]), .Z(n3008) );
  IV U3202 ( .A(o[15]), .Z(n3009) );
  IV U3203 ( .A(o[16]), .Z(n3010) );
  IV U3204 ( .A(o[17]), .Z(n3011) );
  IV U3205 ( .A(o[18]), .Z(n3012) );
  IV U3206 ( .A(o[19]), .Z(n3013) );
  IV U3207 ( .A(o[20]), .Z(n3014) );
  IV U3208 ( .A(o[21]), .Z(n3015) );
  IV U3209 ( .A(o[22]), .Z(n3016) );
  IV U3210 ( .A(o[23]), .Z(n3017) );
  IV U3211 ( .A(o[24]), .Z(n3018) );
  IV U3212 ( .A(o[25]), .Z(n3019) );
  IV U3213 ( .A(o[26]), .Z(n3020) );
  IV U3214 ( .A(o[28]), .Z(n3021) );
  IV U3215 ( .A(opcode[0]), .Z(n3221) );
  ANDN U3216 ( .B(opcode[0]), .A(opcode[1]), .Z(n3153) );
  ANDN U3217 ( .B(n3153), .A(opcode[2]), .Z(n3219) );
  IV U3218 ( .A(opcode[2]), .Z(n3220) );
  NANDN U3219 ( .A(opcode[0]), .B(opcode[1]), .Z(n15051) );
  OR U3220 ( .A(opcode[2]), .B(n15051), .Z(n3152) );
  NANDN U3221 ( .A(n3219), .B(n3152), .Z(n3148) );
  AND U3222 ( .A(o[63]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_63 ) );
  AND U3223 ( .A(o[62]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_62 ) );
  AND U3224 ( .A(o[61]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_61 ) );
  AND U3225 ( .A(o[60]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_60 ) );
  AND U3226 ( .A(o[59]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_59 ) );
  AND U3227 ( .A(o[58]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_58 ) );
  AND U3228 ( .A(o[57]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_57 ) );
  AND U3229 ( .A(o[56]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_56 ) );
  AND U3230 ( .A(o[55]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_55 ) );
  AND U3231 ( .A(o[54]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_54 ) );
  AND U3232 ( .A(o[53]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_53 ) );
  AND U3233 ( .A(o[52]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_52 ) );
  AND U3234 ( .A(o[51]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_51 ) );
  AND U3235 ( .A(o[50]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_50 ) );
  AND U3236 ( .A(o[49]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_49 ) );
  AND U3237 ( .A(o[48]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_48 ) );
  AND U3238 ( .A(o[47]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_47 ) );
  AND U3239 ( .A(o[46]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_46 ) );
  AND U3240 ( .A(o[45]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_45 ) );
  AND U3241 ( .A(o[44]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_44 ) );
  AND U3242 ( .A(o[43]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_43 ) );
  AND U3243 ( .A(o[42]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_42 ) );
  AND U3244 ( .A(o[41]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_41 ) );
  AND U3245 ( .A(o[40]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_40 ) );
  AND U3246 ( .A(o[39]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_39 ) );
  AND U3247 ( .A(o[38]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_38 ) );
  AND U3248 ( .A(o[37]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_37 ) );
  AND U3249 ( .A(o[36]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_36 ) );
  AND U3250 ( .A(o[35]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_35 ) );
  AND U3251 ( .A(o[34]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_34 ) );
  AND U3252 ( .A(o[33]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_33 ) );
  AND U3253 ( .A(o[32]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_32 ) );
  AND U3254 ( .A(o[31]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_31 ) );
  AND U3255 ( .A(o[30]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_30 ) );
  AND U3256 ( .A(o[29]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_29 ) );
  AND U3257 ( .A(o[28]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_28 ) );
  AND U3258 ( .A(o[27]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_27 ) );
  AND U3259 ( .A(o[26]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_26 ) );
  AND U3260 ( .A(o[25]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_25 ) );
  AND U3261 ( .A(o[24]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_24 ) );
  AND U3262 ( .A(o[23]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_23 ) );
  AND U3263 ( .A(o[22]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_22 ) );
  AND U3264 ( .A(o[21]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_21 ) );
  AND U3265 ( .A(o[20]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_20 ) );
  AND U3266 ( .A(o[19]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_19 ) );
  AND U3267 ( .A(o[18]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_18 ) );
  AND U3268 ( .A(o[17]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_17 ) );
  AND U3269 ( .A(o[16]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_16 ) );
  AND U3270 ( .A(o[15]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_15 ) );
  AND U3271 ( .A(o[14]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_14 ) );
  AND U3272 ( .A(o[13]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_13 ) );
  AND U3273 ( .A(o[12]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_12 ) );
  AND U3274 ( .A(o[11]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_11 ) );
  AND U3275 ( .A(o[10]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_10 ) );
  AND U3276 ( .A(o[9]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_9 ) );
  AND U3277 ( .A(o[8]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_8 ) );
  AND U3278 ( .A(o[7]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_7 ) );
  AND U3279 ( .A(o[6]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_6 ) );
  AND U3280 ( .A(o[5]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_5 ) );
  AND U3281 ( .A(o[4]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_4 ) );
  AND U3282 ( .A(o[3]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_3 ) );
  AND U3283 ( .A(o[2]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_2 ) );
  AND U3284 ( .A(o[1]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_1 ) );
  AND U3285 ( .A(o[0]), .B(n3148), .Z(\U1/RSOP_16/C2/Z_0 ) );
  AND U3286 ( .A(n3153), .B(opcode[2]), .Z(n3151) );
  NAND U3287 ( .A(n3151), .B(o[63]), .Z(n3023) );
  NAND U3288 ( .A(\stack[1][63] ), .B(n3148), .Z(n3022) );
  NAND U3289 ( .A(n3023), .B(n3022), .Z(\U1/RSOP_16/C3/Z_63 ) );
  NAND U3290 ( .A(n3151), .B(o[62]), .Z(n3025) );
  NAND U3291 ( .A(\stack[1][62] ), .B(n3148), .Z(n3024) );
  NAND U3292 ( .A(n3025), .B(n3024), .Z(\U1/RSOP_16/C3/Z_62 ) );
  NAND U3293 ( .A(n3151), .B(o[61]), .Z(n3027) );
  NAND U3294 ( .A(\stack[1][61] ), .B(n3148), .Z(n3026) );
  NAND U3295 ( .A(n3027), .B(n3026), .Z(\U1/RSOP_16/C3/Z_61 ) );
  NAND U3296 ( .A(n3151), .B(o[60]), .Z(n3029) );
  NAND U3297 ( .A(\stack[1][60] ), .B(n3148), .Z(n3028) );
  NAND U3298 ( .A(n3029), .B(n3028), .Z(\U1/RSOP_16/C3/Z_60 ) );
  NAND U3299 ( .A(n3151), .B(o[59]), .Z(n3031) );
  NAND U3300 ( .A(\stack[1][59] ), .B(n3148), .Z(n3030) );
  NAND U3301 ( .A(n3031), .B(n3030), .Z(\U1/RSOP_16/C3/Z_59 ) );
  NAND U3302 ( .A(n3151), .B(o[58]), .Z(n3033) );
  NAND U3303 ( .A(\stack[1][58] ), .B(n3148), .Z(n3032) );
  NAND U3304 ( .A(n3033), .B(n3032), .Z(\U1/RSOP_16/C3/Z_58 ) );
  NAND U3305 ( .A(n3151), .B(o[57]), .Z(n3035) );
  NAND U3306 ( .A(\stack[1][57] ), .B(n3148), .Z(n3034) );
  NAND U3307 ( .A(n3035), .B(n3034), .Z(\U1/RSOP_16/C3/Z_57 ) );
  NAND U3308 ( .A(n3151), .B(o[56]), .Z(n3037) );
  NAND U3309 ( .A(\stack[1][56] ), .B(n3148), .Z(n3036) );
  NAND U3310 ( .A(n3037), .B(n3036), .Z(\U1/RSOP_16/C3/Z_56 ) );
  NAND U3311 ( .A(n3151), .B(o[55]), .Z(n3039) );
  NAND U3312 ( .A(\stack[1][55] ), .B(n3148), .Z(n3038) );
  NAND U3313 ( .A(n3039), .B(n3038), .Z(\U1/RSOP_16/C3/Z_55 ) );
  NAND U3314 ( .A(n3151), .B(o[54]), .Z(n3041) );
  NAND U3315 ( .A(\stack[1][54] ), .B(n3148), .Z(n3040) );
  NAND U3316 ( .A(n3041), .B(n3040), .Z(\U1/RSOP_16/C3/Z_54 ) );
  NAND U3317 ( .A(n3151), .B(o[53]), .Z(n3043) );
  NAND U3318 ( .A(\stack[1][53] ), .B(n3148), .Z(n3042) );
  NAND U3319 ( .A(n3043), .B(n3042), .Z(\U1/RSOP_16/C3/Z_53 ) );
  NAND U3320 ( .A(n3151), .B(o[52]), .Z(n3045) );
  NAND U3321 ( .A(\stack[1][52] ), .B(n3148), .Z(n3044) );
  NAND U3322 ( .A(n3045), .B(n3044), .Z(\U1/RSOP_16/C3/Z_52 ) );
  NAND U3323 ( .A(n3151), .B(o[51]), .Z(n3047) );
  NAND U3324 ( .A(\stack[1][51] ), .B(n3148), .Z(n3046) );
  NAND U3325 ( .A(n3047), .B(n3046), .Z(\U1/RSOP_16/C3/Z_51 ) );
  NAND U3326 ( .A(n3151), .B(o[50]), .Z(n3049) );
  NAND U3327 ( .A(\stack[1][50] ), .B(n3148), .Z(n3048) );
  NAND U3328 ( .A(n3049), .B(n3048), .Z(\U1/RSOP_16/C3/Z_50 ) );
  NAND U3329 ( .A(n3151), .B(o[49]), .Z(n3051) );
  NAND U3330 ( .A(\stack[1][49] ), .B(n3148), .Z(n3050) );
  NAND U3331 ( .A(n3051), .B(n3050), .Z(\U1/RSOP_16/C3/Z_49 ) );
  NAND U3332 ( .A(n3151), .B(o[48]), .Z(n3053) );
  NAND U3333 ( .A(\stack[1][48] ), .B(n3148), .Z(n3052) );
  NAND U3334 ( .A(n3053), .B(n3052), .Z(\U1/RSOP_16/C3/Z_48 ) );
  NAND U3335 ( .A(n3151), .B(o[47]), .Z(n3055) );
  NAND U3336 ( .A(\stack[1][47] ), .B(n3148), .Z(n3054) );
  NAND U3337 ( .A(n3055), .B(n3054), .Z(\U1/RSOP_16/C3/Z_47 ) );
  NAND U3338 ( .A(n3151), .B(o[46]), .Z(n3057) );
  NAND U3339 ( .A(\stack[1][46] ), .B(n3148), .Z(n3056) );
  NAND U3340 ( .A(n3057), .B(n3056), .Z(\U1/RSOP_16/C3/Z_46 ) );
  NAND U3341 ( .A(n3151), .B(o[45]), .Z(n3059) );
  NAND U3342 ( .A(\stack[1][45] ), .B(n3148), .Z(n3058) );
  NAND U3343 ( .A(n3059), .B(n3058), .Z(\U1/RSOP_16/C3/Z_45 ) );
  NAND U3344 ( .A(n3151), .B(o[44]), .Z(n3061) );
  NAND U3345 ( .A(\stack[1][44] ), .B(n3148), .Z(n3060) );
  NAND U3346 ( .A(n3061), .B(n3060), .Z(\U1/RSOP_16/C3/Z_44 ) );
  NAND U3347 ( .A(n3151), .B(o[43]), .Z(n3063) );
  NAND U3348 ( .A(\stack[1][43] ), .B(n3148), .Z(n3062) );
  NAND U3349 ( .A(n3063), .B(n3062), .Z(\U1/RSOP_16/C3/Z_43 ) );
  NAND U3350 ( .A(n3151), .B(o[42]), .Z(n3065) );
  NAND U3351 ( .A(\stack[1][42] ), .B(n3148), .Z(n3064) );
  NAND U3352 ( .A(n3065), .B(n3064), .Z(\U1/RSOP_16/C3/Z_42 ) );
  NAND U3353 ( .A(n3151), .B(o[41]), .Z(n3067) );
  NAND U3354 ( .A(\stack[1][41] ), .B(n3148), .Z(n3066) );
  NAND U3355 ( .A(n3067), .B(n3066), .Z(\U1/RSOP_16/C3/Z_41 ) );
  NAND U3356 ( .A(n3151), .B(o[40]), .Z(n3069) );
  NAND U3357 ( .A(\stack[1][40] ), .B(n3148), .Z(n3068) );
  NAND U3358 ( .A(n3069), .B(n3068), .Z(\U1/RSOP_16/C3/Z_40 ) );
  NAND U3359 ( .A(n3151), .B(o[39]), .Z(n3071) );
  NAND U3360 ( .A(\stack[1][39] ), .B(n3148), .Z(n3070) );
  NAND U3361 ( .A(n3071), .B(n3070), .Z(\U1/RSOP_16/C3/Z_39 ) );
  NAND U3362 ( .A(n3151), .B(o[38]), .Z(n3073) );
  NAND U3363 ( .A(\stack[1][38] ), .B(n3148), .Z(n3072) );
  NAND U3364 ( .A(n3073), .B(n3072), .Z(\U1/RSOP_16/C3/Z_38 ) );
  NAND U3365 ( .A(n3151), .B(o[37]), .Z(n3075) );
  NAND U3366 ( .A(\stack[1][37] ), .B(n3148), .Z(n3074) );
  NAND U3367 ( .A(n3075), .B(n3074), .Z(\U1/RSOP_16/C3/Z_37 ) );
  NAND U3368 ( .A(n3151), .B(o[36]), .Z(n3077) );
  NAND U3369 ( .A(\stack[1][36] ), .B(n3148), .Z(n3076) );
  NAND U3370 ( .A(n3077), .B(n3076), .Z(\U1/RSOP_16/C3/Z_36 ) );
  NAND U3371 ( .A(n3151), .B(o[35]), .Z(n3079) );
  NAND U3372 ( .A(\stack[1][35] ), .B(n3148), .Z(n3078) );
  NAND U3373 ( .A(n3079), .B(n3078), .Z(\U1/RSOP_16/C3/Z_35 ) );
  NAND U3374 ( .A(n3151), .B(o[34]), .Z(n3081) );
  NAND U3375 ( .A(\stack[1][34] ), .B(n3148), .Z(n3080) );
  NAND U3376 ( .A(n3081), .B(n3080), .Z(\U1/RSOP_16/C3/Z_34 ) );
  NAND U3377 ( .A(n3151), .B(o[33]), .Z(n3083) );
  NAND U3378 ( .A(\stack[1][33] ), .B(n3148), .Z(n3082) );
  NAND U3379 ( .A(n3083), .B(n3082), .Z(\U1/RSOP_16/C3/Z_33 ) );
  NAND U3380 ( .A(n3151), .B(o[32]), .Z(n3085) );
  NAND U3381 ( .A(\stack[1][32] ), .B(n3148), .Z(n3084) );
  NAND U3382 ( .A(n3085), .B(n3084), .Z(\U1/RSOP_16/C3/Z_32 ) );
  NAND U3383 ( .A(n3151), .B(o[31]), .Z(n3087) );
  NAND U3384 ( .A(\stack[1][31] ), .B(n3148), .Z(n3086) );
  NAND U3385 ( .A(n3087), .B(n3086), .Z(\U1/RSOP_16/C3/Z_31 ) );
  NAND U3386 ( .A(n3151), .B(o[30]), .Z(n3089) );
  NAND U3387 ( .A(\stack[1][30] ), .B(n3148), .Z(n3088) );
  NAND U3388 ( .A(n3089), .B(n3088), .Z(\U1/RSOP_16/C3/Z_30 ) );
  NAND U3389 ( .A(n3151), .B(o[29]), .Z(n3091) );
  NAND U3390 ( .A(\stack[1][29] ), .B(n3148), .Z(n3090) );
  NAND U3391 ( .A(n3091), .B(n3090), .Z(\U1/RSOP_16/C3/Z_29 ) );
  NAND U3392 ( .A(n3151), .B(o[28]), .Z(n3093) );
  NAND U3393 ( .A(\stack[1][28] ), .B(n3148), .Z(n3092) );
  NAND U3394 ( .A(n3093), .B(n3092), .Z(\U1/RSOP_16/C3/Z_28 ) );
  NAND U3395 ( .A(n3151), .B(o[27]), .Z(n3095) );
  NAND U3396 ( .A(\stack[1][27] ), .B(n3148), .Z(n3094) );
  NAND U3397 ( .A(n3095), .B(n3094), .Z(\U1/RSOP_16/C3/Z_27 ) );
  NAND U3398 ( .A(n3151), .B(o[26]), .Z(n3097) );
  NAND U3399 ( .A(\stack[1][26] ), .B(n3148), .Z(n3096) );
  NAND U3400 ( .A(n3097), .B(n3096), .Z(\U1/RSOP_16/C3/Z_26 ) );
  NAND U3401 ( .A(n3151), .B(o[25]), .Z(n3099) );
  NAND U3402 ( .A(\stack[1][25] ), .B(n3148), .Z(n3098) );
  NAND U3403 ( .A(n3099), .B(n3098), .Z(\U1/RSOP_16/C3/Z_25 ) );
  NAND U3404 ( .A(n3151), .B(o[24]), .Z(n3101) );
  NAND U3405 ( .A(\stack[1][24] ), .B(n3148), .Z(n3100) );
  NAND U3406 ( .A(n3101), .B(n3100), .Z(\U1/RSOP_16/C3/Z_24 ) );
  NAND U3407 ( .A(n3151), .B(o[23]), .Z(n3103) );
  NAND U3408 ( .A(\stack[1][23] ), .B(n3148), .Z(n3102) );
  NAND U3409 ( .A(n3103), .B(n3102), .Z(\U1/RSOP_16/C3/Z_23 ) );
  NAND U3410 ( .A(n3151), .B(o[22]), .Z(n3105) );
  NAND U3411 ( .A(\stack[1][22] ), .B(n3148), .Z(n3104) );
  NAND U3412 ( .A(n3105), .B(n3104), .Z(\U1/RSOP_16/C3/Z_22 ) );
  NAND U3413 ( .A(n3151), .B(o[21]), .Z(n3107) );
  NAND U3414 ( .A(\stack[1][21] ), .B(n3148), .Z(n3106) );
  NAND U3415 ( .A(n3107), .B(n3106), .Z(\U1/RSOP_16/C3/Z_21 ) );
  NAND U3416 ( .A(n3151), .B(o[20]), .Z(n3109) );
  NAND U3417 ( .A(\stack[1][20] ), .B(n3148), .Z(n3108) );
  NAND U3418 ( .A(n3109), .B(n3108), .Z(\U1/RSOP_16/C3/Z_20 ) );
  NAND U3419 ( .A(n3151), .B(o[19]), .Z(n3111) );
  NAND U3420 ( .A(\stack[1][19] ), .B(n3148), .Z(n3110) );
  NAND U3421 ( .A(n3111), .B(n3110), .Z(\U1/RSOP_16/C3/Z_19 ) );
  NAND U3422 ( .A(n3151), .B(o[18]), .Z(n3113) );
  NAND U3423 ( .A(\stack[1][18] ), .B(n3148), .Z(n3112) );
  NAND U3424 ( .A(n3113), .B(n3112), .Z(\U1/RSOP_16/C3/Z_18 ) );
  NAND U3425 ( .A(n3151), .B(o[17]), .Z(n3115) );
  NAND U3426 ( .A(\stack[1][17] ), .B(n3148), .Z(n3114) );
  NAND U3427 ( .A(n3115), .B(n3114), .Z(\U1/RSOP_16/C3/Z_17 ) );
  NAND U3428 ( .A(n3151), .B(o[16]), .Z(n3117) );
  NAND U3429 ( .A(\stack[1][16] ), .B(n3148), .Z(n3116) );
  NAND U3430 ( .A(n3117), .B(n3116), .Z(\U1/RSOP_16/C3/Z_16 ) );
  NAND U3431 ( .A(n3151), .B(o[15]), .Z(n3119) );
  NAND U3432 ( .A(\stack[1][15] ), .B(n3148), .Z(n3118) );
  NAND U3433 ( .A(n3119), .B(n3118), .Z(\U1/RSOP_16/C3/Z_15 ) );
  NAND U3434 ( .A(n3151), .B(o[14]), .Z(n3121) );
  NAND U3435 ( .A(\stack[1][14] ), .B(n3148), .Z(n3120) );
  NAND U3436 ( .A(n3121), .B(n3120), .Z(\U1/RSOP_16/C3/Z_14 ) );
  NAND U3437 ( .A(n3151), .B(o[13]), .Z(n3123) );
  NAND U3438 ( .A(\stack[1][13] ), .B(n3148), .Z(n3122) );
  NAND U3439 ( .A(n3123), .B(n3122), .Z(\U1/RSOP_16/C3/Z_13 ) );
  NAND U3440 ( .A(n3151), .B(o[12]), .Z(n3125) );
  NAND U3441 ( .A(\stack[1][12] ), .B(n3148), .Z(n3124) );
  NAND U3442 ( .A(n3125), .B(n3124), .Z(\U1/RSOP_16/C3/Z_12 ) );
  NAND U3443 ( .A(n3151), .B(o[11]), .Z(n3127) );
  NAND U3444 ( .A(\stack[1][11] ), .B(n3148), .Z(n3126) );
  NAND U3445 ( .A(n3127), .B(n3126), .Z(\U1/RSOP_16/C3/Z_11 ) );
  NAND U3446 ( .A(n3151), .B(o[10]), .Z(n3129) );
  NAND U3447 ( .A(\stack[1][10] ), .B(n3148), .Z(n3128) );
  NAND U3448 ( .A(n3129), .B(n3128), .Z(\U1/RSOP_16/C3/Z_10 ) );
  NAND U3449 ( .A(n3151), .B(o[9]), .Z(n3131) );
  NAND U3450 ( .A(\stack[1][9] ), .B(n3148), .Z(n3130) );
  NAND U3451 ( .A(n3131), .B(n3130), .Z(\U1/RSOP_16/C3/Z_9 ) );
  NAND U3452 ( .A(n3151), .B(o[8]), .Z(n3133) );
  NAND U3453 ( .A(\stack[1][8] ), .B(n3148), .Z(n3132) );
  NAND U3454 ( .A(n3133), .B(n3132), .Z(\U1/RSOP_16/C3/Z_8 ) );
  NAND U3455 ( .A(n3151), .B(o[7]), .Z(n3135) );
  NAND U3456 ( .A(\stack[1][7] ), .B(n3148), .Z(n3134) );
  NAND U3457 ( .A(n3135), .B(n3134), .Z(\U1/RSOP_16/C3/Z_7 ) );
  NAND U3458 ( .A(n3151), .B(o[6]), .Z(n3137) );
  NAND U3459 ( .A(\stack[1][6] ), .B(n3148), .Z(n3136) );
  NAND U3460 ( .A(n3137), .B(n3136), .Z(\U1/RSOP_16/C3/Z_6 ) );
  NAND U3461 ( .A(n3151), .B(o[5]), .Z(n3139) );
  NAND U3462 ( .A(\stack[1][5] ), .B(n3148), .Z(n3138) );
  NAND U3463 ( .A(n3139), .B(n3138), .Z(\U1/RSOP_16/C3/Z_5 ) );
  NAND U3464 ( .A(n3151), .B(o[4]), .Z(n3141) );
  NAND U3465 ( .A(\stack[1][4] ), .B(n3148), .Z(n3140) );
  NAND U3466 ( .A(n3141), .B(n3140), .Z(\U1/RSOP_16/C3/Z_4 ) );
  NAND U3467 ( .A(n3151), .B(o[3]), .Z(n3143) );
  NAND U3468 ( .A(\stack[1][3] ), .B(n3148), .Z(n3142) );
  NAND U3469 ( .A(n3143), .B(n3142), .Z(\U1/RSOP_16/C3/Z_3 ) );
  NAND U3470 ( .A(n3151), .B(o[2]), .Z(n3145) );
  NAND U3471 ( .A(\stack[1][2] ), .B(n3148), .Z(n3144) );
  NAND U3472 ( .A(n3145), .B(n3144), .Z(\U1/RSOP_16/C3/Z_2 ) );
  NAND U3473 ( .A(n3151), .B(o[1]), .Z(n3147) );
  NAND U3474 ( .A(\stack[1][1] ), .B(n3148), .Z(n3146) );
  NAND U3475 ( .A(n3147), .B(n3146), .Z(\U1/RSOP_16/C3/Z_1 ) );
  NAND U3476 ( .A(n3151), .B(o[0]), .Z(n3150) );
  NAND U3477 ( .A(\stack[1][0] ), .B(n3148), .Z(n3149) );
  NAND U3478 ( .A(n3150), .B(n3149), .Z(\U1/RSOP_16/C3/Z_0 ) );
  NANDN U3479 ( .A(n3151), .B(n3152), .Z(\C1/Z_0 ) );
  NANDN U3480 ( .A(n3153), .B(n3152), .Z(n3217) );
  NAND U3481 ( .A(\C3/DATA5_63 ), .B(n3217), .Z(n3154) );
  AND U3482 ( .A(n15046), .B(n3154), .Z(n15050) );
  NAND U3483 ( .A(\C3/DATA5_36 ), .B(n3217), .Z(n3155) );
  AND U3484 ( .A(n16093), .B(n3155), .Z(n16094) );
  NAND U3485 ( .A(\C3/DATA5_34 ), .B(n3217), .Z(n3156) );
  AND U3486 ( .A(n16169), .B(n3156), .Z(n16170) );
  NAND U3487 ( .A(\C3/DATA5_32 ), .B(n3217), .Z(n3157) );
  AND U3488 ( .A(n16245), .B(n3157), .Z(n16246) );
  NAND U3489 ( .A(\C3/DATA5_31 ), .B(n3217), .Z(n3158) );
  AND U3490 ( .A(n16284), .B(n3158), .Z(n16285) );
  NAND U3491 ( .A(\C3/DATA5_30 ), .B(n3217), .Z(n3159) );
  AND U3492 ( .A(n16323), .B(n3159), .Z(n16324) );
  NAND U3493 ( .A(\C3/DATA5_28 ), .B(n3217), .Z(n3160) );
  AND U3494 ( .A(n16400), .B(n3160), .Z(n16401) );
  NAND U3495 ( .A(\C3/DATA5_27 ), .B(n3217), .Z(n3161) );
  NAND U3496 ( .A(n16436), .B(n3161), .Z(n16441) );
  NAND U3497 ( .A(\C3/DATA5_26 ), .B(n3217), .Z(n3162) );
  AND U3498 ( .A(n16478), .B(n3162), .Z(n16479) );
  NAND U3499 ( .A(\C3/DATA5_24 ), .B(n3217), .Z(n3163) );
  AND U3500 ( .A(n16556), .B(n3163), .Z(n16557) );
  NAND U3501 ( .A(\C3/DATA5_23 ), .B(n3217), .Z(n3164) );
  AND U3502 ( .A(n16595), .B(n3164), .Z(n16596) );
  NAND U3503 ( .A(\C3/DATA5_22 ), .B(n3217), .Z(n3165) );
  AND U3504 ( .A(n16634), .B(n3165), .Z(n16635) );
  NAND U3505 ( .A(\C3/DATA5_21 ), .B(n3217), .Z(n3166) );
  AND U3506 ( .A(n16673), .B(n3166), .Z(n16674) );
  NAND U3507 ( .A(\C3/DATA5_20 ), .B(n3217), .Z(n3167) );
  AND U3508 ( .A(n16713), .B(n3167), .Z(n16714) );
  NAND U3509 ( .A(\C3/DATA5_19 ), .B(n3217), .Z(n3168) );
  AND U3510 ( .A(n16753), .B(n3168), .Z(n16754) );
  NAND U3511 ( .A(\C3/DATA5_18 ), .B(n3217), .Z(n3169) );
  AND U3512 ( .A(n16793), .B(n3169), .Z(n16794) );
  NAND U3513 ( .A(\C3/DATA5_17 ), .B(n3217), .Z(n3170) );
  AND U3514 ( .A(n16833), .B(n3170), .Z(n16834) );
  NAND U3515 ( .A(\C3/DATA5_15 ), .B(n3217), .Z(n3171) );
  AND U3516 ( .A(n16911), .B(n3171), .Z(n16912) );
  NAND U3517 ( .A(\C3/DATA5_14 ), .B(n3217), .Z(n3172) );
  AND U3518 ( .A(n16950), .B(n3172), .Z(n16951) );
  NAND U3519 ( .A(\C3/DATA5_13 ), .B(n3217), .Z(n3173) );
  AND U3520 ( .A(n16989), .B(n3173), .Z(n16990) );
  NAND U3521 ( .A(\C3/DATA5_12 ), .B(n3217), .Z(n3174) );
  AND U3522 ( .A(n17028), .B(n3174), .Z(n17029) );
  NAND U3523 ( .A(\C3/DATA5_11 ), .B(n3217), .Z(n3175) );
  AND U3524 ( .A(n17067), .B(n3175), .Z(n17068) );
  NAND U3525 ( .A(\C3/DATA5_10 ), .B(n3217), .Z(n3176) );
  AND U3526 ( .A(n17106), .B(n3176), .Z(n17107) );
  NAND U3527 ( .A(\C3/DATA5_9 ), .B(n3217), .Z(n3177) );
  AND U3528 ( .A(n17146), .B(n3177), .Z(n17147) );
  NAND U3529 ( .A(\C3/DATA5_8 ), .B(n3217), .Z(n3178) );
  AND U3530 ( .A(n17186), .B(n3178), .Z(n17187) );
  NAND U3531 ( .A(\C3/DATA5_6 ), .B(n3217), .Z(n3179) );
  AND U3532 ( .A(n17259), .B(n3179), .Z(n17264) );
  NAND U3533 ( .A(\C3/DATA5_5 ), .B(n3217), .Z(n3180) );
  NAND U3534 ( .A(n17303), .B(n3180), .Z(n17304) );
  NAND U3535 ( .A(\C3/DATA5_4 ), .B(n3217), .Z(n3181) );
  AND U3536 ( .A(n17344), .B(n3181), .Z(n17345) );
  NAND U3537 ( .A(\C3/DATA5_3 ), .B(n3217), .Z(n3182) );
  AND U3538 ( .A(n17378), .B(n3182), .Z(n17383) );
  NAND U3539 ( .A(\C3/DATA5_2 ), .B(n3217), .Z(n3183) );
  NAND U3540 ( .A(n17421), .B(n3183), .Z(n17425) );
  NAND U3541 ( .A(\C3/DATA5_1 ), .B(n3217), .Z(n3184) );
  AND U3542 ( .A(n17468), .B(n3184), .Z(n17469) );
  NAND U3543 ( .A(\C3/DATA5_0 ), .B(n3217), .Z(n3185) );
  AND U3544 ( .A(n17487), .B(n3185), .Z(n17488) );
  NAND U3545 ( .A(\C3/DATA5_62 ), .B(n3217), .Z(n3186) );
  NAND U3546 ( .A(n15095), .B(n3186), .Z(n2142) );
  NAND U3547 ( .A(\C3/DATA5_61 ), .B(n3217), .Z(n3187) );
  NAND U3548 ( .A(n15133), .B(n3187), .Z(n2150) );
  NAND U3549 ( .A(\C3/DATA5_60 ), .B(n3217), .Z(n3188) );
  NAND U3550 ( .A(n15172), .B(n3188), .Z(n2158) );
  NAND U3551 ( .A(\C3/DATA5_59 ), .B(n3217), .Z(n3189) );
  NAND U3552 ( .A(n15211), .B(n3189), .Z(n2166) );
  NAND U3553 ( .A(\C3/DATA5_58 ), .B(n3217), .Z(n3190) );
  NAND U3554 ( .A(n15250), .B(n3190), .Z(n2174) );
  NAND U3555 ( .A(\C3/DATA5_57 ), .B(n3217), .Z(n3191) );
  NAND U3556 ( .A(n15288), .B(n3191), .Z(n2182) );
  NAND U3557 ( .A(\C3/DATA5_56 ), .B(n3217), .Z(n3192) );
  NAND U3558 ( .A(n15327), .B(n3192), .Z(n2190) );
  NAND U3559 ( .A(\C3/DATA5_55 ), .B(n3217), .Z(n3193) );
  NAND U3560 ( .A(n15365), .B(n3193), .Z(n2198) );
  NAND U3561 ( .A(\C3/DATA5_54 ), .B(n3217), .Z(n3194) );
  NAND U3562 ( .A(n15403), .B(n3194), .Z(n2206) );
  NAND U3563 ( .A(\C3/DATA5_53 ), .B(n3217), .Z(n3195) );
  NAND U3564 ( .A(n15441), .B(n3195), .Z(n2214) );
  NAND U3565 ( .A(\C3/DATA5_52 ), .B(n3217), .Z(n3196) );
  NAND U3566 ( .A(n15480), .B(n3196), .Z(n2222) );
  NAND U3567 ( .A(\C3/DATA5_51 ), .B(n3217), .Z(n3197) );
  NAND U3568 ( .A(n15519), .B(n3197), .Z(n2230) );
  NAND U3569 ( .A(\C3/DATA5_50 ), .B(n3217), .Z(n3198) );
  NAND U3570 ( .A(n15558), .B(n3198), .Z(n2238) );
  NAND U3571 ( .A(\C3/DATA5_49 ), .B(n3217), .Z(n3199) );
  NAND U3572 ( .A(n15596), .B(n3199), .Z(n2246) );
  NAND U3573 ( .A(\C3/DATA5_48 ), .B(n3217), .Z(n3200) );
  NAND U3574 ( .A(n15635), .B(n3200), .Z(n2254) );
  NAND U3575 ( .A(\C3/DATA5_47 ), .B(n3217), .Z(n3201) );
  NAND U3576 ( .A(n15674), .B(n3201), .Z(n2262) );
  NAND U3577 ( .A(\C3/DATA5_46 ), .B(n3217), .Z(n3202) );
  NAND U3578 ( .A(n15713), .B(n3202), .Z(n2270) );
  NAND U3579 ( .A(\C3/DATA5_45 ), .B(n3217), .Z(n3203) );
  NAND U3580 ( .A(n15752), .B(n3203), .Z(n2278) );
  NAND U3581 ( .A(\C3/DATA5_44 ), .B(n3217), .Z(n3204) );
  NAND U3582 ( .A(n15791), .B(n3204), .Z(n2286) );
  NAND U3583 ( .A(\C3/DATA5_43 ), .B(n3217), .Z(n3205) );
  NAND U3584 ( .A(n15830), .B(n3205), .Z(n2294) );
  NAND U3585 ( .A(\C3/DATA5_42 ), .B(n3217), .Z(n3206) );
  NAND U3586 ( .A(n15869), .B(n3206), .Z(n2302) );
  NAND U3587 ( .A(\C3/DATA5_41 ), .B(n3217), .Z(n3207) );
  NAND U3588 ( .A(n15908), .B(n3207), .Z(n2310) );
  NAND U3589 ( .A(\C3/DATA5_40 ), .B(n3217), .Z(n3208) );
  NAND U3590 ( .A(n15947), .B(n3208), .Z(n2318) );
  NAND U3591 ( .A(\C3/DATA5_39 ), .B(n3217), .Z(n3209) );
  NAND U3592 ( .A(n15985), .B(n3209), .Z(n2326) );
  NAND U3593 ( .A(\C3/DATA5_38 ), .B(n3217), .Z(n3210) );
  NAND U3594 ( .A(n16023), .B(n3210), .Z(n2334) );
  NAND U3595 ( .A(\C3/DATA5_37 ), .B(n3217), .Z(n3211) );
  NAND U3596 ( .A(n16061), .B(n3211), .Z(n2342) );
  NAND U3597 ( .A(\C3/DATA5_35 ), .B(n3217), .Z(n3212) );
  NAND U3598 ( .A(n16137), .B(n3212), .Z(n2358) );
  NAND U3599 ( .A(\C3/DATA5_33 ), .B(n3217), .Z(n3213) );
  NAND U3600 ( .A(n16213), .B(n3213), .Z(n2374) );
  NAND U3601 ( .A(\C3/DATA5_29 ), .B(n3217), .Z(n3214) );
  NAND U3602 ( .A(n16367), .B(n3214), .Z(n2406) );
  NAND U3603 ( .A(\C3/DATA5_25 ), .B(n3217), .Z(n3215) );
  NAND U3604 ( .A(n16523), .B(n3215), .Z(n2438) );
  NAND U3605 ( .A(\C3/DATA5_16 ), .B(n3217), .Z(n3216) );
  NAND U3606 ( .A(n16878), .B(n3216), .Z(n2510) );
  NAND U3607 ( .A(\C3/DATA5_7 ), .B(n3217), .Z(n3218) );
  NAND U3608 ( .A(n17231), .B(n3218), .Z(n2582) );
  ANDN U3609 ( .B(n3221), .A(opcode[1]), .Z(n3222) );
  AND U3610 ( .A(n3222), .B(opcode[2]), .Z(n17471) );
  NANDN U3611 ( .A(n2967), .B(\stack[6][0] ), .Z(n3224) );
  NANDN U3612 ( .A(n17471), .B(\stack[7][0] ), .Z(n3223) );
  NAND U3613 ( .A(n3224), .B(n3223), .Z(n2121) );
  NANDN U3614 ( .A(n2967), .B(\stack[5][0] ), .Z(n3226) );
  NOR U3615 ( .A(opcode[1]), .B(n3219), .Z(n17472) );
  NANDN U3616 ( .A(n17472), .B(\stack[7][0] ), .Z(n3225) );
  AND U3617 ( .A(n3226), .B(n3225), .Z(n3229) );
  XOR U3618 ( .A(n3220), .B(opcode[0]), .Z(n3227) );
  NANDN U3619 ( .A(opcode[1]), .B(n3227), .Z(n17475) );
  NANDN U3620 ( .A(n17475), .B(\stack[6][0] ), .Z(n3228) );
  NAND U3621 ( .A(n3229), .B(n3228), .Z(n2122) );
  NANDN U3622 ( .A(n2967), .B(\stack[4][0] ), .Z(n3231) );
  NANDN U3623 ( .A(n17472), .B(\stack[6][0] ), .Z(n3230) );
  AND U3624 ( .A(n3231), .B(n3230), .Z(n3233) );
  NANDN U3625 ( .A(n17475), .B(\stack[5][0] ), .Z(n3232) );
  NAND U3626 ( .A(n3233), .B(n3232), .Z(n2123) );
  NANDN U3627 ( .A(n2967), .B(\stack[3][0] ), .Z(n3235) );
  NANDN U3628 ( .A(n17472), .B(\stack[5][0] ), .Z(n3234) );
  AND U3629 ( .A(n3235), .B(n3234), .Z(n3237) );
  NANDN U3630 ( .A(n17475), .B(\stack[4][0] ), .Z(n3236) );
  NAND U3631 ( .A(n3237), .B(n3236), .Z(n2124) );
  NANDN U3632 ( .A(n2967), .B(\stack[2][0] ), .Z(n3239) );
  NANDN U3633 ( .A(n17472), .B(\stack[4][0] ), .Z(n3238) );
  AND U3634 ( .A(n3239), .B(n3238), .Z(n3241) );
  NANDN U3635 ( .A(n17475), .B(\stack[3][0] ), .Z(n3240) );
  NAND U3636 ( .A(n3241), .B(n3240), .Z(n2125) );
  NANDN U3637 ( .A(n2968), .B(n17471), .Z(n3243) );
  NANDN U3638 ( .A(n17472), .B(\stack[3][0] ), .Z(n3242) );
  AND U3639 ( .A(n3243), .B(n3242), .Z(n3245) );
  NANDN U3640 ( .A(n17475), .B(\stack[2][0] ), .Z(n3244) );
  NAND U3641 ( .A(n3245), .B(n3244), .Z(n2126) );
  NANDN U3642 ( .A(n2967), .B(\stack[6][63] ), .Z(n3247) );
  NANDN U3643 ( .A(n17471), .B(\stack[7][63] ), .Z(n3246) );
  NAND U3644 ( .A(n3247), .B(n3246), .Z(n2127) );
  NANDN U3645 ( .A(n2967), .B(\stack[5][63] ), .Z(n3249) );
  NANDN U3646 ( .A(n17472), .B(\stack[7][63] ), .Z(n3248) );
  AND U3647 ( .A(n3249), .B(n3248), .Z(n3251) );
  NANDN U3648 ( .A(n17475), .B(\stack[6][63] ), .Z(n3250) );
  NAND U3649 ( .A(n3251), .B(n3250), .Z(n2128) );
  NANDN U3650 ( .A(n2967), .B(\stack[4][63] ), .Z(n3253) );
  NANDN U3651 ( .A(n17472), .B(\stack[6][63] ), .Z(n3252) );
  AND U3652 ( .A(n3253), .B(n3252), .Z(n3255) );
  NANDN U3653 ( .A(n17475), .B(\stack[5][63] ), .Z(n3254) );
  NAND U3654 ( .A(n3255), .B(n3254), .Z(n2129) );
  NANDN U3655 ( .A(n2967), .B(\stack[3][63] ), .Z(n3257) );
  NANDN U3656 ( .A(n17472), .B(\stack[5][63] ), .Z(n3256) );
  AND U3657 ( .A(n3257), .B(n3256), .Z(n3259) );
  NANDN U3658 ( .A(n17475), .B(\stack[4][63] ), .Z(n3258) );
  NAND U3659 ( .A(n3259), .B(n3258), .Z(n2130) );
  NANDN U3660 ( .A(n2967), .B(\stack[2][63] ), .Z(n3261) );
  NANDN U3661 ( .A(n17472), .B(\stack[4][63] ), .Z(n3260) );
  AND U3662 ( .A(n3261), .B(n3260), .Z(n3263) );
  NANDN U3663 ( .A(n17475), .B(\stack[3][63] ), .Z(n3262) );
  NAND U3664 ( .A(n3263), .B(n3262), .Z(n2131) );
  NANDN U3665 ( .A(n2967), .B(\stack[1][63] ), .Z(n3265) );
  NANDN U3666 ( .A(n17472), .B(\stack[3][63] ), .Z(n3264) );
  AND U3667 ( .A(n3265), .B(n3264), .Z(n3267) );
  NANDN U3668 ( .A(n17475), .B(\stack[2][63] ), .Z(n3266) );
  NAND U3669 ( .A(n3267), .B(n3266), .Z(n2132) );
  NANDN U3670 ( .A(n2967), .B(o[63]), .Z(n3269) );
  NANDN U3671 ( .A(n17472), .B(\stack[2][63] ), .Z(n3268) );
  AND U3672 ( .A(n3269), .B(n3268), .Z(n3271) );
  NANDN U3673 ( .A(n17475), .B(\stack[1][63] ), .Z(n3270) );
  NAND U3674 ( .A(n3271), .B(n3270), .Z(n2133) );
  AND U3675 ( .A(o[61]), .B(\stack[1][0] ), .Z(n13715) );
  AND U3676 ( .A(o[59]), .B(\stack[1][0] ), .Z(n13021) );
  AND U3677 ( .A(o[57]), .B(\stack[1][0] ), .Z(n12351) );
  AND U3678 ( .A(o[55]), .B(\stack[1][0] ), .Z(n11706) );
  AND U3679 ( .A(o[53]), .B(\stack[1][0] ), .Z(n11084) );
  AND U3680 ( .A(o[51]), .B(\stack[1][0] ), .Z(n10487) );
  AND U3681 ( .A(o[49]), .B(\stack[1][0] ), .Z(n9914) );
  AND U3682 ( .A(o[47]), .B(\stack[1][0] ), .Z(n9365) );
  AND U3683 ( .A(o[45]), .B(\stack[1][0] ), .Z(n8839) );
  AND U3684 ( .A(o[43]), .B(\stack[1][0] ), .Z(n8337) );
  AND U3685 ( .A(o[41]), .B(\stack[1][0] ), .Z(n7858) );
  AND U3686 ( .A(o[39]), .B(\stack[1][0] ), .Z(n7404) );
  AND U3687 ( .A(o[37]), .B(\stack[1][0] ), .Z(n6972) );
  AND U3688 ( .A(o[35]), .B(\stack[1][0] ), .Z(n6563) );
  AND U3689 ( .A(o[33]), .B(\stack[1][0] ), .Z(n6177) );
  AND U3690 ( .A(o[31]), .B(\stack[1][0] ), .Z(n5816) );
  AND U3691 ( .A(o[29]), .B(\stack[1][0] ), .Z(n5640) );
  AND U3692 ( .A(o[27]), .B(\stack[1][0] ), .Z(n5314) );
  AND U3693 ( .A(o[25]), .B(\stack[1][0] ), .Z(n4876) );
  AND U3694 ( .A(o[23]), .B(\stack[1][0] ), .Z(n4611) );
  AND U3695 ( .A(o[21]), .B(\stack[1][0] ), .Z(n4483) );
  AND U3696 ( .A(o[19]), .B(\stack[1][0] ), .Z(n4152) );
  AND U3697 ( .A(o[17]), .B(\stack[1][0] ), .Z(n3959) );
  AND U3698 ( .A(o[15]), .B(\stack[1][0] ), .Z(n3789) );
  AND U3699 ( .A(o[13]), .B(\stack[1][0] ), .Z(n3643) );
  AND U3700 ( .A(o[11]), .B(\stack[1][0] ), .Z(n3522) );
  AND U3701 ( .A(o[9]), .B(\stack[1][0] ), .Z(n3425) );
  AND U3702 ( .A(o[7]), .B(\stack[1][0] ), .Z(n3352) );
  AND U3703 ( .A(o[5]), .B(\stack[1][0] ), .Z(n3303) );
  AND U3704 ( .A(o[3]), .B(\stack[1][0] ), .Z(n3280) );
  AND U3705 ( .A(\stack[1][1] ), .B(o[0]), .Z(n17456) );
  NANDN U3706 ( .A(n2995), .B(n17456), .Z(n3272) );
  XOR U3707 ( .A(n2996), .B(n3272), .Z(n3273) );
  NANDN U3708 ( .A(n2968), .B(n3273), .Z(n17417) );
  ANDN U3709 ( .B(o[0]), .A(n2970), .Z(n3275) );
  ANDN U3710 ( .B(o[1]), .A(n2969), .Z(n3274) );
  XOR U3711 ( .A(n3275), .B(n3274), .Z(n17418) );
  OR U3712 ( .A(n17417), .B(n17418), .Z(n3279) );
  NANDN U3713 ( .A(n2968), .B(o[1]), .Z(n17457) );
  NANDN U3714 ( .A(n17457), .B(n17456), .Z(n3277) );
  NANDN U3715 ( .A(n2968), .B(o[2]), .Z(n3276) );
  AND U3716 ( .A(n3277), .B(n3276), .Z(n3278) );
  ANDN U3717 ( .B(n3279), .A(n3278), .Z(n3281) );
  OR U3718 ( .A(n3280), .B(n3281), .Z(n3287) );
  XNOR U3719 ( .A(n3281), .B(n3280), .Z(n17380) );
  IV U3720 ( .A(\stack[1][3] ), .Z(n17375) );
  ANDN U3721 ( .B(o[0]), .A(n17375), .Z(n3283) );
  ANDN U3722 ( .B(o[1]), .A(n2970), .Z(n3282) );
  XOR U3723 ( .A(n3283), .B(n3282), .Z(n3288) );
  NANDN U3724 ( .A(n2995), .B(\stack[1][2] ), .Z(n3290) );
  OR U3725 ( .A(n3290), .B(n2994), .Z(n3284) );
  XOR U3726 ( .A(n2996), .B(n3284), .Z(n3285) );
  NANDN U3727 ( .A(n2969), .B(n3285), .Z(n3289) );
  XNOR U3728 ( .A(n3288), .B(n3289), .Z(n17379) );
  OR U3729 ( .A(n17380), .B(n17379), .Z(n3286) );
  AND U3730 ( .A(n3287), .B(n3286), .Z(n3300) );
  OR U3731 ( .A(n3289), .B(n3288), .Z(n3294) );
  NANDN U3732 ( .A(n3290), .B(n17456), .Z(n3292) );
  NANDN U3733 ( .A(n2996), .B(\stack[1][1] ), .Z(n3291) );
  AND U3734 ( .A(n3292), .B(n3291), .Z(n3293) );
  ANDN U3735 ( .B(n3294), .A(n3293), .Z(n3305) );
  AND U3736 ( .A(o[3]), .B(\stack[1][1] ), .Z(n3306) );
  XNOR U3737 ( .A(n3305), .B(n3306), .Z(n3308) );
  ANDN U3738 ( .B(o[0]), .A(n2971), .Z(n3296) );
  ANDN U3739 ( .B(o[1]), .A(n17375), .Z(n3295) );
  XOR U3740 ( .A(n3296), .B(n3295), .Z(n3314) );
  NANDN U3741 ( .A(n2995), .B(\stack[1][3] ), .Z(n3312) );
  OR U3742 ( .A(n3312), .B(n2994), .Z(n3297) );
  XOR U3743 ( .A(n2996), .B(n3297), .Z(n3298) );
  NANDN U3744 ( .A(n2970), .B(n3298), .Z(n3315) );
  XNOR U3745 ( .A(n3314), .B(n3315), .Z(n3307) );
  XOR U3746 ( .A(n3308), .B(n3307), .Z(n3299) );
  NANDN U3747 ( .A(n3300), .B(n3299), .Z(n3302) );
  XOR U3748 ( .A(n3300), .B(n3299), .Z(n17341) );
  AND U3749 ( .A(o[4]), .B(\stack[1][0] ), .Z(n17342) );
  OR U3750 ( .A(n17341), .B(n17342), .Z(n3301) );
  AND U3751 ( .A(n3302), .B(n3301), .Z(n3304) );
  OR U3752 ( .A(n3303), .B(n3304), .Z(n3323) );
  XNOR U3753 ( .A(n3304), .B(n3303), .Z(n17299) );
  OR U3754 ( .A(n3306), .B(n3305), .Z(n3310) );
  OR U3755 ( .A(n3308), .B(n3307), .Z(n3309) );
  NAND U3756 ( .A(n3310), .B(n3309), .Z(n3343) );
  ANDN U3757 ( .B(\stack[1][2] ), .A(n2994), .Z(n3311) );
  NANDN U3758 ( .A(n3312), .B(n3311), .Z(n3313) );
  NANDN U3759 ( .A(n2970), .B(o[2]), .Z(n17420) );
  NAND U3760 ( .A(n3313), .B(n17420), .Z(n3317) );
  OR U3761 ( .A(n3315), .B(n3314), .Z(n3316) );
  AND U3762 ( .A(n3317), .B(n3316), .Z(n3324) );
  AND U3763 ( .A(o[3]), .B(\stack[1][2] ), .Z(n3325) );
  XNOR U3764 ( .A(n3324), .B(n3325), .Z(n3327) );
  IV U3765 ( .A(\stack[1][5] ), .Z(n17296) );
  ANDN U3766 ( .B(o[0]), .A(n17296), .Z(n3319) );
  ANDN U3767 ( .B(o[1]), .A(n2971), .Z(n3318) );
  XOR U3768 ( .A(n3319), .B(n3318), .Z(n3330) );
  NANDN U3769 ( .A(n2995), .B(\stack[1][4] ), .Z(n3333) );
  OR U3770 ( .A(n3333), .B(n2994), .Z(n3320) );
  XOR U3771 ( .A(n2996), .B(n3320), .Z(n3321) );
  NANDN U3772 ( .A(n17375), .B(n3321), .Z(n3331) );
  XNOR U3773 ( .A(n3330), .B(n3331), .Z(n3326) );
  XOR U3774 ( .A(n3327), .B(n3326), .Z(n3342) );
  XOR U3775 ( .A(n3343), .B(n3342), .Z(n3344) );
  NANDN U3776 ( .A(n2969), .B(o[4]), .Z(n3345) );
  XNOR U3777 ( .A(n3344), .B(n3345), .Z(n17300) );
  OR U3778 ( .A(n17299), .B(n17300), .Z(n3322) );
  AND U3779 ( .A(n3323), .B(n3322), .Z(n3349) );
  NANDN U3780 ( .A(n2970), .B(o[4]), .Z(n3380) );
  OR U3781 ( .A(n3325), .B(n3324), .Z(n3329) );
  OR U3782 ( .A(n3327), .B(n3326), .Z(n3328) );
  NAND U3783 ( .A(n3329), .B(n3328), .Z(n3378) );
  AND U3784 ( .A(\stack[1][3] ), .B(o[3]), .Z(n17384) );
  OR U3785 ( .A(n3331), .B(n3330), .Z(n3337) );
  ANDN U3786 ( .B(\stack[1][3] ), .A(n2994), .Z(n3332) );
  NANDN U3787 ( .A(n3333), .B(n3332), .Z(n3335) );
  NANDN U3788 ( .A(n17375), .B(o[2]), .Z(n3334) );
  AND U3789 ( .A(n3335), .B(n3334), .Z(n3336) );
  ANDN U3790 ( .B(n3337), .A(n3336), .Z(n3360) );
  XNOR U3791 ( .A(n17384), .B(n3360), .Z(n3362) );
  IV U3792 ( .A(\stack[1][6] ), .Z(n17256) );
  ANDN U3793 ( .B(o[0]), .A(n17256), .Z(n3339) );
  ANDN U3794 ( .B(o[1]), .A(n17296), .Z(n3338) );
  XOR U3795 ( .A(n3339), .B(n3338), .Z(n3365) );
  NANDN U3796 ( .A(n2995), .B(\stack[1][5] ), .Z(n3368) );
  OR U3797 ( .A(n3368), .B(n2994), .Z(n3340) );
  XOR U3798 ( .A(n2996), .B(n3340), .Z(n3341) );
  NANDN U3799 ( .A(n2971), .B(n3341), .Z(n3366) );
  XNOR U3800 ( .A(n3365), .B(n3366), .Z(n3361) );
  XOR U3801 ( .A(n3362), .B(n3361), .Z(n3377) );
  XNOR U3802 ( .A(n3378), .B(n3377), .Z(n3379) );
  AND U3803 ( .A(o[5]), .B(\stack[1][1] ), .Z(n3354) );
  OR U3804 ( .A(n3343), .B(n3342), .Z(n3347) );
  NANDN U3805 ( .A(n3345), .B(n3344), .Z(n3346) );
  NAND U3806 ( .A(n3347), .B(n3346), .Z(n3355) );
  XNOR U3807 ( .A(n3354), .B(n3355), .Z(n3357) );
  XOR U3808 ( .A(n3356), .B(n3357), .Z(n3348) );
  NANDN U3809 ( .A(n3349), .B(n3348), .Z(n3351) );
  XOR U3810 ( .A(n3349), .B(n3348), .Z(n17260) );
  AND U3811 ( .A(o[6]), .B(\stack[1][0] ), .Z(n17261) );
  OR U3812 ( .A(n17260), .B(n17261), .Z(n3350) );
  AND U3813 ( .A(n3351), .B(n3350), .Z(n3353) );
  OR U3814 ( .A(n3352), .B(n3353), .Z(n3384) );
  XNOR U3815 ( .A(n3353), .B(n3352), .Z(n17222) );
  NANDN U3816 ( .A(n2969), .B(o[6]), .Z(n3388) );
  OR U3817 ( .A(n3355), .B(n3354), .Z(n3359) );
  OR U3818 ( .A(n3357), .B(n3356), .Z(n3358) );
  NAND U3819 ( .A(n3359), .B(n3358), .Z(n3386) );
  OR U3820 ( .A(n3360), .B(n17384), .Z(n3364) );
  OR U3821 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U3822 ( .A(n3364), .B(n3363), .Z(n3416) );
  OR U3823 ( .A(n3366), .B(n3365), .Z(n3372) );
  ANDN U3824 ( .B(\stack[1][4] ), .A(n2994), .Z(n3367) );
  NANDN U3825 ( .A(n3368), .B(n3367), .Z(n3370) );
  NANDN U3826 ( .A(n2971), .B(o[2]), .Z(n3369) );
  AND U3827 ( .A(n3370), .B(n3369), .Z(n3371) );
  ANDN U3828 ( .B(n3372), .A(n3371), .Z(n3397) );
  AND U3829 ( .A(\stack[1][4] ), .B(o[3]), .Z(n3398) );
  XNOR U3830 ( .A(n3397), .B(n3398), .Z(n3400) );
  IV U3831 ( .A(\stack[1][7] ), .Z(n17219) );
  ANDN U3832 ( .B(o[0]), .A(n17219), .Z(n3374) );
  ANDN U3833 ( .B(o[1]), .A(n17256), .Z(n3373) );
  XOR U3834 ( .A(n3374), .B(n3373), .Z(n3403) );
  NANDN U3835 ( .A(n2995), .B(\stack[1][6] ), .Z(n3406) );
  OR U3836 ( .A(n3406), .B(n2994), .Z(n3375) );
  XOR U3837 ( .A(n2996), .B(n3375), .Z(n3376) );
  NANDN U3838 ( .A(n17296), .B(n3376), .Z(n3404) );
  XNOR U3839 ( .A(n3403), .B(n3404), .Z(n3399) );
  XOR U3840 ( .A(n3400), .B(n3399), .Z(n3415) );
  XNOR U3841 ( .A(n3416), .B(n3415), .Z(n3417) );
  NANDN U3842 ( .A(n17375), .B(o[4]), .Z(n3418) );
  AND U3843 ( .A(o[5]), .B(\stack[1][2] ), .Z(n3391) );
  OR U3844 ( .A(n3378), .B(n3377), .Z(n3382) );
  OR U3845 ( .A(n3380), .B(n3379), .Z(n3381) );
  NAND U3846 ( .A(n3382), .B(n3381), .Z(n3392) );
  XOR U3847 ( .A(n3391), .B(n3392), .Z(n3393) );
  XNOR U3848 ( .A(n3394), .B(n3393), .Z(n3385) );
  XNOR U3849 ( .A(n3386), .B(n3385), .Z(n3387) );
  XOR U3850 ( .A(n3388), .B(n3387), .Z(n17223) );
  OR U3851 ( .A(n17222), .B(n17223), .Z(n3383) );
  AND U3852 ( .A(n3384), .B(n3383), .Z(n3422) );
  AND U3853 ( .A(o[7]), .B(\stack[1][1] ), .Z(n3427) );
  OR U3854 ( .A(n3386), .B(n3385), .Z(n3390) );
  OR U3855 ( .A(n3388), .B(n3387), .Z(n3389) );
  NAND U3856 ( .A(n3390), .B(n3389), .Z(n3428) );
  XNOR U3857 ( .A(n3427), .B(n3428), .Z(n3430) );
  OR U3858 ( .A(n3392), .B(n3391), .Z(n3396) );
  NANDN U3859 ( .A(n3394), .B(n3393), .Z(n3395) );
  AND U3860 ( .A(n3396), .B(n3395), .Z(n3434) );
  AND U3861 ( .A(o[4]), .B(\stack[1][4] ), .Z(n17338) );
  OR U3862 ( .A(n3398), .B(n3397), .Z(n3402) );
  OR U3863 ( .A(n3400), .B(n3399), .Z(n3401) );
  NAND U3864 ( .A(n3402), .B(n3401), .Z(n3464) );
  OR U3865 ( .A(n3404), .B(n3403), .Z(n3410) );
  ANDN U3866 ( .B(\stack[1][5] ), .A(n2994), .Z(n3405) );
  NANDN U3867 ( .A(n3406), .B(n3405), .Z(n3408) );
  NANDN U3868 ( .A(n17296), .B(o[2]), .Z(n3407) );
  AND U3869 ( .A(n3408), .B(n3407), .Z(n3409) );
  ANDN U3870 ( .B(n3410), .A(n3409), .Z(n3445) );
  AND U3871 ( .A(\stack[1][5] ), .B(o[3]), .Z(n3446) );
  XNOR U3872 ( .A(n3445), .B(n3446), .Z(n3448) );
  IV U3873 ( .A(\stack[1][8] ), .Z(n17179) );
  ANDN U3874 ( .B(o[0]), .A(n17179), .Z(n3412) );
  ANDN U3875 ( .B(o[1]), .A(n17219), .Z(n3411) );
  XOR U3876 ( .A(n3412), .B(n3411), .Z(n3451) );
  NANDN U3877 ( .A(n2995), .B(\stack[1][7] ), .Z(n3454) );
  OR U3878 ( .A(n3454), .B(n2994), .Z(n3413) );
  XOR U3879 ( .A(n2996), .B(n3413), .Z(n3414) );
  NANDN U3880 ( .A(n17256), .B(n3414), .Z(n3452) );
  XNOR U3881 ( .A(n3451), .B(n3452), .Z(n3447) );
  XOR U3882 ( .A(n3448), .B(n3447), .Z(n3463) );
  XNOR U3883 ( .A(n3464), .B(n3463), .Z(n3465) );
  AND U3884 ( .A(o[5]), .B(\stack[1][3] ), .Z(n3439) );
  OR U3885 ( .A(n3416), .B(n3415), .Z(n3420) );
  OR U3886 ( .A(n3418), .B(n3417), .Z(n3419) );
  NAND U3887 ( .A(n3420), .B(n3419), .Z(n3440) );
  XNOR U3888 ( .A(n3439), .B(n3440), .Z(n3442) );
  XOR U3889 ( .A(n3441), .B(n3442), .Z(n3433) );
  XOR U3890 ( .A(n3434), .B(n3433), .Z(n3436) );
  AND U3891 ( .A(o[6]), .B(\stack[1][2] ), .Z(n3435) );
  XNOR U3892 ( .A(n3436), .B(n3435), .Z(n3429) );
  NANDN U3893 ( .A(n3422), .B(n3421), .Z(n3424) );
  XOR U3894 ( .A(n3422), .B(n3421), .Z(n17183) );
  AND U3895 ( .A(o[8]), .B(\stack[1][0] ), .Z(n17184) );
  OR U3896 ( .A(n17183), .B(n17184), .Z(n3423) );
  AND U3897 ( .A(n3424), .B(n3423), .Z(n3426) );
  OR U3898 ( .A(n3425), .B(n3426), .Z(n3469) );
  XNOR U3899 ( .A(n3426), .B(n3425), .Z(n17142) );
  NANDN U3900 ( .A(n2969), .B(o[8]), .Z(n3515) );
  OR U3901 ( .A(n3428), .B(n3427), .Z(n3432) );
  OR U3902 ( .A(n3430), .B(n3429), .Z(n3431) );
  NAND U3903 ( .A(n3432), .B(n3431), .Z(n3513) );
  NANDN U3904 ( .A(n3434), .B(n3433), .Z(n3438) );
  OR U3905 ( .A(n3436), .B(n3435), .Z(n3437) );
  AND U3906 ( .A(n3438), .B(n3437), .Z(n3470) );
  AND U3907 ( .A(o[7]), .B(\stack[1][2] ), .Z(n3471) );
  XNOR U3908 ( .A(n3470), .B(n3471), .Z(n3473) );
  OR U3909 ( .A(n3440), .B(n3439), .Z(n3444) );
  OR U3910 ( .A(n3442), .B(n3441), .Z(n3443) );
  AND U3911 ( .A(n3444), .B(n3443), .Z(n3477) );
  OR U3912 ( .A(n3446), .B(n3445), .Z(n3450) );
  OR U3913 ( .A(n3448), .B(n3447), .Z(n3449) );
  NAND U3914 ( .A(n3450), .B(n3449), .Z(n3507) );
  OR U3915 ( .A(n3452), .B(n3451), .Z(n3458) );
  ANDN U3916 ( .B(\stack[1][6] ), .A(n2994), .Z(n3453) );
  NANDN U3917 ( .A(n3454), .B(n3453), .Z(n3456) );
  NANDN U3918 ( .A(n17256), .B(o[2]), .Z(n3455) );
  AND U3919 ( .A(n3456), .B(n3455), .Z(n3457) );
  ANDN U3920 ( .B(n3458), .A(n3457), .Z(n3488) );
  AND U3921 ( .A(\stack[1][6] ), .B(o[3]), .Z(n3489) );
  XNOR U3922 ( .A(n3488), .B(n3489), .Z(n3491) );
  IV U3923 ( .A(\stack[1][9] ), .Z(n17145) );
  ANDN U3924 ( .B(o[0]), .A(n17145), .Z(n3460) );
  ANDN U3925 ( .B(o[1]), .A(n17179), .Z(n3459) );
  XOR U3926 ( .A(n3460), .B(n3459), .Z(n3494) );
  NANDN U3927 ( .A(n2995), .B(\stack[1][8] ), .Z(n3497) );
  OR U3928 ( .A(n3497), .B(n2994), .Z(n3461) );
  XOR U3929 ( .A(n2996), .B(n3461), .Z(n3462) );
  NANDN U3930 ( .A(n17219), .B(n3462), .Z(n3495) );
  XNOR U3931 ( .A(n3494), .B(n3495), .Z(n3490) );
  XOR U3932 ( .A(n3491), .B(n3490), .Z(n3506) );
  XNOR U3933 ( .A(n3507), .B(n3506), .Z(n3508) );
  NANDN U3934 ( .A(n2998), .B(\stack[1][5] ), .Z(n3509) );
  AND U3935 ( .A(o[5]), .B(\stack[1][4] ), .Z(n3482) );
  OR U3936 ( .A(n3464), .B(n3463), .Z(n3467) );
  NANDN U3937 ( .A(n3465), .B(n17338), .Z(n3466) );
  NAND U3938 ( .A(n3467), .B(n3466), .Z(n3483) );
  XNOR U3939 ( .A(n3482), .B(n3483), .Z(n3485) );
  XOR U3940 ( .A(n3484), .B(n3485), .Z(n3476) );
  XOR U3941 ( .A(n3477), .B(n3476), .Z(n3479) );
  AND U3942 ( .A(o[6]), .B(\stack[1][3] ), .Z(n3478) );
  XNOR U3943 ( .A(n3479), .B(n3478), .Z(n3472) );
  XOR U3944 ( .A(n3473), .B(n3472), .Z(n3512) );
  XOR U3945 ( .A(n3513), .B(n3512), .Z(n3514) );
  XNOR U3946 ( .A(n3515), .B(n3514), .Z(n17143) );
  OR U3947 ( .A(n17142), .B(n17143), .Z(n3468) );
  AND U3948 ( .A(n3469), .B(n3468), .Z(n3519) );
  NANDN U3949 ( .A(n2970), .B(o[8]), .Z(n3574) );
  OR U3950 ( .A(n3471), .B(n3470), .Z(n3475) );
  OR U3951 ( .A(n3473), .B(n3472), .Z(n3474) );
  NAND U3952 ( .A(n3475), .B(n3474), .Z(n3572) );
  NANDN U3953 ( .A(n3477), .B(n3476), .Z(n3481) );
  OR U3954 ( .A(n3479), .B(n3478), .Z(n3480) );
  AND U3955 ( .A(n3481), .B(n3480), .Z(n3530) );
  AND U3956 ( .A(o[7]), .B(\stack[1][3] ), .Z(n3531) );
  XNOR U3957 ( .A(n3530), .B(n3531), .Z(n3533) );
  OR U3958 ( .A(n3483), .B(n3482), .Z(n3487) );
  OR U3959 ( .A(n3485), .B(n3484), .Z(n3486) );
  AND U3960 ( .A(n3487), .B(n3486), .Z(n3537) );
  OR U3961 ( .A(n3489), .B(n3488), .Z(n3493) );
  OR U3962 ( .A(n3491), .B(n3490), .Z(n3492) );
  NAND U3963 ( .A(n3493), .B(n3492), .Z(n3566) );
  OR U3964 ( .A(n3495), .B(n3494), .Z(n3501) );
  ANDN U3965 ( .B(\stack[1][7] ), .A(n2994), .Z(n3496) );
  NANDN U3966 ( .A(n3497), .B(n3496), .Z(n3499) );
  NANDN U3967 ( .A(n17219), .B(o[2]), .Z(n3498) );
  AND U3968 ( .A(n3499), .B(n3498), .Z(n3500) );
  ANDN U3969 ( .B(n3501), .A(n3500), .Z(n3547) );
  AND U3970 ( .A(\stack[1][7] ), .B(o[3]), .Z(n3548) );
  XNOR U3971 ( .A(n3547), .B(n3548), .Z(n3550) );
  IV U3972 ( .A(\stack[1][10] ), .Z(n17101) );
  ANDN U3973 ( .B(o[0]), .A(n17101), .Z(n3503) );
  ANDN U3974 ( .B(o[1]), .A(n17145), .Z(n3502) );
  XOR U3975 ( .A(n3503), .B(n3502), .Z(n3553) );
  NANDN U3976 ( .A(n2995), .B(\stack[1][9] ), .Z(n3556) );
  OR U3977 ( .A(n3556), .B(n2994), .Z(n3504) );
  XOR U3978 ( .A(n2996), .B(n3504), .Z(n3505) );
  NANDN U3979 ( .A(n17179), .B(n3505), .Z(n3554) );
  XNOR U3980 ( .A(n3553), .B(n3554), .Z(n3549) );
  XOR U3981 ( .A(n3550), .B(n3549), .Z(n3565) );
  XNOR U3982 ( .A(n3566), .B(n3565), .Z(n3567) );
  NANDN U3983 ( .A(n2998), .B(\stack[1][6] ), .Z(n3568) );
  AND U3984 ( .A(\stack[1][5] ), .B(o[5]), .Z(n17302) );
  OR U3985 ( .A(n3507), .B(n3506), .Z(n3511) );
  OR U3986 ( .A(n3509), .B(n3508), .Z(n3510) );
  NAND U3987 ( .A(n3511), .B(n3510), .Z(n3542) );
  XNOR U3988 ( .A(n17302), .B(n3542), .Z(n3544) );
  XOR U3989 ( .A(n3543), .B(n3544), .Z(n3536) );
  XOR U3990 ( .A(n3537), .B(n3536), .Z(n3539) );
  AND U3991 ( .A(o[6]), .B(\stack[1][4] ), .Z(n3538) );
  XNOR U3992 ( .A(n3539), .B(n3538), .Z(n3532) );
  XOR U3993 ( .A(n3533), .B(n3532), .Z(n3571) );
  XNOR U3994 ( .A(n3572), .B(n3571), .Z(n3573) );
  AND U3995 ( .A(o[9]), .B(\stack[1][1] ), .Z(n3524) );
  OR U3996 ( .A(n3513), .B(n3512), .Z(n3517) );
  NANDN U3997 ( .A(n3515), .B(n3514), .Z(n3516) );
  NAND U3998 ( .A(n3517), .B(n3516), .Z(n3525) );
  XNOR U3999 ( .A(n3524), .B(n3525), .Z(n3527) );
  XOR U4000 ( .A(n3526), .B(n3527), .Z(n3518) );
  NANDN U4001 ( .A(n3519), .B(n3518), .Z(n3521) );
  XOR U4002 ( .A(n3519), .B(n3518), .Z(n17103) );
  AND U4003 ( .A(o[10]), .B(\stack[1][0] ), .Z(n17104) );
  OR U4004 ( .A(n17103), .B(n17104), .Z(n3520) );
  AND U4005 ( .A(n3521), .B(n3520), .Z(n3523) );
  OR U4006 ( .A(n3522), .B(n3523), .Z(n3578) );
  XNOR U4007 ( .A(n3523), .B(n3522), .Z(n17064) );
  NANDN U4008 ( .A(n2969), .B(o[10]), .Z(n3636) );
  OR U4009 ( .A(n3525), .B(n3524), .Z(n3529) );
  OR U4010 ( .A(n3527), .B(n3526), .Z(n3528) );
  NAND U4011 ( .A(n3529), .B(n3528), .Z(n3634) );
  NANDN U4012 ( .A(n17375), .B(o[8]), .Z(n3630) );
  OR U4013 ( .A(n3531), .B(n3530), .Z(n3535) );
  OR U4014 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U4015 ( .A(n3535), .B(n3534), .Z(n3628) );
  NANDN U4016 ( .A(n3537), .B(n3536), .Z(n3541) );
  OR U4017 ( .A(n3539), .B(n3538), .Z(n3540) );
  AND U4018 ( .A(n3541), .B(n3540), .Z(n3585) );
  AND U4019 ( .A(o[7]), .B(\stack[1][4] ), .Z(n3586) );
  XNOR U4020 ( .A(n3585), .B(n3586), .Z(n3588) );
  OR U4021 ( .A(n3542), .B(n17302), .Z(n3546) );
  OR U4022 ( .A(n3544), .B(n3543), .Z(n3545) );
  AND U4023 ( .A(n3546), .B(n3545), .Z(n3592) );
  OR U4024 ( .A(n3548), .B(n3547), .Z(n3552) );
  OR U4025 ( .A(n3550), .B(n3549), .Z(n3551) );
  NAND U4026 ( .A(n3552), .B(n3551), .Z(n3622) );
  OR U4027 ( .A(n3554), .B(n3553), .Z(n3560) );
  ANDN U4028 ( .B(\stack[1][8] ), .A(n2994), .Z(n3555) );
  NANDN U4029 ( .A(n3556), .B(n3555), .Z(n3558) );
  NANDN U4030 ( .A(n17179), .B(o[2]), .Z(n3557) );
  AND U4031 ( .A(n3558), .B(n3557), .Z(n3559) );
  ANDN U4032 ( .B(n3560), .A(n3559), .Z(n3603) );
  AND U4033 ( .A(\stack[1][8] ), .B(o[3]), .Z(n3604) );
  XNOR U4034 ( .A(n3603), .B(n3604), .Z(n3606) );
  ANDN U4035 ( .B(o[0]), .A(n2972), .Z(n3562) );
  ANDN U4036 ( .B(o[1]), .A(n17101), .Z(n3561) );
  XOR U4037 ( .A(n3562), .B(n3561), .Z(n3609) );
  NANDN U4038 ( .A(n2995), .B(\stack[1][10] ), .Z(n3612) );
  OR U4039 ( .A(n3612), .B(n2994), .Z(n3563) );
  XOR U4040 ( .A(n2996), .B(n3563), .Z(n3564) );
  NANDN U4041 ( .A(n17145), .B(n3564), .Z(n3610) );
  XNOR U4042 ( .A(n3609), .B(n3610), .Z(n3605) );
  XOR U4043 ( .A(n3606), .B(n3605), .Z(n3621) );
  XNOR U4044 ( .A(n3622), .B(n3621), .Z(n3623) );
  NANDN U4045 ( .A(n2998), .B(\stack[1][7] ), .Z(n3624) );
  AND U4046 ( .A(\stack[1][6] ), .B(o[5]), .Z(n3597) );
  OR U4047 ( .A(n3566), .B(n3565), .Z(n3570) );
  OR U4048 ( .A(n3568), .B(n3567), .Z(n3569) );
  NAND U4049 ( .A(n3570), .B(n3569), .Z(n3598) );
  XNOR U4050 ( .A(n3597), .B(n3598), .Z(n3600) );
  XOR U4051 ( .A(n3599), .B(n3600), .Z(n3591) );
  XOR U4052 ( .A(n3592), .B(n3591), .Z(n3594) );
  AND U4053 ( .A(o[6]), .B(\stack[1][5] ), .Z(n3593) );
  XNOR U4054 ( .A(n3594), .B(n3593), .Z(n3587) );
  XOR U4055 ( .A(n3588), .B(n3587), .Z(n3627) );
  XNOR U4056 ( .A(n3628), .B(n3627), .Z(n3629) );
  AND U4057 ( .A(o[9]), .B(\stack[1][2] ), .Z(n3579) );
  OR U4058 ( .A(n3572), .B(n3571), .Z(n3576) );
  OR U4059 ( .A(n3574), .B(n3573), .Z(n3575) );
  NAND U4060 ( .A(n3576), .B(n3575), .Z(n3580) );
  XOR U4061 ( .A(n3579), .B(n3580), .Z(n3581) );
  XNOR U4062 ( .A(n3582), .B(n3581), .Z(n3633) );
  XNOR U4063 ( .A(n3634), .B(n3633), .Z(n3635) );
  XOR U4064 ( .A(n3636), .B(n3635), .Z(n17065) );
  OR U4065 ( .A(n17064), .B(n17065), .Z(n3577) );
  AND U4066 ( .A(n3578), .B(n3577), .Z(n3640) );
  NANDN U4067 ( .A(n2970), .B(o[10]), .Z(n3707) );
  OR U4068 ( .A(n3580), .B(n3579), .Z(n3584) );
  NANDN U4069 ( .A(n3582), .B(n3581), .Z(n3583) );
  NAND U4070 ( .A(n3584), .B(n3583), .Z(n3705) );
  NANDN U4071 ( .A(n2971), .B(o[8]), .Z(n3701) );
  OR U4072 ( .A(n3586), .B(n3585), .Z(n3590) );
  OR U4073 ( .A(n3588), .B(n3587), .Z(n3589) );
  NAND U4074 ( .A(n3590), .B(n3589), .Z(n3699) );
  NANDN U4075 ( .A(n3592), .B(n3591), .Z(n3596) );
  OR U4076 ( .A(n3594), .B(n3593), .Z(n3595) );
  AND U4077 ( .A(n3596), .B(n3595), .Z(n3657) );
  AND U4078 ( .A(o[7]), .B(\stack[1][5] ), .Z(n3658) );
  XNOR U4079 ( .A(n3657), .B(n3658), .Z(n3660) );
  AND U4080 ( .A(o[6]), .B(\stack[1][6] ), .Z(n17265) );
  OR U4081 ( .A(n3598), .B(n3597), .Z(n3602) );
  OR U4082 ( .A(n3600), .B(n3599), .Z(n3601) );
  AND U4083 ( .A(n3602), .B(n3601), .Z(n3664) );
  OR U4084 ( .A(n3604), .B(n3603), .Z(n3608) );
  OR U4085 ( .A(n3606), .B(n3605), .Z(n3607) );
  NAND U4086 ( .A(n3608), .B(n3607), .Z(n3693) );
  OR U4087 ( .A(n3610), .B(n3609), .Z(n3616) );
  ANDN U4088 ( .B(\stack[1][9] ), .A(n2994), .Z(n3611) );
  NANDN U4089 ( .A(n3612), .B(n3611), .Z(n3614) );
  NANDN U4090 ( .A(n17145), .B(o[2]), .Z(n3613) );
  AND U4091 ( .A(n3614), .B(n3613), .Z(n3615) );
  ANDN U4092 ( .B(n3616), .A(n3615), .Z(n3674) );
  AND U4093 ( .A(\stack[1][9] ), .B(o[3]), .Z(n3675) );
  XNOR U4094 ( .A(n3674), .B(n3675), .Z(n3677) );
  ANDN U4095 ( .B(o[0]), .A(n2973), .Z(n3618) );
  ANDN U4096 ( .B(o[1]), .A(n2972), .Z(n3617) );
  XOR U4097 ( .A(n3618), .B(n3617), .Z(n3680) );
  NANDN U4098 ( .A(n2995), .B(\stack[1][11] ), .Z(n3683) );
  OR U4099 ( .A(n3683), .B(n2994), .Z(n3619) );
  XOR U4100 ( .A(n2996), .B(n3619), .Z(n3620) );
  NANDN U4101 ( .A(n17101), .B(n3620), .Z(n3681) );
  XNOR U4102 ( .A(n3680), .B(n3681), .Z(n3676) );
  XOR U4103 ( .A(n3677), .B(n3676), .Z(n3692) );
  XNOR U4104 ( .A(n3693), .B(n3692), .Z(n3694) );
  NANDN U4105 ( .A(n2998), .B(\stack[1][8] ), .Z(n3695) );
  AND U4106 ( .A(\stack[1][7] ), .B(o[5]), .Z(n3668) );
  OR U4107 ( .A(n3622), .B(n3621), .Z(n3626) );
  OR U4108 ( .A(n3624), .B(n3623), .Z(n3625) );
  NAND U4109 ( .A(n3626), .B(n3625), .Z(n3669) );
  XNOR U4110 ( .A(n3668), .B(n3669), .Z(n3671) );
  XOR U4111 ( .A(n3670), .B(n3671), .Z(n3663) );
  XOR U4112 ( .A(n3664), .B(n3663), .Z(n3665) );
  XNOR U4113 ( .A(n17265), .B(n3665), .Z(n3659) );
  XOR U4114 ( .A(n3660), .B(n3659), .Z(n3698) );
  XNOR U4115 ( .A(n3699), .B(n3698), .Z(n3700) );
  AND U4116 ( .A(o[9]), .B(\stack[1][3] ), .Z(n3651) );
  OR U4117 ( .A(n3628), .B(n3627), .Z(n3632) );
  OR U4118 ( .A(n3630), .B(n3629), .Z(n3631) );
  NAND U4119 ( .A(n3632), .B(n3631), .Z(n3652) );
  XOR U4120 ( .A(n3651), .B(n3652), .Z(n3653) );
  XNOR U4121 ( .A(n3654), .B(n3653), .Z(n3704) );
  XNOR U4122 ( .A(n3705), .B(n3704), .Z(n3706) );
  XOR U4123 ( .A(n3707), .B(n3706), .Z(n3647) );
  AND U4124 ( .A(o[11]), .B(\stack[1][1] ), .Z(n3645) );
  OR U4125 ( .A(n3634), .B(n3633), .Z(n3638) );
  OR U4126 ( .A(n3636), .B(n3635), .Z(n3637) );
  NAND U4127 ( .A(n3638), .B(n3637), .Z(n3646) );
  XNOR U4128 ( .A(n3645), .B(n3646), .Z(n3648) );
  XOR U4129 ( .A(n3647), .B(n3648), .Z(n3639) );
  NANDN U4130 ( .A(n3640), .B(n3639), .Z(n3642) );
  XOR U4131 ( .A(n3640), .B(n3639), .Z(n17024) );
  AND U4132 ( .A(o[12]), .B(\stack[1][0] ), .Z(n17025) );
  OR U4133 ( .A(n17024), .B(n17025), .Z(n3641) );
  AND U4134 ( .A(n3642), .B(n3641), .Z(n3644) );
  OR U4135 ( .A(n3643), .B(n3644), .Z(n3711) );
  XNOR U4136 ( .A(n3644), .B(n3643), .Z(n16986) );
  NANDN U4137 ( .A(n2969), .B(o[12]), .Z(n3782) );
  OR U4138 ( .A(n3646), .B(n3645), .Z(n3650) );
  OR U4139 ( .A(n3648), .B(n3647), .Z(n3649) );
  NAND U4140 ( .A(n3650), .B(n3649), .Z(n3780) );
  NANDN U4141 ( .A(n17375), .B(o[10]), .Z(n3776) );
  OR U4142 ( .A(n3652), .B(n3651), .Z(n3656) );
  NANDN U4143 ( .A(n3654), .B(n3653), .Z(n3655) );
  NAND U4144 ( .A(n3656), .B(n3655), .Z(n3774) );
  NANDN U4145 ( .A(n17296), .B(o[8]), .Z(n3770) );
  OR U4146 ( .A(n3658), .B(n3657), .Z(n3662) );
  OR U4147 ( .A(n3660), .B(n3659), .Z(n3661) );
  NAND U4148 ( .A(n3662), .B(n3661), .Z(n3768) );
  NANDN U4149 ( .A(n3664), .B(n3663), .Z(n3667) );
  OR U4150 ( .A(n3665), .B(n17265), .Z(n3666) );
  AND U4151 ( .A(n3667), .B(n3666), .Z(n3724) );
  AND U4152 ( .A(o[7]), .B(\stack[1][6] ), .Z(n3725) );
  XNOR U4153 ( .A(n3724), .B(n3725), .Z(n3727) );
  OR U4154 ( .A(n3669), .B(n3668), .Z(n3673) );
  OR U4155 ( .A(n3671), .B(n3670), .Z(n3672) );
  AND U4156 ( .A(n3673), .B(n3672), .Z(n3731) );
  OR U4157 ( .A(n3675), .B(n3674), .Z(n3679) );
  OR U4158 ( .A(n3677), .B(n3676), .Z(n3678) );
  NAND U4159 ( .A(n3679), .B(n3678), .Z(n3762) );
  OR U4160 ( .A(n3681), .B(n3680), .Z(n3687) );
  ANDN U4161 ( .B(\stack[1][10] ), .A(n2994), .Z(n3682) );
  NANDN U4162 ( .A(n3683), .B(n3682), .Z(n3685) );
  NANDN U4163 ( .A(n17101), .B(o[2]), .Z(n3684) );
  AND U4164 ( .A(n3685), .B(n3684), .Z(n3686) );
  ANDN U4165 ( .B(n3687), .A(n3686), .Z(n3742) );
  AND U4166 ( .A(\stack[1][10] ), .B(o[3]), .Z(n3743) );
  XNOR U4167 ( .A(n3742), .B(n3743), .Z(n3745) );
  ANDN U4168 ( .B(o[0]), .A(n2974), .Z(n3689) );
  ANDN U4169 ( .B(o[1]), .A(n2973), .Z(n3688) );
  XOR U4170 ( .A(n3689), .B(n3688), .Z(n3748) );
  NANDN U4171 ( .A(n2995), .B(\stack[1][12] ), .Z(n3751) );
  OR U4172 ( .A(n3751), .B(n2994), .Z(n3690) );
  XOR U4173 ( .A(n2996), .B(n3690), .Z(n3691) );
  NANDN U4174 ( .A(n2972), .B(n3691), .Z(n3749) );
  XNOR U4175 ( .A(n3748), .B(n3749), .Z(n3744) );
  XOR U4176 ( .A(n3745), .B(n3744), .Z(n3761) );
  XNOR U4177 ( .A(n3762), .B(n3761), .Z(n3763) );
  NANDN U4178 ( .A(n2998), .B(\stack[1][9] ), .Z(n3764) );
  AND U4179 ( .A(\stack[1][8] ), .B(o[5]), .Z(n3736) );
  OR U4180 ( .A(n3693), .B(n3692), .Z(n3697) );
  OR U4181 ( .A(n3695), .B(n3694), .Z(n3696) );
  NAND U4182 ( .A(n3697), .B(n3696), .Z(n3737) );
  XNOR U4183 ( .A(n3736), .B(n3737), .Z(n3739) );
  XOR U4184 ( .A(n3738), .B(n3739), .Z(n3730) );
  XOR U4185 ( .A(n3731), .B(n3730), .Z(n3733) );
  AND U4186 ( .A(\stack[1][7] ), .B(o[6]), .Z(n3732) );
  XNOR U4187 ( .A(n3733), .B(n3732), .Z(n3726) );
  XOR U4188 ( .A(n3727), .B(n3726), .Z(n3767) );
  XNOR U4189 ( .A(n3768), .B(n3767), .Z(n3769) );
  AND U4190 ( .A(o[9]), .B(\stack[1][4] ), .Z(n3718) );
  OR U4191 ( .A(n3699), .B(n3698), .Z(n3703) );
  OR U4192 ( .A(n3701), .B(n3700), .Z(n3702) );
  NAND U4193 ( .A(n3703), .B(n3702), .Z(n3719) );
  XOR U4194 ( .A(n3718), .B(n3719), .Z(n3720) );
  XNOR U4195 ( .A(n3721), .B(n3720), .Z(n3773) );
  XNOR U4196 ( .A(n3774), .B(n3773), .Z(n3775) );
  XOR U4197 ( .A(n3776), .B(n3775), .Z(n3715) );
  AND U4198 ( .A(o[11]), .B(\stack[1][2] ), .Z(n3712) );
  OR U4199 ( .A(n3705), .B(n3704), .Z(n3709) );
  OR U4200 ( .A(n3707), .B(n3706), .Z(n3708) );
  NAND U4201 ( .A(n3709), .B(n3708), .Z(n3713) );
  XOR U4202 ( .A(n3712), .B(n3713), .Z(n3714) );
  XNOR U4203 ( .A(n3715), .B(n3714), .Z(n3779) );
  XNOR U4204 ( .A(n3780), .B(n3779), .Z(n3781) );
  XOR U4205 ( .A(n3782), .B(n3781), .Z(n16987) );
  OR U4206 ( .A(n16986), .B(n16987), .Z(n3710) );
  AND U4207 ( .A(n3711), .B(n3710), .Z(n3786) );
  NANDN U4208 ( .A(n2970), .B(o[12]), .Z(n3866) );
  OR U4209 ( .A(n3713), .B(n3712), .Z(n3717) );
  NANDN U4210 ( .A(n3715), .B(n3714), .Z(n3716) );
  NAND U4211 ( .A(n3717), .B(n3716), .Z(n3864) );
  NANDN U4212 ( .A(n2971), .B(o[10]), .Z(n3860) );
  OR U4213 ( .A(n3719), .B(n3718), .Z(n3723) );
  NANDN U4214 ( .A(n3721), .B(n3720), .Z(n3722) );
  NAND U4215 ( .A(n3723), .B(n3722), .Z(n3858) );
  NANDN U4216 ( .A(n17256), .B(o[8]), .Z(n3854) );
  OR U4217 ( .A(n3725), .B(n3724), .Z(n3729) );
  OR U4218 ( .A(n3727), .B(n3726), .Z(n3728) );
  NAND U4219 ( .A(n3729), .B(n3728), .Z(n3852) );
  AND U4220 ( .A(\stack[1][7] ), .B(o[7]), .Z(n3809) );
  NANDN U4221 ( .A(n3731), .B(n3730), .Z(n3735) );
  OR U4222 ( .A(n3733), .B(n3732), .Z(n3734) );
  AND U4223 ( .A(n3735), .B(n3734), .Z(n3810) );
  XNOR U4224 ( .A(n3809), .B(n3810), .Z(n3812) );
  OR U4225 ( .A(n3737), .B(n3736), .Z(n3741) );
  OR U4226 ( .A(n3739), .B(n3738), .Z(n3740) );
  AND U4227 ( .A(n3741), .B(n3740), .Z(n3816) );
  OR U4228 ( .A(n3743), .B(n3742), .Z(n3747) );
  OR U4229 ( .A(n3745), .B(n3744), .Z(n3746) );
  NAND U4230 ( .A(n3747), .B(n3746), .Z(n3846) );
  OR U4231 ( .A(n3749), .B(n3748), .Z(n3755) );
  ANDN U4232 ( .B(\stack[1][11] ), .A(n2994), .Z(n3750) );
  NANDN U4233 ( .A(n3751), .B(n3750), .Z(n3753) );
  NANDN U4234 ( .A(n2972), .B(o[2]), .Z(n3752) );
  AND U4235 ( .A(n3753), .B(n3752), .Z(n3754) );
  ANDN U4236 ( .B(n3755), .A(n3754), .Z(n3827) );
  AND U4237 ( .A(\stack[1][11] ), .B(o[3]), .Z(n3828) );
  XNOR U4238 ( .A(n3827), .B(n3828), .Z(n3830) );
  ANDN U4239 ( .B(o[0]), .A(n2975), .Z(n3757) );
  ANDN U4240 ( .B(o[1]), .A(n2974), .Z(n3756) );
  XOR U4241 ( .A(n3757), .B(n3756), .Z(n3833) );
  NANDN U4242 ( .A(n2995), .B(\stack[1][13] ), .Z(n3836) );
  OR U4243 ( .A(n3836), .B(n2994), .Z(n3758) );
  XOR U4244 ( .A(n2996), .B(n3758), .Z(n3759) );
  NANDN U4245 ( .A(n2973), .B(n3759), .Z(n3834) );
  XNOR U4246 ( .A(n3833), .B(n3834), .Z(n3829) );
  XOR U4247 ( .A(n3830), .B(n3829), .Z(n3845) );
  XNOR U4248 ( .A(n3846), .B(n3845), .Z(n3847) );
  IV U4249 ( .A(n3847), .Z(n3760) );
  NANDN U4250 ( .A(n2998), .B(\stack[1][10] ), .Z(n3848) );
  XNOR U4251 ( .A(n3760), .B(n3848), .Z(n3823) );
  AND U4252 ( .A(\stack[1][9] ), .B(o[5]), .Z(n3821) );
  OR U4253 ( .A(n3762), .B(n3761), .Z(n3766) );
  OR U4254 ( .A(n3764), .B(n3763), .Z(n3765) );
  NAND U4255 ( .A(n3766), .B(n3765), .Z(n3822) );
  XNOR U4256 ( .A(n3821), .B(n3822), .Z(n3824) );
  XOR U4257 ( .A(n3823), .B(n3824), .Z(n3815) );
  XOR U4258 ( .A(n3816), .B(n3815), .Z(n3818) );
  AND U4259 ( .A(\stack[1][8] ), .B(o[6]), .Z(n3817) );
  XNOR U4260 ( .A(n3818), .B(n3817), .Z(n3811) );
  XOR U4261 ( .A(n3812), .B(n3811), .Z(n3851) );
  XNOR U4262 ( .A(n3852), .B(n3851), .Z(n3853) );
  AND U4263 ( .A(o[9]), .B(\stack[1][5] ), .Z(n3803) );
  OR U4264 ( .A(n3768), .B(n3767), .Z(n3772) );
  OR U4265 ( .A(n3770), .B(n3769), .Z(n3771) );
  NAND U4266 ( .A(n3772), .B(n3771), .Z(n3804) );
  XOR U4267 ( .A(n3803), .B(n3804), .Z(n3805) );
  XNOR U4268 ( .A(n3806), .B(n3805), .Z(n3857) );
  XNOR U4269 ( .A(n3858), .B(n3857), .Z(n3859) );
  XOR U4270 ( .A(n3860), .B(n3859), .Z(n3800) );
  AND U4271 ( .A(o[11]), .B(\stack[1][3] ), .Z(n3797) );
  OR U4272 ( .A(n3774), .B(n3773), .Z(n3778) );
  OR U4273 ( .A(n3776), .B(n3775), .Z(n3777) );
  NAND U4274 ( .A(n3778), .B(n3777), .Z(n3798) );
  XOR U4275 ( .A(n3797), .B(n3798), .Z(n3799) );
  XNOR U4276 ( .A(n3800), .B(n3799), .Z(n3863) );
  XNOR U4277 ( .A(n3864), .B(n3863), .Z(n3865) );
  XOR U4278 ( .A(n3866), .B(n3865), .Z(n3793) );
  AND U4279 ( .A(o[13]), .B(\stack[1][1] ), .Z(n3791) );
  OR U4280 ( .A(n3780), .B(n3779), .Z(n3784) );
  OR U4281 ( .A(n3782), .B(n3781), .Z(n3783) );
  NAND U4282 ( .A(n3784), .B(n3783), .Z(n3792) );
  XNOR U4283 ( .A(n3791), .B(n3792), .Z(n3794) );
  XOR U4284 ( .A(n3793), .B(n3794), .Z(n3785) );
  NANDN U4285 ( .A(n3786), .B(n3785), .Z(n3788) );
  XOR U4286 ( .A(n3786), .B(n3785), .Z(n16947) );
  AND U4287 ( .A(o[14]), .B(\stack[1][0] ), .Z(n16948) );
  OR U4288 ( .A(n16947), .B(n16948), .Z(n3787) );
  AND U4289 ( .A(n3788), .B(n3787), .Z(n3790) );
  OR U4290 ( .A(n3789), .B(n3790), .Z(n3870) );
  XNOR U4291 ( .A(n3790), .B(n3789), .Z(n16908) );
  NANDN U4292 ( .A(n2969), .B(o[14]), .Z(n3952) );
  OR U4293 ( .A(n3792), .B(n3791), .Z(n3796) );
  OR U4294 ( .A(n3794), .B(n3793), .Z(n3795) );
  NAND U4295 ( .A(n3796), .B(n3795), .Z(n3950) );
  NANDN U4296 ( .A(n17375), .B(o[12]), .Z(n3946) );
  OR U4297 ( .A(n3798), .B(n3797), .Z(n3802) );
  NANDN U4298 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U4299 ( .A(n3802), .B(n3801), .Z(n3944) );
  NANDN U4300 ( .A(n17296), .B(o[10]), .Z(n3940) );
  OR U4301 ( .A(n3804), .B(n3803), .Z(n3808) );
  NANDN U4302 ( .A(n3806), .B(n3805), .Z(n3807) );
  NAND U4303 ( .A(n3808), .B(n3807), .Z(n3938) );
  NANDN U4304 ( .A(n17219), .B(o[8]), .Z(n3934) );
  OR U4305 ( .A(n3810), .B(n3809), .Z(n3814) );
  OR U4306 ( .A(n3812), .B(n3811), .Z(n3813) );
  NAND U4307 ( .A(n3814), .B(n3813), .Z(n3932) );
  NANDN U4308 ( .A(n3816), .B(n3815), .Z(n3820) );
  OR U4309 ( .A(n3818), .B(n3817), .Z(n3819) );
  AND U4310 ( .A(n3820), .B(n3819), .Z(n3889) );
  AND U4311 ( .A(\stack[1][8] ), .B(o[7]), .Z(n3890) );
  XNOR U4312 ( .A(n3889), .B(n3890), .Z(n3892) );
  OR U4313 ( .A(n3822), .B(n3821), .Z(n3826) );
  OR U4314 ( .A(n3824), .B(n3823), .Z(n3825) );
  AND U4315 ( .A(n3826), .B(n3825), .Z(n3896) );
  OR U4316 ( .A(n3828), .B(n3827), .Z(n3832) );
  OR U4317 ( .A(n3830), .B(n3829), .Z(n3831) );
  NAND U4318 ( .A(n3832), .B(n3831), .Z(n3926) );
  OR U4319 ( .A(n3834), .B(n3833), .Z(n3840) );
  ANDN U4320 ( .B(\stack[1][12] ), .A(n2994), .Z(n3835) );
  NANDN U4321 ( .A(n3836), .B(n3835), .Z(n3838) );
  NANDN U4322 ( .A(n2973), .B(o[2]), .Z(n3837) );
  AND U4323 ( .A(n3838), .B(n3837), .Z(n3839) );
  ANDN U4324 ( .B(n3840), .A(n3839), .Z(n3907) );
  AND U4325 ( .A(\stack[1][12] ), .B(o[3]), .Z(n3908) );
  XNOR U4326 ( .A(n3907), .B(n3908), .Z(n3910) );
  ANDN U4327 ( .B(o[0]), .A(n2976), .Z(n3841) );
  NANDN U4328 ( .A(n2995), .B(\stack[1][14] ), .Z(n3916) );
  XNOR U4329 ( .A(n3841), .B(n3916), .Z(n3913) );
  OR U4330 ( .A(n3916), .B(n2994), .Z(n3842) );
  XOR U4331 ( .A(n2996), .B(n3842), .Z(n3843) );
  NANDN U4332 ( .A(n2974), .B(n3843), .Z(n3914) );
  XNOR U4333 ( .A(n3913), .B(n3914), .Z(n3909) );
  XNOR U4334 ( .A(n3926), .B(n3925), .Z(n3927) );
  IV U4335 ( .A(n3927), .Z(n3844) );
  NANDN U4336 ( .A(n2998), .B(\stack[1][11] ), .Z(n3928) );
  XNOR U4337 ( .A(n3844), .B(n3928), .Z(n3903) );
  AND U4338 ( .A(\stack[1][10] ), .B(o[5]), .Z(n3901) );
  OR U4339 ( .A(n3846), .B(n3845), .Z(n3850) );
  OR U4340 ( .A(n3848), .B(n3847), .Z(n3849) );
  NAND U4341 ( .A(n3850), .B(n3849), .Z(n3902) );
  XNOR U4342 ( .A(n3901), .B(n3902), .Z(n3904) );
  XOR U4343 ( .A(n3903), .B(n3904), .Z(n3895) );
  XOR U4344 ( .A(n3896), .B(n3895), .Z(n3898) );
  AND U4345 ( .A(\stack[1][9] ), .B(o[6]), .Z(n3897) );
  XNOR U4346 ( .A(n3898), .B(n3897), .Z(n3891) );
  XOR U4347 ( .A(n3892), .B(n3891), .Z(n3931) );
  XNOR U4348 ( .A(n3932), .B(n3931), .Z(n3933) );
  AND U4349 ( .A(o[9]), .B(\stack[1][6] ), .Z(n3883) );
  OR U4350 ( .A(n3852), .B(n3851), .Z(n3856) );
  OR U4351 ( .A(n3854), .B(n3853), .Z(n3855) );
  NAND U4352 ( .A(n3856), .B(n3855), .Z(n3884) );
  XOR U4353 ( .A(n3883), .B(n3884), .Z(n3885) );
  XNOR U4354 ( .A(n3886), .B(n3885), .Z(n3937) );
  XNOR U4355 ( .A(n3938), .B(n3937), .Z(n3939) );
  XOR U4356 ( .A(n3940), .B(n3939), .Z(n3880) );
  AND U4357 ( .A(o[11]), .B(\stack[1][4] ), .Z(n3877) );
  OR U4358 ( .A(n3858), .B(n3857), .Z(n3862) );
  OR U4359 ( .A(n3860), .B(n3859), .Z(n3861) );
  NAND U4360 ( .A(n3862), .B(n3861), .Z(n3878) );
  XOR U4361 ( .A(n3877), .B(n3878), .Z(n3879) );
  XNOR U4362 ( .A(n3880), .B(n3879), .Z(n3943) );
  XNOR U4363 ( .A(n3944), .B(n3943), .Z(n3945) );
  XOR U4364 ( .A(n3946), .B(n3945), .Z(n3874) );
  AND U4365 ( .A(o[13]), .B(\stack[1][2] ), .Z(n3871) );
  OR U4366 ( .A(n3864), .B(n3863), .Z(n3868) );
  OR U4367 ( .A(n3866), .B(n3865), .Z(n3867) );
  NAND U4368 ( .A(n3868), .B(n3867), .Z(n3872) );
  XOR U4369 ( .A(n3871), .B(n3872), .Z(n3873) );
  XNOR U4370 ( .A(n3874), .B(n3873), .Z(n3949) );
  XNOR U4371 ( .A(n3950), .B(n3949), .Z(n3951) );
  XOR U4372 ( .A(n3952), .B(n3951), .Z(n16909) );
  OR U4373 ( .A(n16908), .B(n16909), .Z(n3869) );
  AND U4374 ( .A(n3870), .B(n3869), .Z(n3956) );
  NANDN U4375 ( .A(n2970), .B(o[14]), .Z(n4047) );
  OR U4376 ( .A(n3872), .B(n3871), .Z(n3876) );
  NANDN U4377 ( .A(n3874), .B(n3873), .Z(n3875) );
  NAND U4378 ( .A(n3876), .B(n3875), .Z(n4045) );
  NANDN U4379 ( .A(n2971), .B(o[12]), .Z(n4041) );
  OR U4380 ( .A(n3878), .B(n3877), .Z(n3882) );
  NANDN U4381 ( .A(n3880), .B(n3879), .Z(n3881) );
  NAND U4382 ( .A(n3882), .B(n3881), .Z(n4039) );
  NANDN U4383 ( .A(n17256), .B(o[10]), .Z(n4035) );
  OR U4384 ( .A(n3884), .B(n3883), .Z(n3888) );
  NANDN U4385 ( .A(n3886), .B(n3885), .Z(n3887) );
  NAND U4386 ( .A(n3888), .B(n3887), .Z(n4033) );
  AND U4387 ( .A(o[8]), .B(\stack[1][8] ), .Z(n17180) );
  OR U4388 ( .A(n3890), .B(n3889), .Z(n3894) );
  OR U4389 ( .A(n3892), .B(n3891), .Z(n3893) );
  NAND U4390 ( .A(n3894), .B(n3893), .Z(n4028) );
  NANDN U4391 ( .A(n3896), .B(n3895), .Z(n3900) );
  OR U4392 ( .A(n3898), .B(n3897), .Z(n3899) );
  AND U4393 ( .A(n3900), .B(n3899), .Z(n3985) );
  AND U4394 ( .A(\stack[1][9] ), .B(o[7]), .Z(n3986) );
  XNOR U4395 ( .A(n3985), .B(n3986), .Z(n3988) );
  OR U4396 ( .A(n3902), .B(n3901), .Z(n3906) );
  OR U4397 ( .A(n3904), .B(n3903), .Z(n3905) );
  AND U4398 ( .A(n3906), .B(n3905), .Z(n3991) );
  OR U4399 ( .A(n3908), .B(n3907), .Z(n3912) );
  OR U4400 ( .A(n3910), .B(n3909), .Z(n3911) );
  NAND U4401 ( .A(n3912), .B(n3911), .Z(n4022) );
  OR U4402 ( .A(n3914), .B(n3913), .Z(n3920) );
  ANDN U4403 ( .B(\stack[1][13] ), .A(n2994), .Z(n3915) );
  NANDN U4404 ( .A(n3916), .B(n3915), .Z(n3918) );
  NANDN U4405 ( .A(n2974), .B(o[2]), .Z(n3917) );
  AND U4406 ( .A(n3918), .B(n3917), .Z(n3919) );
  ANDN U4407 ( .B(n3920), .A(n3919), .Z(n4003) );
  AND U4408 ( .A(\stack[1][13] ), .B(o[3]), .Z(n4004) );
  XNOR U4409 ( .A(n4003), .B(n4004), .Z(n4006) );
  ANDN U4410 ( .B(o[0]), .A(n2977), .Z(n3922) );
  NANDN U4411 ( .A(n2995), .B(\stack[1][15] ), .Z(n3921) );
  XNOR U4412 ( .A(n3922), .B(n3921), .Z(n4010) );
  AND U4413 ( .A(\stack[1][15] ), .B(o[1]), .Z(n4011) );
  NANDN U4414 ( .A(n2994), .B(n4011), .Z(n3923) );
  XOR U4415 ( .A(n2996), .B(n3923), .Z(n3924) );
  AND U4416 ( .A(n3924), .B(\stack[1][14] ), .Z(n4009) );
  XOR U4417 ( .A(n4010), .B(n4009), .Z(n4005) );
  XOR U4418 ( .A(n4006), .B(n4005), .Z(n4021) );
  XNOR U4419 ( .A(n4022), .B(n4021), .Z(n4024) );
  AND U4420 ( .A(\stack[1][12] ), .B(o[4]), .Z(n4023) );
  XNOR U4421 ( .A(n4024), .B(n4023), .Z(n3999) );
  AND U4422 ( .A(\stack[1][11] ), .B(o[5]), .Z(n3997) );
  OR U4423 ( .A(n3926), .B(n3925), .Z(n3930) );
  OR U4424 ( .A(n3928), .B(n3927), .Z(n3929) );
  NAND U4425 ( .A(n3930), .B(n3929), .Z(n3998) );
  XNOR U4426 ( .A(n3997), .B(n3998), .Z(n4000) );
  XNOR U4427 ( .A(n3999), .B(n4000), .Z(n3992) );
  XNOR U4428 ( .A(n3991), .B(n3992), .Z(n3994) );
  AND U4429 ( .A(\stack[1][10] ), .B(o[6]), .Z(n3993) );
  XNOR U4430 ( .A(n3994), .B(n3993), .Z(n3987) );
  XOR U4431 ( .A(n3988), .B(n3987), .Z(n4027) );
  XNOR U4432 ( .A(n4028), .B(n4027), .Z(n4029) );
  AND U4433 ( .A(o[9]), .B(\stack[1][7] ), .Z(n3979) );
  OR U4434 ( .A(n3932), .B(n3931), .Z(n3936) );
  OR U4435 ( .A(n3934), .B(n3933), .Z(n3935) );
  NAND U4436 ( .A(n3936), .B(n3935), .Z(n3980) );
  XOR U4437 ( .A(n3979), .B(n3980), .Z(n3981) );
  XNOR U4438 ( .A(n3982), .B(n3981), .Z(n4032) );
  XNOR U4439 ( .A(n4033), .B(n4032), .Z(n4034) );
  XOR U4440 ( .A(n4035), .B(n4034), .Z(n3976) );
  AND U4441 ( .A(o[11]), .B(\stack[1][5] ), .Z(n3973) );
  OR U4442 ( .A(n3938), .B(n3937), .Z(n3942) );
  OR U4443 ( .A(n3940), .B(n3939), .Z(n3941) );
  NAND U4444 ( .A(n3942), .B(n3941), .Z(n3974) );
  XOR U4445 ( .A(n3973), .B(n3974), .Z(n3975) );
  XNOR U4446 ( .A(n3976), .B(n3975), .Z(n4038) );
  XNOR U4447 ( .A(n4039), .B(n4038), .Z(n4040) );
  XOR U4448 ( .A(n4041), .B(n4040), .Z(n3970) );
  AND U4449 ( .A(o[13]), .B(\stack[1][3] ), .Z(n3967) );
  OR U4450 ( .A(n3944), .B(n3943), .Z(n3948) );
  OR U4451 ( .A(n3946), .B(n3945), .Z(n3947) );
  NAND U4452 ( .A(n3948), .B(n3947), .Z(n3968) );
  XOR U4453 ( .A(n3967), .B(n3968), .Z(n3969) );
  XNOR U4454 ( .A(n3970), .B(n3969), .Z(n4044) );
  XNOR U4455 ( .A(n4045), .B(n4044), .Z(n4046) );
  XOR U4456 ( .A(n4047), .B(n4046), .Z(n3963) );
  AND U4457 ( .A(o[15]), .B(\stack[1][1] ), .Z(n3961) );
  OR U4458 ( .A(n3950), .B(n3949), .Z(n3954) );
  OR U4459 ( .A(n3952), .B(n3951), .Z(n3953) );
  NAND U4460 ( .A(n3954), .B(n3953), .Z(n3962) );
  XNOR U4461 ( .A(n3961), .B(n3962), .Z(n3964) );
  XOR U4462 ( .A(n3963), .B(n3964), .Z(n3955) );
  NANDN U4463 ( .A(n3956), .B(n3955), .Z(n3958) );
  XOR U4464 ( .A(n3956), .B(n3955), .Z(n16866) );
  AND U4465 ( .A(o[16]), .B(\stack[1][0] ), .Z(n16867) );
  OR U4466 ( .A(n16866), .B(n16867), .Z(n3957) );
  AND U4467 ( .A(n3958), .B(n3957), .Z(n3960) );
  OR U4468 ( .A(n3959), .B(n3960), .Z(n4051) );
  XNOR U4469 ( .A(n3960), .B(n3959), .Z(n16830) );
  NANDN U4470 ( .A(n2969), .B(o[16]), .Z(n4145) );
  OR U4471 ( .A(n3962), .B(n3961), .Z(n3966) );
  OR U4472 ( .A(n3964), .B(n3963), .Z(n3965) );
  NAND U4473 ( .A(n3966), .B(n3965), .Z(n4143) );
  NANDN U4474 ( .A(n17375), .B(o[14]), .Z(n4139) );
  OR U4475 ( .A(n3968), .B(n3967), .Z(n3972) );
  NANDN U4476 ( .A(n3970), .B(n3969), .Z(n3971) );
  NAND U4477 ( .A(n3972), .B(n3971), .Z(n4137) );
  NANDN U4478 ( .A(n17296), .B(o[12]), .Z(n4133) );
  OR U4479 ( .A(n3974), .B(n3973), .Z(n3978) );
  NANDN U4480 ( .A(n3976), .B(n3975), .Z(n3977) );
  NAND U4481 ( .A(n3978), .B(n3977), .Z(n4131) );
  NANDN U4482 ( .A(n17219), .B(o[10]), .Z(n4073) );
  OR U4483 ( .A(n3980), .B(n3979), .Z(n3984) );
  NANDN U4484 ( .A(n3982), .B(n3981), .Z(n3983) );
  NAND U4485 ( .A(n3984), .B(n3983), .Z(n4071) );
  NANDN U4486 ( .A(n3002), .B(\stack[1][9] ), .Z(n4127) );
  OR U4487 ( .A(n3986), .B(n3985), .Z(n3990) );
  OR U4488 ( .A(n3988), .B(n3987), .Z(n3989) );
  NAND U4489 ( .A(n3990), .B(n3989), .Z(n4125) );
  OR U4490 ( .A(n3992), .B(n3991), .Z(n3996) );
  OR U4491 ( .A(n3994), .B(n3993), .Z(n3995) );
  AND U4492 ( .A(n3996), .B(n3995), .Z(n4082) );
  AND U4493 ( .A(\stack[1][10] ), .B(o[7]), .Z(n4083) );
  XNOR U4494 ( .A(n4082), .B(n4083), .Z(n4085) );
  OR U4495 ( .A(n3998), .B(n3997), .Z(n4002) );
  OR U4496 ( .A(n4000), .B(n3999), .Z(n4001) );
  AND U4497 ( .A(n4002), .B(n4001), .Z(n4088) );
  OR U4498 ( .A(n4004), .B(n4003), .Z(n4008) );
  OR U4499 ( .A(n4006), .B(n4005), .Z(n4007) );
  NAND U4500 ( .A(n4008), .B(n4007), .Z(n4119) );
  NANDN U4501 ( .A(n4010), .B(n4009), .Z(n4016) );
  ANDN U4502 ( .B(\stack[1][14] ), .A(n2994), .Z(n4012) );
  NAND U4503 ( .A(n4012), .B(n4011), .Z(n4014) );
  NANDN U4504 ( .A(n2975), .B(o[2]), .Z(n4013) );
  AND U4505 ( .A(n4014), .B(n4013), .Z(n4015) );
  ANDN U4506 ( .B(n4016), .A(n4015), .Z(n4100) );
  AND U4507 ( .A(\stack[1][14] ), .B(o[3]), .Z(n4101) );
  XNOR U4508 ( .A(n4100), .B(n4101), .Z(n4103) );
  IV U4509 ( .A(\stack[1][17] ), .Z(n16826) );
  ANDN U4510 ( .B(o[0]), .A(n16826), .Z(n4018) );
  NANDN U4511 ( .A(n2995), .B(\stack[1][16] ), .Z(n4017) );
  XNOR U4512 ( .A(n4018), .B(n4017), .Z(n4107) );
  AND U4513 ( .A(\stack[1][16] ), .B(o[1]), .Z(n4108) );
  NANDN U4514 ( .A(n2994), .B(n4108), .Z(n4019) );
  XOR U4515 ( .A(n2996), .B(n4019), .Z(n4020) );
  AND U4516 ( .A(n4020), .B(\stack[1][15] ), .Z(n4106) );
  XOR U4517 ( .A(n4107), .B(n4106), .Z(n4102) );
  XOR U4518 ( .A(n4103), .B(n4102), .Z(n4118) );
  XNOR U4519 ( .A(n4119), .B(n4118), .Z(n4121) );
  AND U4520 ( .A(\stack[1][13] ), .B(o[4]), .Z(n4120) );
  XNOR U4521 ( .A(n4121), .B(n4120), .Z(n4096) );
  AND U4522 ( .A(\stack[1][12] ), .B(o[5]), .Z(n4094) );
  OR U4523 ( .A(n4022), .B(n4021), .Z(n4026) );
  NANDN U4524 ( .A(n4024), .B(n4023), .Z(n4025) );
  NAND U4525 ( .A(n4026), .B(n4025), .Z(n4095) );
  XNOR U4526 ( .A(n4094), .B(n4095), .Z(n4097) );
  XNOR U4527 ( .A(n4096), .B(n4097), .Z(n4089) );
  XOR U4528 ( .A(n4088), .B(n4089), .Z(n4090) );
  AND U4529 ( .A(\stack[1][11] ), .B(o[6]), .Z(n4091) );
  XOR U4530 ( .A(n4090), .B(n4091), .Z(n4084) );
  XOR U4531 ( .A(n4085), .B(n4084), .Z(n4124) );
  XNOR U4532 ( .A(n4125), .B(n4124), .Z(n4126) );
  AND U4533 ( .A(o[9]), .B(\stack[1][8] ), .Z(n4076) );
  OR U4534 ( .A(n4028), .B(n4027), .Z(n4031) );
  NANDN U4535 ( .A(n4029), .B(n17180), .Z(n4030) );
  NAND U4536 ( .A(n4031), .B(n4030), .Z(n4077) );
  XOR U4537 ( .A(n4076), .B(n4077), .Z(n4078) );
  XNOR U4538 ( .A(n4079), .B(n4078), .Z(n4070) );
  XNOR U4539 ( .A(n4071), .B(n4070), .Z(n4072) );
  XOR U4540 ( .A(n4073), .B(n4072), .Z(n4067) );
  AND U4541 ( .A(o[11]), .B(\stack[1][6] ), .Z(n4064) );
  OR U4542 ( .A(n4033), .B(n4032), .Z(n4037) );
  OR U4543 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4544 ( .A(n4037), .B(n4036), .Z(n4065) );
  XOR U4545 ( .A(n4064), .B(n4065), .Z(n4066) );
  XNOR U4546 ( .A(n4067), .B(n4066), .Z(n4130) );
  XNOR U4547 ( .A(n4131), .B(n4130), .Z(n4132) );
  XOR U4548 ( .A(n4133), .B(n4132), .Z(n4061) );
  AND U4549 ( .A(o[13]), .B(\stack[1][4] ), .Z(n4058) );
  OR U4550 ( .A(n4039), .B(n4038), .Z(n4043) );
  OR U4551 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U4552 ( .A(n4043), .B(n4042), .Z(n4059) );
  XOR U4553 ( .A(n4058), .B(n4059), .Z(n4060) );
  XNOR U4554 ( .A(n4061), .B(n4060), .Z(n4136) );
  XNOR U4555 ( .A(n4137), .B(n4136), .Z(n4138) );
  XOR U4556 ( .A(n4139), .B(n4138), .Z(n4055) );
  AND U4557 ( .A(o[15]), .B(\stack[1][2] ), .Z(n4052) );
  OR U4558 ( .A(n4045), .B(n4044), .Z(n4049) );
  OR U4559 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4560 ( .A(n4049), .B(n4048), .Z(n4053) );
  XOR U4561 ( .A(n4052), .B(n4053), .Z(n4054) );
  XNOR U4562 ( .A(n4055), .B(n4054), .Z(n4142) );
  XNOR U4563 ( .A(n4143), .B(n4142), .Z(n4144) );
  XOR U4564 ( .A(n4145), .B(n4144), .Z(n16831) );
  OR U4565 ( .A(n16830), .B(n16831), .Z(n4050) );
  AND U4566 ( .A(n4051), .B(n4050), .Z(n4149) );
  NANDN U4567 ( .A(n2970), .B(o[16]), .Z(n4252) );
  OR U4568 ( .A(n4053), .B(n4052), .Z(n4057) );
  NANDN U4569 ( .A(n4055), .B(n4054), .Z(n4056) );
  NAND U4570 ( .A(n4057), .B(n4056), .Z(n4250) );
  NANDN U4571 ( .A(n2971), .B(o[14]), .Z(n4169) );
  OR U4572 ( .A(n4059), .B(n4058), .Z(n4063) );
  NANDN U4573 ( .A(n4061), .B(n4060), .Z(n4062) );
  NAND U4574 ( .A(n4063), .B(n4062), .Z(n4167) );
  AND U4575 ( .A(o[12]), .B(\stack[1][6] ), .Z(n4245) );
  OR U4576 ( .A(n4065), .B(n4064), .Z(n4069) );
  NANDN U4577 ( .A(n4067), .B(n4066), .Z(n4068) );
  AND U4578 ( .A(n4069), .B(n4068), .Z(n4244) );
  AND U4579 ( .A(o[11]), .B(\stack[1][7] ), .Z(n4178) );
  OR U4580 ( .A(n4071), .B(n4070), .Z(n4075) );
  OR U4581 ( .A(n4073), .B(n4072), .Z(n4074) );
  NAND U4582 ( .A(n4075), .B(n4074), .Z(n4179) );
  XNOR U4583 ( .A(n4178), .B(n4179), .Z(n4181) );
  OR U4584 ( .A(n4077), .B(n4076), .Z(n4081) );
  NANDN U4585 ( .A(n4079), .B(n4078), .Z(n4080) );
  AND U4586 ( .A(n4081), .B(n4080), .Z(n4238) );
  OR U4587 ( .A(n4083), .B(n4082), .Z(n4087) );
  OR U4588 ( .A(n4085), .B(n4084), .Z(n4086) );
  NAND U4589 ( .A(n4087), .B(n4086), .Z(n4232) );
  OR U4590 ( .A(n4089), .B(n4088), .Z(n4093) );
  NANDN U4591 ( .A(n4091), .B(n4090), .Z(n4092) );
  AND U4592 ( .A(n4093), .B(n4092), .Z(n4189) );
  AND U4593 ( .A(\stack[1][11] ), .B(o[7]), .Z(n4190) );
  XNOR U4594 ( .A(n4189), .B(n4190), .Z(n4192) );
  OR U4595 ( .A(n4095), .B(n4094), .Z(n4099) );
  OR U4596 ( .A(n4097), .B(n4096), .Z(n4098) );
  AND U4597 ( .A(n4099), .B(n4098), .Z(n4195) );
  OR U4598 ( .A(n4101), .B(n4100), .Z(n4105) );
  OR U4599 ( .A(n4103), .B(n4102), .Z(n4104) );
  NAND U4600 ( .A(n4105), .B(n4104), .Z(n4226) );
  NANDN U4601 ( .A(n4107), .B(n4106), .Z(n4113) );
  ANDN U4602 ( .B(\stack[1][15] ), .A(n2994), .Z(n4109) );
  NAND U4603 ( .A(n4109), .B(n4108), .Z(n4111) );
  NANDN U4604 ( .A(n2976), .B(o[2]), .Z(n4110) );
  AND U4605 ( .A(n4111), .B(n4110), .Z(n4112) );
  ANDN U4606 ( .B(n4113), .A(n4112), .Z(n4207) );
  AND U4607 ( .A(\stack[1][15] ), .B(o[3]), .Z(n4208) );
  XNOR U4608 ( .A(n4207), .B(n4208), .Z(n4210) );
  IV U4609 ( .A(\stack[1][18] ), .Z(n16786) );
  ANDN U4610 ( .B(o[0]), .A(n16786), .Z(n4115) );
  NANDN U4611 ( .A(n2995), .B(\stack[1][17] ), .Z(n4114) );
  XNOR U4612 ( .A(n4115), .B(n4114), .Z(n4214) );
  AND U4613 ( .A(\stack[1][17] ), .B(o[1]), .Z(n4215) );
  NANDN U4614 ( .A(n2994), .B(n4215), .Z(n4116) );
  XOR U4615 ( .A(n2996), .B(n4116), .Z(n4117) );
  AND U4616 ( .A(n4117), .B(\stack[1][16] ), .Z(n4213) );
  XOR U4617 ( .A(n4214), .B(n4213), .Z(n4209) );
  XOR U4618 ( .A(n4210), .B(n4209), .Z(n4225) );
  XNOR U4619 ( .A(n4226), .B(n4225), .Z(n4228) );
  AND U4620 ( .A(\stack[1][14] ), .B(o[4]), .Z(n4227) );
  XNOR U4621 ( .A(n4228), .B(n4227), .Z(n4203) );
  AND U4622 ( .A(\stack[1][13] ), .B(o[5]), .Z(n4201) );
  OR U4623 ( .A(n4119), .B(n4118), .Z(n4123) );
  NANDN U4624 ( .A(n4121), .B(n4120), .Z(n4122) );
  NAND U4625 ( .A(n4123), .B(n4122), .Z(n4202) );
  XNOR U4626 ( .A(n4201), .B(n4202), .Z(n4204) );
  XNOR U4627 ( .A(n4203), .B(n4204), .Z(n4196) );
  XOR U4628 ( .A(n4195), .B(n4196), .Z(n4197) );
  AND U4629 ( .A(\stack[1][12] ), .B(o[6]), .Z(n4198) );
  XOR U4630 ( .A(n4197), .B(n4198), .Z(n4191) );
  XOR U4631 ( .A(n4192), .B(n4191), .Z(n4231) );
  XNOR U4632 ( .A(n4232), .B(n4231), .Z(n4233) );
  NANDN U4633 ( .A(n3002), .B(\stack[1][10] ), .Z(n4234) );
  AND U4634 ( .A(\stack[1][9] ), .B(o[9]), .Z(n17139) );
  OR U4635 ( .A(n4125), .B(n4124), .Z(n4129) );
  OR U4636 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND U4637 ( .A(n4129), .B(n4128), .Z(n4184) );
  XNOR U4638 ( .A(n17139), .B(n4184), .Z(n4186) );
  XOR U4639 ( .A(n4185), .B(n4186), .Z(n4237) );
  XOR U4640 ( .A(n4238), .B(n4237), .Z(n4240) );
  AND U4641 ( .A(o[10]), .B(\stack[1][8] ), .Z(n4239) );
  XNOR U4642 ( .A(n4240), .B(n4239), .Z(n4180) );
  XOR U4643 ( .A(n4244), .B(n4243), .Z(n4246) );
  XNOR U4644 ( .A(n4245), .B(n4246), .Z(n4175) );
  AND U4645 ( .A(o[13]), .B(\stack[1][5] ), .Z(n4172) );
  OR U4646 ( .A(n4131), .B(n4130), .Z(n4135) );
  OR U4647 ( .A(n4133), .B(n4132), .Z(n4134) );
  NAND U4648 ( .A(n4135), .B(n4134), .Z(n4173) );
  XNOR U4649 ( .A(n4172), .B(n4173), .Z(n4174) );
  XOR U4650 ( .A(n4175), .B(n4174), .Z(n4166) );
  XNOR U4651 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U4652 ( .A(o[15]), .B(\stack[1][3] ), .Z(n4160) );
  OR U4653 ( .A(n4137), .B(n4136), .Z(n4141) );
  OR U4654 ( .A(n4139), .B(n4138), .Z(n4140) );
  NAND U4655 ( .A(n4141), .B(n4140), .Z(n4161) );
  XOR U4656 ( .A(n4160), .B(n4161), .Z(n4162) );
  XNOR U4657 ( .A(n4163), .B(n4162), .Z(n4249) );
  XNOR U4658 ( .A(n4250), .B(n4249), .Z(n4251) );
  XOR U4659 ( .A(n4252), .B(n4251), .Z(n4156) );
  AND U4660 ( .A(o[17]), .B(\stack[1][1] ), .Z(n4154) );
  OR U4661 ( .A(n4143), .B(n4142), .Z(n4147) );
  OR U4662 ( .A(n4145), .B(n4144), .Z(n4146) );
  NAND U4663 ( .A(n4147), .B(n4146), .Z(n4155) );
  XNOR U4664 ( .A(n4154), .B(n4155), .Z(n4157) );
  XOR U4665 ( .A(n4156), .B(n4157), .Z(n4148) );
  NANDN U4666 ( .A(n4149), .B(n4148), .Z(n4151) );
  XOR U4667 ( .A(n4149), .B(n4148), .Z(n16790) );
  AND U4668 ( .A(o[18]), .B(\stack[1][0] ), .Z(n16791) );
  OR U4669 ( .A(n16790), .B(n16791), .Z(n4150) );
  AND U4670 ( .A(n4151), .B(n4150), .Z(n4153) );
  OR U4671 ( .A(n4152), .B(n4153), .Z(n4256) );
  XNOR U4672 ( .A(n4153), .B(n4152), .Z(n16750) );
  NANDN U4673 ( .A(n2969), .B(o[18]), .Z(n4260) );
  OR U4674 ( .A(n4155), .B(n4154), .Z(n4159) );
  OR U4675 ( .A(n4157), .B(n4156), .Z(n4158) );
  NAND U4676 ( .A(n4159), .B(n4158), .Z(n4258) );
  AND U4677 ( .A(o[16]), .B(\stack[1][3] ), .Z(n4361) );
  OR U4678 ( .A(n4161), .B(n4160), .Z(n4165) );
  NANDN U4679 ( .A(n4163), .B(n4162), .Z(n4164) );
  AND U4680 ( .A(n4165), .B(n4164), .Z(n4360) );
  AND U4681 ( .A(o[15]), .B(\stack[1][4] ), .Z(n4269) );
  OR U4682 ( .A(n4167), .B(n4166), .Z(n4171) );
  OR U4683 ( .A(n4169), .B(n4168), .Z(n4170) );
  NAND U4684 ( .A(n4171), .B(n4170), .Z(n4270) );
  XNOR U4685 ( .A(n4269), .B(n4270), .Z(n4272) );
  OR U4686 ( .A(n4173), .B(n4172), .Z(n4177) );
  OR U4687 ( .A(n4175), .B(n4174), .Z(n4176) );
  AND U4688 ( .A(n4177), .B(n4176), .Z(n4354) );
  OR U4689 ( .A(n4179), .B(n4178), .Z(n4183) );
  OR U4690 ( .A(n4181), .B(n4180), .Z(n4182) );
  NAND U4691 ( .A(n4183), .B(n4182), .Z(n4348) );
  NANDN U4692 ( .A(n17145), .B(o[10]), .Z(n4344) );
  OR U4693 ( .A(n4184), .B(n17139), .Z(n4188) );
  OR U4694 ( .A(n4186), .B(n4185), .Z(n4187) );
  NAND U4695 ( .A(n4188), .B(n4187), .Z(n4342) );
  NANDN U4696 ( .A(n3002), .B(\stack[1][11] ), .Z(n4338) );
  OR U4697 ( .A(n4190), .B(n4189), .Z(n4194) );
  OR U4698 ( .A(n4192), .B(n4191), .Z(n4193) );
  NAND U4699 ( .A(n4194), .B(n4193), .Z(n4336) );
  OR U4700 ( .A(n4196), .B(n4195), .Z(n4200) );
  NANDN U4701 ( .A(n4198), .B(n4197), .Z(n4199) );
  AND U4702 ( .A(n4200), .B(n4199), .Z(n4293) );
  AND U4703 ( .A(\stack[1][12] ), .B(o[7]), .Z(n4294) );
  XNOR U4704 ( .A(n4293), .B(n4294), .Z(n4296) );
  OR U4705 ( .A(n4202), .B(n4201), .Z(n4206) );
  OR U4706 ( .A(n4204), .B(n4203), .Z(n4205) );
  AND U4707 ( .A(n4206), .B(n4205), .Z(n4299) );
  OR U4708 ( .A(n4208), .B(n4207), .Z(n4212) );
  OR U4709 ( .A(n4210), .B(n4209), .Z(n4211) );
  NAND U4710 ( .A(n4212), .B(n4211), .Z(n4330) );
  NANDN U4711 ( .A(n4214), .B(n4213), .Z(n4220) );
  ANDN U4712 ( .B(\stack[1][16] ), .A(n2994), .Z(n4216) );
  NAND U4713 ( .A(n4216), .B(n4215), .Z(n4218) );
  NANDN U4714 ( .A(n2977), .B(o[2]), .Z(n4217) );
  AND U4715 ( .A(n4218), .B(n4217), .Z(n4219) );
  ANDN U4716 ( .B(n4220), .A(n4219), .Z(n4311) );
  AND U4717 ( .A(\stack[1][16] ), .B(o[3]), .Z(n4312) );
  XNOR U4718 ( .A(n4311), .B(n4312), .Z(n4314) );
  IV U4719 ( .A(\stack[1][19] ), .Z(n16746) );
  ANDN U4720 ( .B(o[0]), .A(n16746), .Z(n4222) );
  NANDN U4721 ( .A(n2995), .B(\stack[1][18] ), .Z(n4221) );
  XNOR U4722 ( .A(n4222), .B(n4221), .Z(n4318) );
  AND U4723 ( .A(\stack[1][18] ), .B(o[1]), .Z(n4319) );
  NANDN U4724 ( .A(n2994), .B(n4319), .Z(n4223) );
  XOR U4725 ( .A(n2996), .B(n4223), .Z(n4224) );
  AND U4726 ( .A(n4224), .B(\stack[1][17] ), .Z(n4317) );
  XOR U4727 ( .A(n4318), .B(n4317), .Z(n4313) );
  XOR U4728 ( .A(n4314), .B(n4313), .Z(n4329) );
  XNOR U4729 ( .A(n4330), .B(n4329), .Z(n4332) );
  AND U4730 ( .A(\stack[1][15] ), .B(o[4]), .Z(n4331) );
  XNOR U4731 ( .A(n4332), .B(n4331), .Z(n4307) );
  AND U4732 ( .A(\stack[1][14] ), .B(o[5]), .Z(n4305) );
  OR U4733 ( .A(n4226), .B(n4225), .Z(n4230) );
  NANDN U4734 ( .A(n4228), .B(n4227), .Z(n4229) );
  NAND U4735 ( .A(n4230), .B(n4229), .Z(n4306) );
  XNOR U4736 ( .A(n4305), .B(n4306), .Z(n4308) );
  XNOR U4737 ( .A(n4307), .B(n4308), .Z(n4300) );
  XNOR U4738 ( .A(n4299), .B(n4300), .Z(n4301) );
  AND U4739 ( .A(\stack[1][13] ), .B(o[6]), .Z(n4302) );
  XNOR U4740 ( .A(n4296), .B(n4295), .Z(n4335) );
  XOR U4741 ( .A(n4336), .B(n4335), .Z(n4337) );
  XOR U4742 ( .A(n4338), .B(n4337), .Z(n4290) );
  AND U4743 ( .A(\stack[1][10] ), .B(o[9]), .Z(n4287) );
  OR U4744 ( .A(n4232), .B(n4231), .Z(n4236) );
  OR U4745 ( .A(n4234), .B(n4233), .Z(n4235) );
  NAND U4746 ( .A(n4236), .B(n4235), .Z(n4288) );
  XOR U4747 ( .A(n4287), .B(n4288), .Z(n4289) );
  XNOR U4748 ( .A(n4290), .B(n4289), .Z(n4341) );
  XNOR U4749 ( .A(n4342), .B(n4341), .Z(n4343) );
  XOR U4750 ( .A(n4344), .B(n4343), .Z(n4284) );
  NANDN U4751 ( .A(n4238), .B(n4237), .Z(n4242) );
  OR U4752 ( .A(n4240), .B(n4239), .Z(n4241) );
  AND U4753 ( .A(n4242), .B(n4241), .Z(n4281) );
  AND U4754 ( .A(o[11]), .B(\stack[1][8] ), .Z(n4282) );
  XOR U4755 ( .A(n4281), .B(n4282), .Z(n4283) );
  XNOR U4756 ( .A(n4284), .B(n4283), .Z(n4347) );
  XNOR U4757 ( .A(n4348), .B(n4347), .Z(n4350) );
  NANDN U4758 ( .A(n17219), .B(o[12]), .Z(n4349) );
  XOR U4759 ( .A(n4350), .B(n4349), .Z(n4277) );
  NANDN U4760 ( .A(n4244), .B(n4243), .Z(n4248) );
  OR U4761 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U4762 ( .A(n4248), .B(n4247), .Z(n4275) );
  AND U4763 ( .A(o[13]), .B(\stack[1][6] ), .Z(n4276) );
  XNOR U4764 ( .A(n4275), .B(n4276), .Z(n4278) );
  XOR U4765 ( .A(n4277), .B(n4278), .Z(n4353) );
  XOR U4766 ( .A(n4354), .B(n4353), .Z(n4356) );
  AND U4767 ( .A(o[14]), .B(\stack[1][5] ), .Z(n4355) );
  XNOR U4768 ( .A(n4356), .B(n4355), .Z(n4271) );
  XOR U4769 ( .A(n4360), .B(n4359), .Z(n4362) );
  XNOR U4770 ( .A(n4361), .B(n4362), .Z(n4266) );
  AND U4771 ( .A(o[17]), .B(\stack[1][2] ), .Z(n4263) );
  OR U4772 ( .A(n4250), .B(n4249), .Z(n4254) );
  OR U4773 ( .A(n4252), .B(n4251), .Z(n4253) );
  NAND U4774 ( .A(n4254), .B(n4253), .Z(n4264) );
  XNOR U4775 ( .A(n4263), .B(n4264), .Z(n4265) );
  XOR U4776 ( .A(n4266), .B(n4265), .Z(n4257) );
  XOR U4777 ( .A(n4258), .B(n4257), .Z(n4259) );
  XNOR U4778 ( .A(n4260), .B(n4259), .Z(n16751) );
  OR U4779 ( .A(n16750), .B(n16751), .Z(n4255) );
  AND U4780 ( .A(n4256), .B(n4255), .Z(n4366) );
  AND U4781 ( .A(o[19]), .B(\stack[1][1] ), .Z(n4477) );
  OR U4782 ( .A(n4258), .B(n4257), .Z(n4262) );
  NANDN U4783 ( .A(n4260), .B(n4259), .Z(n4261) );
  NAND U4784 ( .A(n4262), .B(n4261), .Z(n4478) );
  XNOR U4785 ( .A(n4477), .B(n4478), .Z(n4480) );
  OR U4786 ( .A(n4264), .B(n4263), .Z(n4268) );
  OR U4787 ( .A(n4266), .B(n4265), .Z(n4267) );
  AND U4788 ( .A(n4268), .B(n4267), .Z(n4370) );
  OR U4789 ( .A(n4270), .B(n4269), .Z(n4274) );
  OR U4790 ( .A(n4272), .B(n4271), .Z(n4273) );
  NAND U4791 ( .A(n4274), .B(n4273), .Z(n4472) );
  NANDN U4792 ( .A(n17256), .B(o[14]), .Z(n4468) );
  OR U4793 ( .A(n4276), .B(n4275), .Z(n4280) );
  OR U4794 ( .A(n4278), .B(n4277), .Z(n4279) );
  NAND U4795 ( .A(n4280), .B(n4279), .Z(n4466) );
  NANDN U4796 ( .A(n17179), .B(o[12]), .Z(n4462) );
  OR U4797 ( .A(n4282), .B(n4281), .Z(n4286) );
  NANDN U4798 ( .A(n4284), .B(n4283), .Z(n4285) );
  NAND U4799 ( .A(n4286), .B(n4285), .Z(n4460) );
  OR U4800 ( .A(n4288), .B(n4287), .Z(n4292) );
  NANDN U4801 ( .A(n4290), .B(n4289), .Z(n4291) );
  NAND U4802 ( .A(n4292), .B(n4291), .Z(n4400) );
  NANDN U4803 ( .A(n3002), .B(\stack[1][12] ), .Z(n4456) );
  OR U4804 ( .A(n4294), .B(n4293), .Z(n4298) );
  OR U4805 ( .A(n4296), .B(n4295), .Z(n4297) );
  NAND U4806 ( .A(n4298), .B(n4297), .Z(n4454) );
  OR U4807 ( .A(n4300), .B(n4299), .Z(n4304) );
  OR U4808 ( .A(n4302), .B(n4301), .Z(n4303) );
  AND U4809 ( .A(n4304), .B(n4303), .Z(n4411) );
  AND U4810 ( .A(\stack[1][13] ), .B(o[7]), .Z(n4412) );
  XNOR U4811 ( .A(n4411), .B(n4412), .Z(n4414) );
  OR U4812 ( .A(n4306), .B(n4305), .Z(n4310) );
  OR U4813 ( .A(n4308), .B(n4307), .Z(n4309) );
  AND U4814 ( .A(n4310), .B(n4309), .Z(n4417) );
  OR U4815 ( .A(n4312), .B(n4311), .Z(n4316) );
  OR U4816 ( .A(n4314), .B(n4313), .Z(n4315) );
  NAND U4817 ( .A(n4316), .B(n4315), .Z(n4448) );
  NANDN U4818 ( .A(n4318), .B(n4317), .Z(n4324) );
  ANDN U4819 ( .B(\stack[1][17] ), .A(n2994), .Z(n4320) );
  NAND U4820 ( .A(n4320), .B(n4319), .Z(n4322) );
  NANDN U4821 ( .A(n16826), .B(o[2]), .Z(n4321) );
  AND U4822 ( .A(n4322), .B(n4321), .Z(n4323) );
  ANDN U4823 ( .B(n4324), .A(n4323), .Z(n4429) );
  AND U4824 ( .A(\stack[1][17] ), .B(o[3]), .Z(n4430) );
  XNOR U4825 ( .A(n4429), .B(n4430), .Z(n4432) );
  IV U4826 ( .A(\stack[1][20] ), .Z(n16712) );
  ANDN U4827 ( .B(o[0]), .A(n16712), .Z(n4326) );
  NANDN U4828 ( .A(n2995), .B(\stack[1][19] ), .Z(n4325) );
  XNOR U4829 ( .A(n4326), .B(n4325), .Z(n4436) );
  AND U4830 ( .A(\stack[1][19] ), .B(o[1]), .Z(n4437) );
  NANDN U4831 ( .A(n2994), .B(n4437), .Z(n4327) );
  XOR U4832 ( .A(n2996), .B(n4327), .Z(n4328) );
  AND U4833 ( .A(n4328), .B(\stack[1][18] ), .Z(n4435) );
  XOR U4834 ( .A(n4436), .B(n4435), .Z(n4431) );
  XOR U4835 ( .A(n4432), .B(n4431), .Z(n4447) );
  XNOR U4836 ( .A(n4448), .B(n4447), .Z(n4450) );
  AND U4837 ( .A(\stack[1][16] ), .B(o[4]), .Z(n4449) );
  XNOR U4838 ( .A(n4450), .B(n4449), .Z(n4425) );
  AND U4839 ( .A(\stack[1][15] ), .B(o[5]), .Z(n4423) );
  OR U4840 ( .A(n4330), .B(n4329), .Z(n4334) );
  NANDN U4841 ( .A(n4332), .B(n4331), .Z(n4333) );
  NAND U4842 ( .A(n4334), .B(n4333), .Z(n4424) );
  XNOR U4843 ( .A(n4423), .B(n4424), .Z(n4426) );
  XNOR U4844 ( .A(n4425), .B(n4426), .Z(n4418) );
  XOR U4845 ( .A(n4417), .B(n4418), .Z(n4419) );
  AND U4846 ( .A(\stack[1][14] ), .B(o[6]), .Z(n4420) );
  XOR U4847 ( .A(n4419), .B(n4420), .Z(n4413) );
  XOR U4848 ( .A(n4414), .B(n4413), .Z(n4453) );
  XNOR U4849 ( .A(n4454), .B(n4453), .Z(n4455) );
  XNOR U4850 ( .A(n4456), .B(n4455), .Z(n4407) );
  NANDN U4851 ( .A(n2972), .B(o[9]), .Z(n4405) );
  NANDN U4852 ( .A(n4336), .B(n4335), .Z(n4340) );
  OR U4853 ( .A(n4338), .B(n4337), .Z(n4339) );
  NAND U4854 ( .A(n4340), .B(n4339), .Z(n4406) );
  XOR U4855 ( .A(n4405), .B(n4406), .Z(n4408) );
  XNOR U4856 ( .A(n4407), .B(n4408), .Z(n4399) );
  XNOR U4857 ( .A(n4400), .B(n4399), .Z(n4401) );
  NANDN U4858 ( .A(n17101), .B(o[10]), .Z(n4402) );
  AND U4859 ( .A(o[11]), .B(\stack[1][9] ), .Z(n4393) );
  OR U4860 ( .A(n4342), .B(n4341), .Z(n4346) );
  OR U4861 ( .A(n4344), .B(n4343), .Z(n4345) );
  NAND U4862 ( .A(n4346), .B(n4345), .Z(n4394) );
  XOR U4863 ( .A(n4393), .B(n4394), .Z(n4395) );
  XNOR U4864 ( .A(n4396), .B(n4395), .Z(n4459) );
  XNOR U4865 ( .A(n4460), .B(n4459), .Z(n4461) );
  XOR U4866 ( .A(n4462), .B(n4461), .Z(n4390) );
  AND U4867 ( .A(o[13]), .B(\stack[1][7] ), .Z(n4387) );
  OR U4868 ( .A(n4348), .B(n4347), .Z(n4352) );
  OR U4869 ( .A(n4350), .B(n4349), .Z(n4351) );
  NAND U4870 ( .A(n4352), .B(n4351), .Z(n4388) );
  XOR U4871 ( .A(n4387), .B(n4388), .Z(n4389) );
  XNOR U4872 ( .A(n4390), .B(n4389), .Z(n4465) );
  XNOR U4873 ( .A(n4466), .B(n4465), .Z(n4467) );
  XOR U4874 ( .A(n4468), .B(n4467), .Z(n4384) );
  NANDN U4875 ( .A(n4354), .B(n4353), .Z(n4358) );
  OR U4876 ( .A(n4356), .B(n4355), .Z(n4357) );
  AND U4877 ( .A(n4358), .B(n4357), .Z(n4381) );
  AND U4878 ( .A(o[15]), .B(\stack[1][5] ), .Z(n4382) );
  XOR U4879 ( .A(n4381), .B(n4382), .Z(n4383) );
  XNOR U4880 ( .A(n4384), .B(n4383), .Z(n4471) );
  XNOR U4881 ( .A(n4472), .B(n4471), .Z(n4474) );
  NANDN U4882 ( .A(n2971), .B(o[16]), .Z(n4473) );
  XOR U4883 ( .A(n4474), .B(n4473), .Z(n4377) );
  NANDN U4884 ( .A(n4360), .B(n4359), .Z(n4364) );
  OR U4885 ( .A(n4362), .B(n4361), .Z(n4363) );
  AND U4886 ( .A(n4364), .B(n4363), .Z(n4375) );
  AND U4887 ( .A(o[17]), .B(\stack[1][3] ), .Z(n4376) );
  XNOR U4888 ( .A(n4375), .B(n4376), .Z(n4378) );
  XOR U4889 ( .A(n4377), .B(n4378), .Z(n4369) );
  XOR U4890 ( .A(n4370), .B(n4369), .Z(n4372) );
  AND U4891 ( .A(o[18]), .B(\stack[1][2] ), .Z(n4371) );
  XNOR U4892 ( .A(n4372), .B(n4371), .Z(n4479) );
  NANDN U4893 ( .A(n4366), .B(n4365), .Z(n4368) );
  XOR U4894 ( .A(n4366), .B(n4365), .Z(n16709) );
  AND U4895 ( .A(o[20]), .B(\stack[1][0] ), .Z(n16710) );
  OR U4896 ( .A(n16709), .B(n16710), .Z(n4367) );
  AND U4897 ( .A(n4368), .B(n4367), .Z(n4484) );
  OR U4898 ( .A(n4483), .B(n4484), .Z(n4486) );
  NANDN U4899 ( .A(n4370), .B(n4369), .Z(n4374) );
  OR U4900 ( .A(n4372), .B(n4371), .Z(n4373) );
  NAND U4901 ( .A(n4374), .B(n4373), .Z(n4488) );
  ANDN U4902 ( .B(\stack[1][2] ), .A(n3013), .Z(n4487) );
  XOR U4903 ( .A(n4488), .B(n4487), .Z(n4490) );
  NANDN U4904 ( .A(n17375), .B(o[18]), .Z(n4598) );
  OR U4905 ( .A(n4376), .B(n4375), .Z(n4380) );
  OR U4906 ( .A(n4378), .B(n4377), .Z(n4379) );
  NAND U4907 ( .A(n4380), .B(n4379), .Z(n4596) );
  NANDN U4908 ( .A(n17296), .B(o[16]), .Z(n4592) );
  OR U4909 ( .A(n4382), .B(n4381), .Z(n4386) );
  NANDN U4910 ( .A(n4384), .B(n4383), .Z(n4385) );
  NAND U4911 ( .A(n4386), .B(n4385), .Z(n4590) );
  NANDN U4912 ( .A(n17219), .B(o[14]), .Z(n4586) );
  OR U4913 ( .A(n4388), .B(n4387), .Z(n4392) );
  NANDN U4914 ( .A(n4390), .B(n4389), .Z(n4391) );
  NAND U4915 ( .A(n4392), .B(n4391), .Z(n4584) );
  AND U4916 ( .A(o[12]), .B(\stack[1][9] ), .Z(n4513) );
  OR U4917 ( .A(n4394), .B(n4393), .Z(n4398) );
  NANDN U4918 ( .A(n4396), .B(n4395), .Z(n4397) );
  AND U4919 ( .A(n4398), .B(n4397), .Z(n4511) );
  AND U4920 ( .A(o[11]), .B(\stack[1][10] ), .Z(n4577) );
  OR U4921 ( .A(n4400), .B(n4399), .Z(n4404) );
  OR U4922 ( .A(n4402), .B(n4401), .Z(n4403) );
  NAND U4923 ( .A(n4404), .B(n4403), .Z(n4578) );
  XNOR U4924 ( .A(n4577), .B(n4578), .Z(n4580) );
  NANDN U4925 ( .A(n4406), .B(n4405), .Z(n4410) );
  NANDN U4926 ( .A(n4408), .B(n4407), .Z(n4409) );
  AND U4927 ( .A(n4410), .B(n4409), .Z(n4517) );
  OR U4928 ( .A(n4412), .B(n4411), .Z(n4416) );
  OR U4929 ( .A(n4414), .B(n4413), .Z(n4415) );
  NAND U4930 ( .A(n4416), .B(n4415), .Z(n4572) );
  OR U4931 ( .A(n4418), .B(n4417), .Z(n4422) );
  NANDN U4932 ( .A(n4420), .B(n4419), .Z(n4421) );
  AND U4933 ( .A(n4422), .B(n4421), .Z(n4529) );
  AND U4934 ( .A(\stack[1][14] ), .B(o[7]), .Z(n4530) );
  XNOR U4935 ( .A(n4529), .B(n4530), .Z(n4532) );
  OR U4936 ( .A(n4424), .B(n4423), .Z(n4428) );
  OR U4937 ( .A(n4426), .B(n4425), .Z(n4427) );
  AND U4938 ( .A(n4428), .B(n4427), .Z(n4535) );
  OR U4939 ( .A(n4430), .B(n4429), .Z(n4434) );
  OR U4940 ( .A(n4432), .B(n4431), .Z(n4433) );
  NAND U4941 ( .A(n4434), .B(n4433), .Z(n4566) );
  NANDN U4942 ( .A(n4436), .B(n4435), .Z(n4442) );
  ANDN U4943 ( .B(\stack[1][18] ), .A(n2994), .Z(n4438) );
  NAND U4944 ( .A(n4438), .B(n4437), .Z(n4440) );
  NANDN U4945 ( .A(n16786), .B(o[2]), .Z(n4439) );
  AND U4946 ( .A(n4440), .B(n4439), .Z(n4441) );
  ANDN U4947 ( .B(n4442), .A(n4441), .Z(n4547) );
  AND U4948 ( .A(\stack[1][18] ), .B(o[3]), .Z(n4548) );
  XNOR U4949 ( .A(n4547), .B(n4548), .Z(n4550) );
  ANDN U4950 ( .B(o[0]), .A(n2978), .Z(n4444) );
  NANDN U4951 ( .A(n2995), .B(\stack[1][20] ), .Z(n4443) );
  XNOR U4952 ( .A(n4444), .B(n4443), .Z(n4554) );
  AND U4953 ( .A(\stack[1][20] ), .B(o[1]), .Z(n4555) );
  NANDN U4954 ( .A(n2994), .B(n4555), .Z(n4445) );
  XOR U4955 ( .A(n2996), .B(n4445), .Z(n4446) );
  AND U4956 ( .A(n4446), .B(\stack[1][19] ), .Z(n4553) );
  XOR U4957 ( .A(n4554), .B(n4553), .Z(n4549) );
  XOR U4958 ( .A(n4550), .B(n4549), .Z(n4565) );
  XNOR U4959 ( .A(n4566), .B(n4565), .Z(n4568) );
  AND U4960 ( .A(\stack[1][17] ), .B(o[4]), .Z(n4567) );
  XNOR U4961 ( .A(n4568), .B(n4567), .Z(n4543) );
  AND U4962 ( .A(\stack[1][16] ), .B(o[5]), .Z(n4541) );
  OR U4963 ( .A(n4448), .B(n4447), .Z(n4452) );
  NANDN U4964 ( .A(n4450), .B(n4449), .Z(n4451) );
  NAND U4965 ( .A(n4452), .B(n4451), .Z(n4542) );
  XNOR U4966 ( .A(n4541), .B(n4542), .Z(n4544) );
  XNOR U4967 ( .A(n4543), .B(n4544), .Z(n4536) );
  XNOR U4968 ( .A(n4535), .B(n4536), .Z(n4537) );
  AND U4969 ( .A(\stack[1][15] ), .B(o[6]), .Z(n4538) );
  XNOR U4970 ( .A(n4532), .B(n4531), .Z(n4571) );
  XOR U4971 ( .A(n4572), .B(n4571), .Z(n4574) );
  AND U4972 ( .A(\stack[1][13] ), .B(o[8]), .Z(n4573) );
  XNOR U4973 ( .A(n4574), .B(n4573), .Z(n4525) );
  AND U4974 ( .A(\stack[1][12] ), .B(o[9]), .Z(n4523) );
  OR U4975 ( .A(n4454), .B(n4453), .Z(n4458) );
  OR U4976 ( .A(n4456), .B(n4455), .Z(n4457) );
  NAND U4977 ( .A(n4458), .B(n4457), .Z(n4524) );
  XNOR U4978 ( .A(n4523), .B(n4524), .Z(n4526) );
  XNOR U4979 ( .A(n4525), .B(n4526), .Z(n4518) );
  XNOR U4980 ( .A(n4517), .B(n4518), .Z(n4519) );
  AND U4981 ( .A(\stack[1][11] ), .B(o[10]), .Z(n4520) );
  XNOR U4982 ( .A(n4580), .B(n4579), .Z(n4512) );
  XNOR U4983 ( .A(n4511), .B(n4512), .Z(n4514) );
  XNOR U4984 ( .A(n4513), .B(n4514), .Z(n4508) );
  AND U4985 ( .A(o[13]), .B(\stack[1][8] ), .Z(n4505) );
  OR U4986 ( .A(n4460), .B(n4459), .Z(n4464) );
  OR U4987 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U4988 ( .A(n4464), .B(n4463), .Z(n4506) );
  XNOR U4989 ( .A(n4505), .B(n4506), .Z(n4507) );
  XOR U4990 ( .A(n4508), .B(n4507), .Z(n4583) );
  XNOR U4991 ( .A(n4584), .B(n4583), .Z(n4585) );
  AND U4992 ( .A(o[15]), .B(\stack[1][6] ), .Z(n4499) );
  OR U4993 ( .A(n4466), .B(n4465), .Z(n4470) );
  OR U4994 ( .A(n4468), .B(n4467), .Z(n4469) );
  NAND U4995 ( .A(n4470), .B(n4469), .Z(n4500) );
  XOR U4996 ( .A(n4499), .B(n4500), .Z(n4501) );
  XNOR U4997 ( .A(n4502), .B(n4501), .Z(n4589) );
  XNOR U4998 ( .A(n4590), .B(n4589), .Z(n4591) );
  XOR U4999 ( .A(n4592), .B(n4591), .Z(n4496) );
  AND U5000 ( .A(o[17]), .B(\stack[1][4] ), .Z(n4493) );
  OR U5001 ( .A(n4472), .B(n4471), .Z(n4476) );
  OR U5002 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U5003 ( .A(n4476), .B(n4475), .Z(n4494) );
  XOR U5004 ( .A(n4493), .B(n4494), .Z(n4495) );
  XNOR U5005 ( .A(n4496), .B(n4495), .Z(n4595) );
  XNOR U5006 ( .A(n4596), .B(n4595), .Z(n4597) );
  XOR U5007 ( .A(n4598), .B(n4597), .Z(n4489) );
  OR U5008 ( .A(n4478), .B(n4477), .Z(n4482) );
  OR U5009 ( .A(n4480), .B(n4479), .Z(n4481) );
  AND U5010 ( .A(n4482), .B(n4481), .Z(n4602) );
  XNOR U5011 ( .A(n4601), .B(n4602), .Z(n4603) );
  AND U5012 ( .A(o[20]), .B(\stack[1][1] ), .Z(n4604) );
  XOR U5013 ( .A(n4603), .B(n4604), .Z(n16670) );
  XNOR U5014 ( .A(n4484), .B(n4483), .Z(n16669) );
  OR U5015 ( .A(n16670), .B(n16669), .Z(n4485) );
  AND U5016 ( .A(n4486), .B(n4485), .Z(n4608) );
  NANDN U5017 ( .A(n2970), .B(o[20]), .Z(n4735) );
  NANDN U5018 ( .A(n4488), .B(n4487), .Z(n4492) );
  NANDN U5019 ( .A(n4490), .B(n4489), .Z(n4491) );
  AND U5020 ( .A(n4492), .B(n4491), .Z(n4732) );
  NANDN U5021 ( .A(n2971), .B(o[18]), .Z(n4729) );
  OR U5022 ( .A(n4494), .B(n4493), .Z(n4498) );
  NANDN U5023 ( .A(n4496), .B(n4495), .Z(n4497) );
  NAND U5024 ( .A(n4498), .B(n4497), .Z(n4727) );
  NANDN U5025 ( .A(n17256), .B(o[16]), .Z(n4723) );
  OR U5026 ( .A(n4500), .B(n4499), .Z(n4504) );
  NANDN U5027 ( .A(n4502), .B(n4501), .Z(n4503) );
  NAND U5028 ( .A(n4504), .B(n4503), .Z(n4721) );
  AND U5029 ( .A(o[14]), .B(\stack[1][8] ), .Z(n4639) );
  OR U5030 ( .A(n4506), .B(n4505), .Z(n4510) );
  OR U5031 ( .A(n4508), .B(n4507), .Z(n4509) );
  AND U5032 ( .A(n4510), .B(n4509), .Z(n4637) );
  OR U5033 ( .A(n4512), .B(n4511), .Z(n4516) );
  OR U5034 ( .A(n4514), .B(n4513), .Z(n4515) );
  AND U5035 ( .A(n4516), .B(n4515), .Z(n4714) );
  AND U5036 ( .A(o[13]), .B(\stack[1][9] ), .Z(n4715) );
  XNOR U5037 ( .A(n4714), .B(n4715), .Z(n4717) );
  AND U5038 ( .A(\stack[1][11] ), .B(o[11]), .Z(n17061) );
  OR U5039 ( .A(n4518), .B(n4517), .Z(n4522) );
  OR U5040 ( .A(n4520), .B(n4519), .Z(n4521) );
  NAND U5041 ( .A(n4522), .B(n4521), .Z(n4649) );
  XOR U5042 ( .A(n17061), .B(n4649), .Z(n4650) );
  NANDN U5043 ( .A(n3004), .B(\stack[1][12] ), .Z(n4711) );
  OR U5044 ( .A(n4524), .B(n4523), .Z(n4528) );
  OR U5045 ( .A(n4526), .B(n4525), .Z(n4527) );
  NAND U5046 ( .A(n4528), .B(n4527), .Z(n4709) );
  NANDN U5047 ( .A(n3002), .B(\stack[1][14] ), .Z(n4705) );
  OR U5048 ( .A(n4530), .B(n4529), .Z(n4534) );
  OR U5049 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U5050 ( .A(n4534), .B(n4533), .Z(n4703) );
  OR U5051 ( .A(n4536), .B(n4535), .Z(n4540) );
  OR U5052 ( .A(n4538), .B(n4537), .Z(n4539) );
  AND U5053 ( .A(n4540), .B(n4539), .Z(n4660) );
  AND U5054 ( .A(\stack[1][15] ), .B(o[7]), .Z(n4661) );
  XNOR U5055 ( .A(n4660), .B(n4661), .Z(n4663) );
  OR U5056 ( .A(n4542), .B(n4541), .Z(n4546) );
  OR U5057 ( .A(n4544), .B(n4543), .Z(n4545) );
  AND U5058 ( .A(n4546), .B(n4545), .Z(n4666) );
  OR U5059 ( .A(n4548), .B(n4547), .Z(n4552) );
  OR U5060 ( .A(n4550), .B(n4549), .Z(n4551) );
  NAND U5061 ( .A(n4552), .B(n4551), .Z(n4697) );
  NANDN U5062 ( .A(n4554), .B(n4553), .Z(n4560) );
  ANDN U5063 ( .B(\stack[1][19] ), .A(n2994), .Z(n4556) );
  NAND U5064 ( .A(n4556), .B(n4555), .Z(n4558) );
  NANDN U5065 ( .A(n16746), .B(o[2]), .Z(n4557) );
  AND U5066 ( .A(n4558), .B(n4557), .Z(n4559) );
  ANDN U5067 ( .B(n4560), .A(n4559), .Z(n4678) );
  AND U5068 ( .A(\stack[1][19] ), .B(o[3]), .Z(n4679) );
  XNOR U5069 ( .A(n4678), .B(n4679), .Z(n4681) );
  ANDN U5070 ( .B(o[0]), .A(n2979), .Z(n4562) );
  NANDN U5071 ( .A(n2995), .B(\stack[1][21] ), .Z(n4561) );
  XNOR U5072 ( .A(n4562), .B(n4561), .Z(n4685) );
  AND U5073 ( .A(\stack[1][21] ), .B(o[1]), .Z(n4686) );
  NANDN U5074 ( .A(n2994), .B(n4686), .Z(n4563) );
  XOR U5075 ( .A(n2996), .B(n4563), .Z(n4564) );
  AND U5076 ( .A(n4564), .B(\stack[1][20] ), .Z(n4684) );
  XOR U5077 ( .A(n4685), .B(n4684), .Z(n4680) );
  XOR U5078 ( .A(n4681), .B(n4680), .Z(n4696) );
  XNOR U5079 ( .A(n4697), .B(n4696), .Z(n4699) );
  AND U5080 ( .A(\stack[1][18] ), .B(o[4]), .Z(n4698) );
  XNOR U5081 ( .A(n4699), .B(n4698), .Z(n4674) );
  AND U5082 ( .A(\stack[1][17] ), .B(o[5]), .Z(n4672) );
  OR U5083 ( .A(n4566), .B(n4565), .Z(n4570) );
  NANDN U5084 ( .A(n4568), .B(n4567), .Z(n4569) );
  NAND U5085 ( .A(n4570), .B(n4569), .Z(n4673) );
  XNOR U5086 ( .A(n4672), .B(n4673), .Z(n4675) );
  XNOR U5087 ( .A(n4674), .B(n4675), .Z(n4667) );
  XOR U5088 ( .A(n4666), .B(n4667), .Z(n4668) );
  AND U5089 ( .A(\stack[1][16] ), .B(o[6]), .Z(n4669) );
  XOR U5090 ( .A(n4668), .B(n4669), .Z(n4662) );
  XOR U5091 ( .A(n4663), .B(n4662), .Z(n4702) );
  XNOR U5092 ( .A(n4703), .B(n4702), .Z(n4704) );
  XNOR U5093 ( .A(n4705), .B(n4704), .Z(n4656) );
  AND U5094 ( .A(\stack[1][13] ), .B(o[9]), .Z(n4654) );
  NANDN U5095 ( .A(n4572), .B(n4571), .Z(n4576) );
  NANDN U5096 ( .A(n4574), .B(n4573), .Z(n4575) );
  NAND U5097 ( .A(n4576), .B(n4575), .Z(n4655) );
  XNOR U5098 ( .A(n4654), .B(n4655), .Z(n4657) );
  XNOR U5099 ( .A(n4656), .B(n4657), .Z(n4708) );
  XNOR U5100 ( .A(n4709), .B(n4708), .Z(n4710) );
  XNOR U5101 ( .A(n4711), .B(n4710), .Z(n4651) );
  OR U5102 ( .A(n4578), .B(n4577), .Z(n4582) );
  OR U5103 ( .A(n4580), .B(n4579), .Z(n4581) );
  AND U5104 ( .A(n4582), .B(n4581), .Z(n4644) );
  XNOR U5105 ( .A(n4643), .B(n4644), .Z(n4646) );
  AND U5106 ( .A(o[12]), .B(\stack[1][10] ), .Z(n4645) );
  XOR U5107 ( .A(n4646), .B(n4645), .Z(n4716) );
  XOR U5108 ( .A(n4717), .B(n4716), .Z(n4638) );
  XNOR U5109 ( .A(n4637), .B(n4638), .Z(n4640) );
  XNOR U5110 ( .A(n4639), .B(n4640), .Z(n4634) );
  AND U5111 ( .A(o[15]), .B(\stack[1][7] ), .Z(n4631) );
  OR U5112 ( .A(n4584), .B(n4583), .Z(n4588) );
  OR U5113 ( .A(n4586), .B(n4585), .Z(n4587) );
  NAND U5114 ( .A(n4588), .B(n4587), .Z(n4632) );
  XNOR U5115 ( .A(n4631), .B(n4632), .Z(n4633) );
  XOR U5116 ( .A(n4634), .B(n4633), .Z(n4720) );
  XNOR U5117 ( .A(n4721), .B(n4720), .Z(n4722) );
  AND U5118 ( .A(o[17]), .B(\stack[1][5] ), .Z(n4625) );
  OR U5119 ( .A(n4590), .B(n4589), .Z(n4594) );
  OR U5120 ( .A(n4592), .B(n4591), .Z(n4593) );
  NAND U5121 ( .A(n4594), .B(n4593), .Z(n4626) );
  XOR U5122 ( .A(n4625), .B(n4626), .Z(n4627) );
  XNOR U5123 ( .A(n4628), .B(n4627), .Z(n4726) );
  XNOR U5124 ( .A(n4727), .B(n4726), .Z(n4728) );
  XOR U5125 ( .A(n4729), .B(n4728), .Z(n4622) );
  AND U5126 ( .A(o[19]), .B(\stack[1][3] ), .Z(n4619) );
  OR U5127 ( .A(n4596), .B(n4595), .Z(n4600) );
  OR U5128 ( .A(n4598), .B(n4597), .Z(n4599) );
  NAND U5129 ( .A(n4600), .B(n4599), .Z(n4620) );
  XOR U5130 ( .A(n4619), .B(n4620), .Z(n4621) );
  XNOR U5131 ( .A(n4622), .B(n4621), .Z(n4733) );
  XNOR U5132 ( .A(n4732), .B(n4733), .Z(n4734) );
  XOR U5133 ( .A(n4735), .B(n4734), .Z(n4615) );
  NANDN U5134 ( .A(n4602), .B(n4601), .Z(n4606) );
  NANDN U5135 ( .A(n4604), .B(n4603), .Z(n4605) );
  AND U5136 ( .A(n4606), .B(n4605), .Z(n4613) );
  AND U5137 ( .A(o[21]), .B(\stack[1][1] ), .Z(n4614) );
  XNOR U5138 ( .A(n4613), .B(n4614), .Z(n4616) );
  XOR U5139 ( .A(n4615), .B(n4616), .Z(n4607) );
  NANDN U5140 ( .A(n4608), .B(n4607), .Z(n4610) );
  XOR U5141 ( .A(n4608), .B(n4607), .Z(n16630) );
  AND U5142 ( .A(o[22]), .B(\stack[1][0] ), .Z(n16631) );
  OR U5143 ( .A(n16630), .B(n16631), .Z(n4609) );
  AND U5144 ( .A(n4610), .B(n4609), .Z(n4612) );
  OR U5145 ( .A(n4611), .B(n4612), .Z(n4739) );
  XNOR U5146 ( .A(n4612), .B(n4611), .Z(n16592) );
  NANDN U5147 ( .A(n2969), .B(o[22]), .Z(n4869) );
  OR U5148 ( .A(n4614), .B(n4613), .Z(n4618) );
  OR U5149 ( .A(n4616), .B(n4615), .Z(n4617) );
  NAND U5150 ( .A(n4618), .B(n4617), .Z(n4867) );
  NANDN U5151 ( .A(n17375), .B(o[20]), .Z(n4863) );
  OR U5152 ( .A(n4620), .B(n4619), .Z(n4624) );
  NANDN U5153 ( .A(n4622), .B(n4621), .Z(n4623) );
  NAND U5154 ( .A(n4624), .B(n4623), .Z(n4861) );
  NANDN U5155 ( .A(n17296), .B(o[18]), .Z(n4857) );
  OR U5156 ( .A(n4626), .B(n4625), .Z(n4630) );
  NANDN U5157 ( .A(n4628), .B(n4627), .Z(n4629) );
  NAND U5158 ( .A(n4630), .B(n4629), .Z(n4855) );
  AND U5159 ( .A(o[16]), .B(\stack[1][7] ), .Z(n4760) );
  OR U5160 ( .A(n4632), .B(n4631), .Z(n4636) );
  OR U5161 ( .A(n4634), .B(n4633), .Z(n4635) );
  AND U5162 ( .A(n4636), .B(n4635), .Z(n4758) );
  OR U5163 ( .A(n4638), .B(n4637), .Z(n4642) );
  OR U5164 ( .A(n4640), .B(n4639), .Z(n4641) );
  AND U5165 ( .A(n4642), .B(n4641), .Z(n4848) );
  AND U5166 ( .A(o[15]), .B(\stack[1][8] ), .Z(n4849) );
  XNOR U5167 ( .A(n4848), .B(n4849), .Z(n4851) );
  OR U5168 ( .A(n4644), .B(n4643), .Z(n4648) );
  OR U5169 ( .A(n4646), .B(n4645), .Z(n4647) );
  NAND U5170 ( .A(n4648), .B(n4647), .Z(n4771) );
  ANDN U5171 ( .B(\stack[1][10] ), .A(n3007), .Z(n4770) );
  XNOR U5172 ( .A(n4771), .B(n4770), .Z(n4772) );
  NANDN U5173 ( .A(n2972), .B(o[12]), .Z(n4845) );
  NANDN U5174 ( .A(n4649), .B(n17061), .Z(n4653) );
  OR U5175 ( .A(n4651), .B(n4650), .Z(n4652) );
  AND U5176 ( .A(n4653), .B(n4652), .Z(n4842) );
  NANDN U5177 ( .A(n3004), .B(\stack[1][13] ), .Z(n4785) );
  OR U5178 ( .A(n4655), .B(n4654), .Z(n4659) );
  NANDN U5179 ( .A(n4657), .B(n4656), .Z(n4658) );
  NAND U5180 ( .A(n4659), .B(n4658), .Z(n4783) );
  NANDN U5181 ( .A(n3002), .B(\stack[1][15] ), .Z(n4839) );
  OR U5182 ( .A(n4661), .B(n4660), .Z(n4665) );
  OR U5183 ( .A(n4663), .B(n4662), .Z(n4664) );
  NAND U5184 ( .A(n4665), .B(n4664), .Z(n4837) );
  OR U5185 ( .A(n4667), .B(n4666), .Z(n4671) );
  NANDN U5186 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U5187 ( .A(n4671), .B(n4670), .Z(n4794) );
  AND U5188 ( .A(\stack[1][16] ), .B(o[7]), .Z(n4795) );
  XNOR U5189 ( .A(n4794), .B(n4795), .Z(n4797) );
  OR U5190 ( .A(n4673), .B(n4672), .Z(n4677) );
  OR U5191 ( .A(n4675), .B(n4674), .Z(n4676) );
  AND U5192 ( .A(n4677), .B(n4676), .Z(n4800) );
  OR U5193 ( .A(n4679), .B(n4678), .Z(n4683) );
  OR U5194 ( .A(n4681), .B(n4680), .Z(n4682) );
  NAND U5195 ( .A(n4683), .B(n4682), .Z(n4831) );
  NANDN U5196 ( .A(n4685), .B(n4684), .Z(n4691) );
  ANDN U5197 ( .B(\stack[1][20] ), .A(n2994), .Z(n4687) );
  NAND U5198 ( .A(n4687), .B(n4686), .Z(n4689) );
  NANDN U5199 ( .A(n16712), .B(o[2]), .Z(n4688) );
  AND U5200 ( .A(n4689), .B(n4688), .Z(n4690) );
  ANDN U5201 ( .B(n4691), .A(n4690), .Z(n4812) );
  AND U5202 ( .A(\stack[1][20] ), .B(o[3]), .Z(n4813) );
  XNOR U5203 ( .A(n4812), .B(n4813), .Z(n4815) );
  ANDN U5204 ( .B(o[0]), .A(n2980), .Z(n4693) );
  NANDN U5205 ( .A(n2995), .B(\stack[1][22] ), .Z(n4692) );
  XNOR U5206 ( .A(n4693), .B(n4692), .Z(n4819) );
  AND U5207 ( .A(\stack[1][22] ), .B(o[1]), .Z(n4820) );
  NANDN U5208 ( .A(n2994), .B(n4820), .Z(n4694) );
  XOR U5209 ( .A(n2996), .B(n4694), .Z(n4695) );
  AND U5210 ( .A(n4695), .B(\stack[1][21] ), .Z(n4818) );
  XOR U5211 ( .A(n4819), .B(n4818), .Z(n4814) );
  XOR U5212 ( .A(n4815), .B(n4814), .Z(n4830) );
  XNOR U5213 ( .A(n4831), .B(n4830), .Z(n4833) );
  AND U5214 ( .A(\stack[1][19] ), .B(o[4]), .Z(n4832) );
  XNOR U5215 ( .A(n4833), .B(n4832), .Z(n4808) );
  AND U5216 ( .A(\stack[1][18] ), .B(o[5]), .Z(n4806) );
  OR U5217 ( .A(n4697), .B(n4696), .Z(n4701) );
  NANDN U5218 ( .A(n4699), .B(n4698), .Z(n4700) );
  NAND U5219 ( .A(n4701), .B(n4700), .Z(n4807) );
  XNOR U5220 ( .A(n4806), .B(n4807), .Z(n4809) );
  XNOR U5221 ( .A(n4808), .B(n4809), .Z(n4801) );
  XOR U5222 ( .A(n4800), .B(n4801), .Z(n4802) );
  AND U5223 ( .A(\stack[1][17] ), .B(o[6]), .Z(n4803) );
  XOR U5224 ( .A(n4802), .B(n4803), .Z(n4796) );
  XOR U5225 ( .A(n4797), .B(n4796), .Z(n4836) );
  XNOR U5226 ( .A(n4837), .B(n4836), .Z(n4838) );
  XNOR U5227 ( .A(n4839), .B(n4838), .Z(n4790) );
  NANDN U5228 ( .A(n2975), .B(o[9]), .Z(n4788) );
  OR U5229 ( .A(n4703), .B(n4702), .Z(n4707) );
  OR U5230 ( .A(n4705), .B(n4704), .Z(n4706) );
  NAND U5231 ( .A(n4707), .B(n4706), .Z(n4789) );
  XOR U5232 ( .A(n4788), .B(n4789), .Z(n4791) );
  XNOR U5233 ( .A(n4790), .B(n4791), .Z(n4782) );
  XNOR U5234 ( .A(n4783), .B(n4782), .Z(n4784) );
  XNOR U5235 ( .A(n4785), .B(n4784), .Z(n4778) );
  NANDN U5236 ( .A(n2973), .B(o[11]), .Z(n4776) );
  OR U5237 ( .A(n4709), .B(n4708), .Z(n4713) );
  OR U5238 ( .A(n4711), .B(n4710), .Z(n4712) );
  NAND U5239 ( .A(n4713), .B(n4712), .Z(n4777) );
  XOR U5240 ( .A(n4776), .B(n4777), .Z(n4779) );
  XNOR U5241 ( .A(n4778), .B(n4779), .Z(n4843) );
  XNOR U5242 ( .A(n4842), .B(n4843), .Z(n4844) );
  XOR U5243 ( .A(n4772), .B(n4773), .Z(n4764) );
  OR U5244 ( .A(n4715), .B(n4714), .Z(n4719) );
  NANDN U5245 ( .A(n4717), .B(n4716), .Z(n4718) );
  AND U5246 ( .A(n4719), .B(n4718), .Z(n4765) );
  XOR U5247 ( .A(n4764), .B(n4765), .Z(n4767) );
  AND U5248 ( .A(o[14]), .B(\stack[1][9] ), .Z(n4766) );
  XOR U5249 ( .A(n4767), .B(n4766), .Z(n4850) );
  XOR U5250 ( .A(n4851), .B(n4850), .Z(n4759) );
  XNOR U5251 ( .A(n4758), .B(n4759), .Z(n4761) );
  XNOR U5252 ( .A(n4760), .B(n4761), .Z(n4755) );
  AND U5253 ( .A(o[17]), .B(\stack[1][6] ), .Z(n4752) );
  OR U5254 ( .A(n4721), .B(n4720), .Z(n4725) );
  OR U5255 ( .A(n4723), .B(n4722), .Z(n4724) );
  NAND U5256 ( .A(n4725), .B(n4724), .Z(n4753) );
  XNOR U5257 ( .A(n4752), .B(n4753), .Z(n4754) );
  XOR U5258 ( .A(n4755), .B(n4754), .Z(n4854) );
  XNOR U5259 ( .A(n4855), .B(n4854), .Z(n4856) );
  AND U5260 ( .A(o[19]), .B(\stack[1][4] ), .Z(n4746) );
  OR U5261 ( .A(n4727), .B(n4726), .Z(n4731) );
  OR U5262 ( .A(n4729), .B(n4728), .Z(n4730) );
  NAND U5263 ( .A(n4731), .B(n4730), .Z(n4747) );
  XOR U5264 ( .A(n4746), .B(n4747), .Z(n4748) );
  XNOR U5265 ( .A(n4749), .B(n4748), .Z(n4860) );
  XNOR U5266 ( .A(n4861), .B(n4860), .Z(n4862) );
  XOR U5267 ( .A(n4863), .B(n4862), .Z(n4743) );
  AND U5268 ( .A(o[21]), .B(\stack[1][2] ), .Z(n4740) );
  OR U5269 ( .A(n4733), .B(n4732), .Z(n4737) );
  OR U5270 ( .A(n4735), .B(n4734), .Z(n4736) );
  NAND U5271 ( .A(n4737), .B(n4736), .Z(n4741) );
  XOR U5272 ( .A(n4740), .B(n4741), .Z(n4742) );
  XNOR U5273 ( .A(n4743), .B(n4742), .Z(n4866) );
  XNOR U5274 ( .A(n4867), .B(n4866), .Z(n4868) );
  XOR U5275 ( .A(n4869), .B(n4868), .Z(n16593) );
  OR U5276 ( .A(n16592), .B(n16593), .Z(n4738) );
  AND U5277 ( .A(n4739), .B(n4738), .Z(n4873) );
  NANDN U5278 ( .A(n2970), .B(o[22]), .Z(n5012) );
  OR U5279 ( .A(n4741), .B(n4740), .Z(n4745) );
  NANDN U5280 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U5281 ( .A(n4745), .B(n4744), .Z(n5010) );
  NANDN U5282 ( .A(n2971), .B(o[20]), .Z(n5006) );
  OR U5283 ( .A(n4747), .B(n4746), .Z(n4751) );
  NANDN U5284 ( .A(n4749), .B(n4748), .Z(n4750) );
  NAND U5285 ( .A(n4751), .B(n4750), .Z(n5004) );
  AND U5286 ( .A(o[18]), .B(\stack[1][6] ), .Z(n4898) );
  OR U5287 ( .A(n4753), .B(n4752), .Z(n4757) );
  OR U5288 ( .A(n4755), .B(n4754), .Z(n4756) );
  AND U5289 ( .A(n4757), .B(n4756), .Z(n4896) );
  OR U5290 ( .A(n4759), .B(n4758), .Z(n4763) );
  OR U5291 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U5292 ( .A(n4763), .B(n4762), .Z(n4997) );
  AND U5293 ( .A(o[17]), .B(\stack[1][7] ), .Z(n4998) );
  XNOR U5294 ( .A(n4997), .B(n4998), .Z(n5000) );
  NANDN U5295 ( .A(n4765), .B(n4764), .Z(n4769) );
  OR U5296 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U5297 ( .A(n4769), .B(n4768), .Z(n4909) );
  ANDN U5298 ( .B(\stack[1][9] ), .A(n3009), .Z(n4908) );
  XNOR U5299 ( .A(n4909), .B(n4908), .Z(n4910) );
  NANDN U5300 ( .A(n17101), .B(o[14]), .Z(n4994) );
  NANDN U5301 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U5302 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U5303 ( .A(n4775), .B(n4774), .Z(n4991) );
  AND U5304 ( .A(o[12]), .B(\stack[1][12] ), .Z(n17027) );
  NANDN U5305 ( .A(n4777), .B(n4776), .Z(n4781) );
  NANDN U5306 ( .A(n4779), .B(n4778), .Z(n4780) );
  AND U5307 ( .A(n4781), .B(n4780), .Z(n4986) );
  AND U5308 ( .A(\stack[1][13] ), .B(o[11]), .Z(n4920) );
  OR U5309 ( .A(n4783), .B(n4782), .Z(n4787) );
  OR U5310 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U5311 ( .A(n4787), .B(n4786), .Z(n4921) );
  XNOR U5312 ( .A(n4920), .B(n4921), .Z(n4923) );
  NANDN U5313 ( .A(n4789), .B(n4788), .Z(n4793) );
  NANDN U5314 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U5315 ( .A(n4793), .B(n4792), .Z(n4926) );
  OR U5316 ( .A(n4795), .B(n4794), .Z(n4799) );
  OR U5317 ( .A(n4797), .B(n4796), .Z(n4798) );
  NAND U5318 ( .A(n4799), .B(n4798), .Z(n4981) );
  OR U5319 ( .A(n4801), .B(n4800), .Z(n4805) );
  NANDN U5320 ( .A(n4803), .B(n4802), .Z(n4804) );
  AND U5321 ( .A(n4805), .B(n4804), .Z(n4938) );
  AND U5322 ( .A(\stack[1][17] ), .B(o[7]), .Z(n4939) );
  XNOR U5323 ( .A(n4938), .B(n4939), .Z(n4941) );
  OR U5324 ( .A(n4807), .B(n4806), .Z(n4811) );
  OR U5325 ( .A(n4809), .B(n4808), .Z(n4810) );
  AND U5326 ( .A(n4811), .B(n4810), .Z(n4944) );
  OR U5327 ( .A(n4813), .B(n4812), .Z(n4817) );
  OR U5328 ( .A(n4815), .B(n4814), .Z(n4816) );
  NAND U5329 ( .A(n4817), .B(n4816), .Z(n4975) );
  NANDN U5330 ( .A(n4819), .B(n4818), .Z(n4825) );
  ANDN U5331 ( .B(\stack[1][21] ), .A(n2994), .Z(n4821) );
  NAND U5332 ( .A(n4821), .B(n4820), .Z(n4823) );
  NANDN U5333 ( .A(n2978), .B(o[2]), .Z(n4822) );
  AND U5334 ( .A(n4823), .B(n4822), .Z(n4824) );
  ANDN U5335 ( .B(n4825), .A(n4824), .Z(n4956) );
  AND U5336 ( .A(\stack[1][21] ), .B(o[3]), .Z(n4957) );
  XNOR U5337 ( .A(n4956), .B(n4957), .Z(n4959) );
  ANDN U5338 ( .B(o[0]), .A(n2981), .Z(n4827) );
  NANDN U5339 ( .A(n2995), .B(\stack[1][23] ), .Z(n4826) );
  XNOR U5340 ( .A(n4827), .B(n4826), .Z(n4963) );
  AND U5341 ( .A(\stack[1][23] ), .B(o[1]), .Z(n4964) );
  NANDN U5342 ( .A(n2994), .B(n4964), .Z(n4828) );
  XOR U5343 ( .A(n2996), .B(n4828), .Z(n4829) );
  AND U5344 ( .A(n4829), .B(\stack[1][22] ), .Z(n4962) );
  XOR U5345 ( .A(n4963), .B(n4962), .Z(n4958) );
  XOR U5346 ( .A(n4959), .B(n4958), .Z(n4974) );
  XNOR U5347 ( .A(n4975), .B(n4974), .Z(n4977) );
  AND U5348 ( .A(\stack[1][20] ), .B(o[4]), .Z(n4976) );
  XNOR U5349 ( .A(n4977), .B(n4976), .Z(n4952) );
  AND U5350 ( .A(\stack[1][19] ), .B(o[5]), .Z(n4950) );
  OR U5351 ( .A(n4831), .B(n4830), .Z(n4835) );
  NANDN U5352 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U5353 ( .A(n4835), .B(n4834), .Z(n4951) );
  XNOR U5354 ( .A(n4950), .B(n4951), .Z(n4953) );
  XNOR U5355 ( .A(n4952), .B(n4953), .Z(n4945) );
  XNOR U5356 ( .A(n4944), .B(n4945), .Z(n4946) );
  AND U5357 ( .A(\stack[1][18] ), .B(o[6]), .Z(n4947) );
  XNOR U5358 ( .A(n4941), .B(n4940), .Z(n4980) );
  XOR U5359 ( .A(n4981), .B(n4980), .Z(n4983) );
  AND U5360 ( .A(\stack[1][16] ), .B(o[8]), .Z(n4982) );
  XNOR U5361 ( .A(n4983), .B(n4982), .Z(n4934) );
  AND U5362 ( .A(\stack[1][15] ), .B(o[9]), .Z(n4932) );
  OR U5363 ( .A(n4837), .B(n4836), .Z(n4841) );
  OR U5364 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U5365 ( .A(n4841), .B(n4840), .Z(n4933) );
  XNOR U5366 ( .A(n4932), .B(n4933), .Z(n4935) );
  XNOR U5367 ( .A(n4934), .B(n4935), .Z(n4927) );
  XNOR U5368 ( .A(n4926), .B(n4927), .Z(n4928) );
  AND U5369 ( .A(\stack[1][14] ), .B(o[10]), .Z(n4929) );
  XNOR U5370 ( .A(n4923), .B(n4922), .Z(n4987) );
  XOR U5371 ( .A(n4986), .B(n4987), .Z(n4988) );
  XOR U5372 ( .A(n17027), .B(n4988), .Z(n4917) );
  AND U5373 ( .A(o[13]), .B(\stack[1][11] ), .Z(n4914) );
  OR U5374 ( .A(n4843), .B(n4842), .Z(n4847) );
  OR U5375 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5376 ( .A(n4847), .B(n4846), .Z(n4915) );
  XNOR U5377 ( .A(n4914), .B(n4915), .Z(n4916) );
  XOR U5378 ( .A(n4917), .B(n4916), .Z(n4992) );
  XNOR U5379 ( .A(n4991), .B(n4992), .Z(n4993) );
  XOR U5380 ( .A(n4910), .B(n4911), .Z(n4902) );
  OR U5381 ( .A(n4849), .B(n4848), .Z(n4853) );
  NANDN U5382 ( .A(n4851), .B(n4850), .Z(n4852) );
  AND U5383 ( .A(n4853), .B(n4852), .Z(n4903) );
  XOR U5384 ( .A(n4902), .B(n4903), .Z(n4905) );
  AND U5385 ( .A(o[16]), .B(\stack[1][8] ), .Z(n4904) );
  XOR U5386 ( .A(n4905), .B(n4904), .Z(n4999) );
  XOR U5387 ( .A(n5000), .B(n4999), .Z(n4897) );
  XNOR U5388 ( .A(n4896), .B(n4897), .Z(n4899) );
  XNOR U5389 ( .A(n4898), .B(n4899), .Z(n4893) );
  AND U5390 ( .A(o[19]), .B(\stack[1][5] ), .Z(n4890) );
  OR U5391 ( .A(n4855), .B(n4854), .Z(n4859) );
  OR U5392 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U5393 ( .A(n4859), .B(n4858), .Z(n4891) );
  XNOR U5394 ( .A(n4890), .B(n4891), .Z(n4892) );
  XOR U5395 ( .A(n4893), .B(n4892), .Z(n5003) );
  XNOR U5396 ( .A(n5004), .B(n5003), .Z(n5005) );
  AND U5397 ( .A(o[21]), .B(\stack[1][3] ), .Z(n4884) );
  OR U5398 ( .A(n4861), .B(n4860), .Z(n4865) );
  OR U5399 ( .A(n4863), .B(n4862), .Z(n4864) );
  NAND U5400 ( .A(n4865), .B(n4864), .Z(n4885) );
  XOR U5401 ( .A(n4884), .B(n4885), .Z(n4886) );
  XNOR U5402 ( .A(n4887), .B(n4886), .Z(n5009) );
  XNOR U5403 ( .A(n5010), .B(n5009), .Z(n5011) );
  XOR U5404 ( .A(n5012), .B(n5011), .Z(n4880) );
  AND U5405 ( .A(o[23]), .B(\stack[1][1] ), .Z(n4878) );
  OR U5406 ( .A(n4867), .B(n4866), .Z(n4871) );
  OR U5407 ( .A(n4869), .B(n4868), .Z(n4870) );
  NAND U5408 ( .A(n4871), .B(n4870), .Z(n4879) );
  XNOR U5409 ( .A(n4878), .B(n4879), .Z(n4881) );
  XOR U5410 ( .A(n4880), .B(n4881), .Z(n4872) );
  NANDN U5411 ( .A(n4873), .B(n4872), .Z(n4875) );
  XOR U5412 ( .A(n4873), .B(n4872), .Z(n16552) );
  AND U5413 ( .A(o[24]), .B(\stack[1][0] ), .Z(n16553) );
  OR U5414 ( .A(n16552), .B(n16553), .Z(n4874) );
  AND U5415 ( .A(n4875), .B(n4874), .Z(n4877) );
  OR U5416 ( .A(n4876), .B(n4877), .Z(n5016) );
  XNOR U5417 ( .A(n4877), .B(n4876), .Z(n16511) );
  NANDN U5418 ( .A(n2969), .B(o[24]), .Z(n5158) );
  OR U5419 ( .A(n4879), .B(n4878), .Z(n4883) );
  OR U5420 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U5421 ( .A(n4883), .B(n4882), .Z(n5156) );
  NANDN U5422 ( .A(n17375), .B(o[22]), .Z(n5026) );
  OR U5423 ( .A(n4885), .B(n4884), .Z(n4889) );
  NANDN U5424 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U5425 ( .A(n4889), .B(n4888), .Z(n5024) );
  AND U5426 ( .A(o[20]), .B(\stack[1][5] ), .Z(n5151) );
  OR U5427 ( .A(n4891), .B(n4890), .Z(n4895) );
  OR U5428 ( .A(n4893), .B(n4892), .Z(n4894) );
  AND U5429 ( .A(n4895), .B(n4894), .Z(n5150) );
  OR U5430 ( .A(n4897), .B(n4896), .Z(n4901) );
  OR U5431 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U5432 ( .A(n4901), .B(n4900), .Z(n5035) );
  AND U5433 ( .A(o[19]), .B(\stack[1][6] ), .Z(n5036) );
  XNOR U5434 ( .A(n5035), .B(n5036), .Z(n5038) );
  NANDN U5435 ( .A(n4903), .B(n4902), .Z(n4907) );
  OR U5436 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U5437 ( .A(n4907), .B(n4906), .Z(n5042) );
  ANDN U5438 ( .B(\stack[1][8] ), .A(n3011), .Z(n5041) );
  XNOR U5439 ( .A(n5042), .B(n5041), .Z(n5043) );
  NANDN U5440 ( .A(n17145), .B(o[16]), .Z(n5140) );
  NANDN U5441 ( .A(n4909), .B(n4908), .Z(n4913) );
  NANDN U5442 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U5443 ( .A(n4913), .B(n4912), .Z(n5137) );
  NANDN U5444 ( .A(n2972), .B(o[14]), .Z(n5134) );
  OR U5445 ( .A(n4915), .B(n4914), .Z(n4919) );
  OR U5446 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U5447 ( .A(n4919), .B(n4918), .Z(n5132) );
  NANDN U5448 ( .A(n3006), .B(\stack[1][13] ), .Z(n5062) );
  OR U5449 ( .A(n4921), .B(n4920), .Z(n4925) );
  OR U5450 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U5451 ( .A(n4925), .B(n4924), .Z(n5060) );
  OR U5452 ( .A(n4927), .B(n4926), .Z(n4931) );
  OR U5453 ( .A(n4929), .B(n4928), .Z(n4930) );
  AND U5454 ( .A(n4931), .B(n4930), .Z(n5125) );
  AND U5455 ( .A(\stack[1][14] ), .B(o[11]), .Z(n5126) );
  XNOR U5456 ( .A(n5125), .B(n5126), .Z(n5128) );
  OR U5457 ( .A(n4933), .B(n4932), .Z(n4937) );
  OR U5458 ( .A(n4935), .B(n4934), .Z(n4936) );
  AND U5459 ( .A(n4937), .B(n4936), .Z(n5065) );
  OR U5460 ( .A(n4939), .B(n4938), .Z(n4943) );
  OR U5461 ( .A(n4941), .B(n4940), .Z(n4942) );
  NAND U5462 ( .A(n4943), .B(n4942), .Z(n5120) );
  OR U5463 ( .A(n4945), .B(n4944), .Z(n4949) );
  OR U5464 ( .A(n4947), .B(n4946), .Z(n4948) );
  AND U5465 ( .A(n4949), .B(n4948), .Z(n5077) );
  AND U5466 ( .A(\stack[1][18] ), .B(o[7]), .Z(n5078) );
  XNOR U5467 ( .A(n5077), .B(n5078), .Z(n5080) );
  OR U5468 ( .A(n4951), .B(n4950), .Z(n4955) );
  OR U5469 ( .A(n4953), .B(n4952), .Z(n4954) );
  AND U5470 ( .A(n4955), .B(n4954), .Z(n5083) );
  OR U5471 ( .A(n4957), .B(n4956), .Z(n4961) );
  OR U5472 ( .A(n4959), .B(n4958), .Z(n4960) );
  NAND U5473 ( .A(n4961), .B(n4960), .Z(n5114) );
  NANDN U5474 ( .A(n4963), .B(n4962), .Z(n4969) );
  ANDN U5475 ( .B(\stack[1][22] ), .A(n2994), .Z(n4965) );
  NAND U5476 ( .A(n4965), .B(n4964), .Z(n4967) );
  NANDN U5477 ( .A(n2979), .B(o[2]), .Z(n4966) );
  AND U5478 ( .A(n4967), .B(n4966), .Z(n4968) );
  ANDN U5479 ( .B(n4969), .A(n4968), .Z(n5095) );
  AND U5480 ( .A(\stack[1][22] ), .B(o[3]), .Z(n5096) );
  XNOR U5481 ( .A(n5095), .B(n5096), .Z(n5098) );
  ANDN U5482 ( .B(o[0]), .A(n2982), .Z(n4971) );
  NANDN U5483 ( .A(n2995), .B(\stack[1][24] ), .Z(n4970) );
  XNOR U5484 ( .A(n4971), .B(n4970), .Z(n5102) );
  AND U5485 ( .A(\stack[1][24] ), .B(o[1]), .Z(n5103) );
  NANDN U5486 ( .A(n2994), .B(n5103), .Z(n4972) );
  XOR U5487 ( .A(n2996), .B(n4972), .Z(n4973) );
  AND U5488 ( .A(n4973), .B(\stack[1][23] ), .Z(n5101) );
  XOR U5489 ( .A(n5102), .B(n5101), .Z(n5097) );
  XOR U5490 ( .A(n5098), .B(n5097), .Z(n5113) );
  XNOR U5491 ( .A(n5114), .B(n5113), .Z(n5116) );
  AND U5492 ( .A(\stack[1][21] ), .B(o[4]), .Z(n5115) );
  XNOR U5493 ( .A(n5116), .B(n5115), .Z(n5091) );
  AND U5494 ( .A(\stack[1][20] ), .B(o[5]), .Z(n5089) );
  OR U5495 ( .A(n4975), .B(n4974), .Z(n4979) );
  NANDN U5496 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5497 ( .A(n4979), .B(n4978), .Z(n5090) );
  XNOR U5498 ( .A(n5089), .B(n5090), .Z(n5092) );
  XNOR U5499 ( .A(n5091), .B(n5092), .Z(n5084) );
  XNOR U5500 ( .A(n5083), .B(n5084), .Z(n5085) );
  AND U5501 ( .A(\stack[1][19] ), .B(o[6]), .Z(n5086) );
  XNOR U5502 ( .A(n5080), .B(n5079), .Z(n5119) );
  XOR U5503 ( .A(n5120), .B(n5119), .Z(n5122) );
  AND U5504 ( .A(\stack[1][17] ), .B(o[8]), .Z(n5121) );
  XNOR U5505 ( .A(n5122), .B(n5121), .Z(n5073) );
  AND U5506 ( .A(\stack[1][16] ), .B(o[9]), .Z(n5071) );
  NANDN U5507 ( .A(n4981), .B(n4980), .Z(n4985) );
  NANDN U5508 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5509 ( .A(n4985), .B(n4984), .Z(n5072) );
  XNOR U5510 ( .A(n5071), .B(n5072), .Z(n5074) );
  XNOR U5511 ( .A(n5073), .B(n5074), .Z(n5066) );
  XOR U5512 ( .A(n5065), .B(n5066), .Z(n5067) );
  AND U5513 ( .A(\stack[1][15] ), .B(o[10]), .Z(n5068) );
  XOR U5514 ( .A(n5067), .B(n5068), .Z(n5127) );
  XOR U5515 ( .A(n5128), .B(n5127), .Z(n5059) );
  XNOR U5516 ( .A(n5060), .B(n5059), .Z(n5061) );
  XNOR U5517 ( .A(n5062), .B(n5061), .Z(n5055) );
  OR U5518 ( .A(n4987), .B(n4986), .Z(n4990) );
  NANDN U5519 ( .A(n17027), .B(n4988), .Z(n4989) );
  AND U5520 ( .A(n4990), .B(n4989), .Z(n5054) );
  NANDN U5521 ( .A(n3007), .B(\stack[1][12] ), .Z(n5053) );
  XOR U5522 ( .A(n5054), .B(n5053), .Z(n5056) );
  XNOR U5523 ( .A(n5055), .B(n5056), .Z(n5131) );
  XNOR U5524 ( .A(n5132), .B(n5131), .Z(n5133) );
  XNOR U5525 ( .A(n5134), .B(n5133), .Z(n5049) );
  NANDN U5526 ( .A(n3009), .B(\stack[1][10] ), .Z(n5047) );
  OR U5527 ( .A(n4992), .B(n4991), .Z(n4996) );
  OR U5528 ( .A(n4994), .B(n4993), .Z(n4995) );
  NAND U5529 ( .A(n4996), .B(n4995), .Z(n5048) );
  XOR U5530 ( .A(n5047), .B(n5048), .Z(n5050) );
  XNOR U5531 ( .A(n5049), .B(n5050), .Z(n5138) );
  XNOR U5532 ( .A(n5137), .B(n5138), .Z(n5139) );
  XOR U5533 ( .A(n5043), .B(n5044), .Z(n5143) );
  OR U5534 ( .A(n4998), .B(n4997), .Z(n5002) );
  NANDN U5535 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U5536 ( .A(n5002), .B(n5001), .Z(n5144) );
  XOR U5537 ( .A(n5143), .B(n5144), .Z(n5146) );
  AND U5538 ( .A(o[18]), .B(\stack[1][7] ), .Z(n5145) );
  XNOR U5539 ( .A(n5146), .B(n5145), .Z(n5037) );
  XOR U5540 ( .A(n5150), .B(n5149), .Z(n5152) );
  XNOR U5541 ( .A(n5151), .B(n5152), .Z(n5032) );
  AND U5542 ( .A(o[21]), .B(\stack[1][4] ), .Z(n5029) );
  OR U5543 ( .A(n5004), .B(n5003), .Z(n5008) );
  OR U5544 ( .A(n5006), .B(n5005), .Z(n5007) );
  NAND U5545 ( .A(n5008), .B(n5007), .Z(n5030) );
  XNOR U5546 ( .A(n5029), .B(n5030), .Z(n5031) );
  XOR U5547 ( .A(n5032), .B(n5031), .Z(n5023) );
  XNOR U5548 ( .A(n5024), .B(n5023), .Z(n5025) );
  AND U5549 ( .A(o[23]), .B(\stack[1][2] ), .Z(n5017) );
  OR U5550 ( .A(n5010), .B(n5009), .Z(n5014) );
  OR U5551 ( .A(n5012), .B(n5011), .Z(n5013) );
  NAND U5552 ( .A(n5014), .B(n5013), .Z(n5018) );
  XOR U5553 ( .A(n5017), .B(n5018), .Z(n5019) );
  XNOR U5554 ( .A(n5020), .B(n5019), .Z(n5155) );
  XNOR U5555 ( .A(n5156), .B(n5155), .Z(n5157) );
  XOR U5556 ( .A(n5158), .B(n5157), .Z(n16512) );
  OR U5557 ( .A(n16511), .B(n16512), .Z(n5015) );
  AND U5558 ( .A(n5016), .B(n5015), .Z(n5162) );
  AND U5559 ( .A(o[24]), .B(\stack[1][2] ), .Z(n5173) );
  OR U5560 ( .A(n5018), .B(n5017), .Z(n5022) );
  NANDN U5561 ( .A(n5020), .B(n5019), .Z(n5021) );
  AND U5562 ( .A(n5022), .B(n5021), .Z(n5172) );
  AND U5563 ( .A(o[23]), .B(\stack[1][3] ), .Z(n5308) );
  OR U5564 ( .A(n5024), .B(n5023), .Z(n5028) );
  OR U5565 ( .A(n5026), .B(n5025), .Z(n5027) );
  NAND U5566 ( .A(n5028), .B(n5027), .Z(n5309) );
  XNOR U5567 ( .A(n5308), .B(n5309), .Z(n5311) );
  OR U5568 ( .A(n5030), .B(n5029), .Z(n5034) );
  OR U5569 ( .A(n5032), .B(n5031), .Z(n5033) );
  AND U5570 ( .A(n5034), .B(n5033), .Z(n5177) );
  OR U5571 ( .A(n5036), .B(n5035), .Z(n5040) );
  OR U5572 ( .A(n5038), .B(n5037), .Z(n5039) );
  NAND U5573 ( .A(n5040), .B(n5039), .Z(n5303) );
  NANDN U5574 ( .A(n17179), .B(o[18]), .Z(n5299) );
  NANDN U5575 ( .A(n5042), .B(n5041), .Z(n5046) );
  NANDN U5576 ( .A(n5044), .B(n5043), .Z(n5045) );
  AND U5577 ( .A(n5046), .B(n5045), .Z(n5296) );
  NANDN U5578 ( .A(n17101), .B(o[16]), .Z(n5293) );
  NANDN U5579 ( .A(n5048), .B(n5047), .Z(n5052) );
  NANDN U5580 ( .A(n5050), .B(n5049), .Z(n5051) );
  NAND U5581 ( .A(n5052), .B(n5051), .Z(n5291) );
  NANDN U5582 ( .A(n2973), .B(o[14]), .Z(n5210) );
  NANDN U5583 ( .A(n5054), .B(n5053), .Z(n5058) );
  NANDN U5584 ( .A(n5056), .B(n5055), .Z(n5057) );
  NAND U5585 ( .A(n5058), .B(n5057), .Z(n5208) );
  AND U5586 ( .A(\stack[1][13] ), .B(o[13]), .Z(n16983) );
  OR U5587 ( .A(n5060), .B(n5059), .Z(n5064) );
  OR U5588 ( .A(n5062), .B(n5061), .Z(n5063) );
  NAND U5589 ( .A(n5064), .B(n5063), .Z(n5285) );
  XNOR U5590 ( .A(n16983), .B(n5285), .Z(n5287) );
  OR U5591 ( .A(n5066), .B(n5065), .Z(n5070) );
  NANDN U5592 ( .A(n5068), .B(n5067), .Z(n5069) );
  NAND U5593 ( .A(n5070), .B(n5069), .Z(n5220) );
  ANDN U5594 ( .B(o[11]), .A(n2976), .Z(n5219) );
  XOR U5595 ( .A(n5220), .B(n5219), .Z(n5221) );
  NANDN U5596 ( .A(n3004), .B(\stack[1][16] ), .Z(n5282) );
  OR U5597 ( .A(n5072), .B(n5071), .Z(n5076) );
  OR U5598 ( .A(n5074), .B(n5073), .Z(n5075) );
  NAND U5599 ( .A(n5076), .B(n5075), .Z(n5280) );
  NANDN U5600 ( .A(n3002), .B(\stack[1][18] ), .Z(n5276) );
  OR U5601 ( .A(n5078), .B(n5077), .Z(n5082) );
  OR U5602 ( .A(n5080), .B(n5079), .Z(n5081) );
  NAND U5603 ( .A(n5082), .B(n5081), .Z(n5274) );
  OR U5604 ( .A(n5084), .B(n5083), .Z(n5088) );
  OR U5605 ( .A(n5086), .B(n5085), .Z(n5087) );
  AND U5606 ( .A(n5088), .B(n5087), .Z(n5231) );
  AND U5607 ( .A(\stack[1][19] ), .B(o[7]), .Z(n5232) );
  XNOR U5608 ( .A(n5231), .B(n5232), .Z(n5234) );
  OR U5609 ( .A(n5090), .B(n5089), .Z(n5094) );
  OR U5610 ( .A(n5092), .B(n5091), .Z(n5093) );
  AND U5611 ( .A(n5094), .B(n5093), .Z(n5237) );
  OR U5612 ( .A(n5096), .B(n5095), .Z(n5100) );
  OR U5613 ( .A(n5098), .B(n5097), .Z(n5099) );
  NAND U5614 ( .A(n5100), .B(n5099), .Z(n5268) );
  NANDN U5615 ( .A(n5102), .B(n5101), .Z(n5108) );
  ANDN U5616 ( .B(\stack[1][23] ), .A(n2994), .Z(n5104) );
  NAND U5617 ( .A(n5104), .B(n5103), .Z(n5106) );
  NANDN U5618 ( .A(n2980), .B(o[2]), .Z(n5105) );
  AND U5619 ( .A(n5106), .B(n5105), .Z(n5107) );
  ANDN U5620 ( .B(n5108), .A(n5107), .Z(n5249) );
  AND U5621 ( .A(\stack[1][23] ), .B(o[3]), .Z(n5250) );
  XNOR U5622 ( .A(n5249), .B(n5250), .Z(n5252) );
  ANDN U5623 ( .B(o[0]), .A(n2983), .Z(n5110) );
  NANDN U5624 ( .A(n2995), .B(\stack[1][25] ), .Z(n5109) );
  XNOR U5625 ( .A(n5110), .B(n5109), .Z(n5256) );
  AND U5626 ( .A(\stack[1][25] ), .B(o[1]), .Z(n5257) );
  NANDN U5627 ( .A(n2994), .B(n5257), .Z(n5111) );
  XOR U5628 ( .A(n2996), .B(n5111), .Z(n5112) );
  AND U5629 ( .A(n5112), .B(\stack[1][24] ), .Z(n5255) );
  XOR U5630 ( .A(n5256), .B(n5255), .Z(n5251) );
  XOR U5631 ( .A(n5252), .B(n5251), .Z(n5267) );
  XNOR U5632 ( .A(n5268), .B(n5267), .Z(n5270) );
  AND U5633 ( .A(\stack[1][22] ), .B(o[4]), .Z(n5269) );
  XNOR U5634 ( .A(n5270), .B(n5269), .Z(n5245) );
  AND U5635 ( .A(\stack[1][21] ), .B(o[5]), .Z(n5243) );
  OR U5636 ( .A(n5114), .B(n5113), .Z(n5118) );
  NANDN U5637 ( .A(n5116), .B(n5115), .Z(n5117) );
  NAND U5638 ( .A(n5118), .B(n5117), .Z(n5244) );
  XNOR U5639 ( .A(n5243), .B(n5244), .Z(n5246) );
  XNOR U5640 ( .A(n5245), .B(n5246), .Z(n5238) );
  XOR U5641 ( .A(n5237), .B(n5238), .Z(n5239) );
  AND U5642 ( .A(\stack[1][20] ), .B(o[6]), .Z(n5240) );
  XOR U5643 ( .A(n5239), .B(n5240), .Z(n5233) );
  XOR U5644 ( .A(n5234), .B(n5233), .Z(n5273) );
  XNOR U5645 ( .A(n5274), .B(n5273), .Z(n5275) );
  XNOR U5646 ( .A(n5276), .B(n5275), .Z(n5227) );
  AND U5647 ( .A(\stack[1][17] ), .B(o[9]), .Z(n5225) );
  NANDN U5648 ( .A(n5120), .B(n5119), .Z(n5124) );
  NANDN U5649 ( .A(n5122), .B(n5121), .Z(n5123) );
  NAND U5650 ( .A(n5124), .B(n5123), .Z(n5226) );
  XNOR U5651 ( .A(n5225), .B(n5226), .Z(n5228) );
  XNOR U5652 ( .A(n5227), .B(n5228), .Z(n5279) );
  XNOR U5653 ( .A(n5280), .B(n5279), .Z(n5281) );
  XNOR U5654 ( .A(n5282), .B(n5281), .Z(n5222) );
  OR U5655 ( .A(n5126), .B(n5125), .Z(n5130) );
  OR U5656 ( .A(n5128), .B(n5127), .Z(n5129) );
  AND U5657 ( .A(n5130), .B(n5129), .Z(n5214) );
  XNOR U5658 ( .A(n5213), .B(n5214), .Z(n5216) );
  AND U5659 ( .A(\stack[1][14] ), .B(o[12]), .Z(n5215) );
  XNOR U5660 ( .A(n5216), .B(n5215), .Z(n5286) );
  XOR U5661 ( .A(n5287), .B(n5286), .Z(n5207) );
  XNOR U5662 ( .A(n5208), .B(n5207), .Z(n5209) );
  XNOR U5663 ( .A(n5210), .B(n5209), .Z(n5203) );
  NANDN U5664 ( .A(n3009), .B(\stack[1][11] ), .Z(n5201) );
  OR U5665 ( .A(n5132), .B(n5131), .Z(n5136) );
  OR U5666 ( .A(n5134), .B(n5133), .Z(n5135) );
  NAND U5667 ( .A(n5136), .B(n5135), .Z(n5202) );
  XOR U5668 ( .A(n5201), .B(n5202), .Z(n5204) );
  XNOR U5669 ( .A(n5203), .B(n5204), .Z(n5290) );
  XNOR U5670 ( .A(n5291), .B(n5290), .Z(n5292) );
  XOR U5671 ( .A(n5293), .B(n5292), .Z(n5197) );
  AND U5672 ( .A(o[17]), .B(\stack[1][9] ), .Z(n5195) );
  OR U5673 ( .A(n5138), .B(n5137), .Z(n5142) );
  OR U5674 ( .A(n5140), .B(n5139), .Z(n5141) );
  NAND U5675 ( .A(n5142), .B(n5141), .Z(n5196) );
  XNOR U5676 ( .A(n5195), .B(n5196), .Z(n5198) );
  XNOR U5677 ( .A(n5296), .B(n5297), .Z(n5298) );
  XOR U5678 ( .A(n5299), .B(n5298), .Z(n5191) );
  NANDN U5679 ( .A(n5144), .B(n5143), .Z(n5148) );
  OR U5680 ( .A(n5146), .B(n5145), .Z(n5147) );
  AND U5681 ( .A(n5148), .B(n5147), .Z(n5189) );
  AND U5682 ( .A(o[19]), .B(\stack[1][7] ), .Z(n5190) );
  XNOR U5683 ( .A(n5189), .B(n5190), .Z(n5192) );
  XOR U5684 ( .A(n5303), .B(n5302), .Z(n5305) );
  AND U5685 ( .A(o[20]), .B(\stack[1][6] ), .Z(n5304) );
  XNOR U5686 ( .A(n5305), .B(n5304), .Z(n5185) );
  NANDN U5687 ( .A(n5150), .B(n5149), .Z(n5154) );
  OR U5688 ( .A(n5152), .B(n5151), .Z(n5153) );
  AND U5689 ( .A(n5154), .B(n5153), .Z(n5183) );
  AND U5690 ( .A(o[21]), .B(\stack[1][5] ), .Z(n5184) );
  XNOR U5691 ( .A(n5183), .B(n5184), .Z(n5186) );
  XNOR U5692 ( .A(n5185), .B(n5186), .Z(n5178) );
  XNOR U5693 ( .A(n5177), .B(n5178), .Z(n5180) );
  AND U5694 ( .A(o[22]), .B(\stack[1][4] ), .Z(n5179) );
  XNOR U5695 ( .A(n5180), .B(n5179), .Z(n5310) );
  XOR U5696 ( .A(n5172), .B(n5171), .Z(n5174) );
  XNOR U5697 ( .A(n5173), .B(n5174), .Z(n5168) );
  AND U5698 ( .A(o[25]), .B(\stack[1][1] ), .Z(n5165) );
  OR U5699 ( .A(n5156), .B(n5155), .Z(n5160) );
  OR U5700 ( .A(n5158), .B(n5157), .Z(n5159) );
  NAND U5701 ( .A(n5160), .B(n5159), .Z(n5166) );
  XNOR U5702 ( .A(n5165), .B(n5166), .Z(n5167) );
  NANDN U5703 ( .A(n5162), .B(n5161), .Z(n5164) );
  XOR U5704 ( .A(n5162), .B(n5161), .Z(n16475) );
  AND U5705 ( .A(o[26]), .B(\stack[1][0] ), .Z(n16476) );
  OR U5706 ( .A(n16475), .B(n16476), .Z(n5163) );
  AND U5707 ( .A(n5164), .B(n5163), .Z(n5315) );
  OR U5708 ( .A(n5314), .B(n5315), .Z(n5317) );
  AND U5709 ( .A(o[26]), .B(\stack[1][1] ), .Z(n5320) );
  OR U5710 ( .A(n5166), .B(n5165), .Z(n5170) );
  OR U5711 ( .A(n5168), .B(n5167), .Z(n5169) );
  AND U5712 ( .A(n5170), .B(n5169), .Z(n5319) );
  NANDN U5713 ( .A(n5172), .B(n5171), .Z(n5176) );
  OR U5714 ( .A(n5174), .B(n5173), .Z(n5175) );
  AND U5715 ( .A(n5176), .B(n5175), .Z(n5468) );
  AND U5716 ( .A(o[25]), .B(\stack[1][2] ), .Z(n5469) );
  XNOR U5717 ( .A(n5468), .B(n5469), .Z(n5471) );
  OR U5718 ( .A(n5178), .B(n5177), .Z(n5182) );
  OR U5719 ( .A(n5180), .B(n5179), .Z(n5181) );
  NAND U5720 ( .A(n5182), .B(n5181), .Z(n5331) );
  ANDN U5721 ( .B(\stack[1][4] ), .A(n3017), .Z(n5330) );
  XOR U5722 ( .A(n5331), .B(n5330), .Z(n5332) );
  NANDN U5723 ( .A(n17296), .B(o[22]), .Z(n5465) );
  OR U5724 ( .A(n5184), .B(n5183), .Z(n5188) );
  OR U5725 ( .A(n5186), .B(n5185), .Z(n5187) );
  NAND U5726 ( .A(n5188), .B(n5187), .Z(n5463) );
  NANDN U5727 ( .A(n17219), .B(o[20]), .Z(n5459) );
  OR U5728 ( .A(n5190), .B(n5189), .Z(n5194) );
  OR U5729 ( .A(n5192), .B(n5191), .Z(n5193) );
  NAND U5730 ( .A(n5194), .B(n5193), .Z(n5457) );
  NANDN U5731 ( .A(n17145), .B(o[18]), .Z(n5453) );
  OR U5732 ( .A(n5196), .B(n5195), .Z(n5200) );
  OR U5733 ( .A(n5198), .B(n5197), .Z(n5199) );
  NAND U5734 ( .A(n5200), .B(n5199), .Z(n5451) );
  AND U5735 ( .A(o[16]), .B(\stack[1][11] ), .Z(n5447) );
  NANDN U5736 ( .A(n5202), .B(n5201), .Z(n5206) );
  NANDN U5737 ( .A(n5204), .B(n5203), .Z(n5205) );
  AND U5738 ( .A(n5206), .B(n5205), .Z(n5444) );
  AND U5739 ( .A(o[15]), .B(\stack[1][12] ), .Z(n5354) );
  OR U5740 ( .A(n5208), .B(n5207), .Z(n5212) );
  OR U5741 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U5742 ( .A(n5212), .B(n5211), .Z(n5355) );
  XNOR U5743 ( .A(n5354), .B(n5355), .Z(n5357) );
  OR U5744 ( .A(n5214), .B(n5213), .Z(n5218) );
  OR U5745 ( .A(n5216), .B(n5215), .Z(n5217) );
  NAND U5746 ( .A(n5218), .B(n5217), .Z(n5361) );
  ANDN U5747 ( .B(o[13]), .A(n2975), .Z(n5360) );
  XNOR U5748 ( .A(n5361), .B(n5360), .Z(n5362) );
  NANDN U5749 ( .A(n3006), .B(\stack[1][15] ), .Z(n5435) );
  NANDN U5750 ( .A(n5220), .B(n5219), .Z(n5224) );
  OR U5751 ( .A(n5222), .B(n5221), .Z(n5223) );
  AND U5752 ( .A(n5224), .B(n5223), .Z(n5432) );
  NANDN U5753 ( .A(n3004), .B(\stack[1][17] ), .Z(n5429) );
  OR U5754 ( .A(n5226), .B(n5225), .Z(n5230) );
  NANDN U5755 ( .A(n5228), .B(n5227), .Z(n5229) );
  NAND U5756 ( .A(n5230), .B(n5229), .Z(n5427) );
  NANDN U5757 ( .A(n3002), .B(\stack[1][19] ), .Z(n5423) );
  OR U5758 ( .A(n5232), .B(n5231), .Z(n5236) );
  OR U5759 ( .A(n5234), .B(n5233), .Z(n5235) );
  NAND U5760 ( .A(n5236), .B(n5235), .Z(n5421) );
  OR U5761 ( .A(n5238), .B(n5237), .Z(n5242) );
  NANDN U5762 ( .A(n5240), .B(n5239), .Z(n5241) );
  AND U5763 ( .A(n5242), .B(n5241), .Z(n5378) );
  AND U5764 ( .A(\stack[1][20] ), .B(o[7]), .Z(n5379) );
  XNOR U5765 ( .A(n5378), .B(n5379), .Z(n5381) );
  OR U5766 ( .A(n5244), .B(n5243), .Z(n5248) );
  OR U5767 ( .A(n5246), .B(n5245), .Z(n5247) );
  AND U5768 ( .A(n5248), .B(n5247), .Z(n5384) );
  OR U5769 ( .A(n5250), .B(n5249), .Z(n5254) );
  OR U5770 ( .A(n5252), .B(n5251), .Z(n5253) );
  NAND U5771 ( .A(n5254), .B(n5253), .Z(n5415) );
  NANDN U5772 ( .A(n5256), .B(n5255), .Z(n5262) );
  ANDN U5773 ( .B(\stack[1][24] ), .A(n2994), .Z(n5258) );
  NAND U5774 ( .A(n5258), .B(n5257), .Z(n5260) );
  NANDN U5775 ( .A(n2981), .B(o[2]), .Z(n5259) );
  AND U5776 ( .A(n5260), .B(n5259), .Z(n5261) );
  ANDN U5777 ( .B(n5262), .A(n5261), .Z(n5396) );
  AND U5778 ( .A(\stack[1][24] ), .B(o[3]), .Z(n5397) );
  XNOR U5779 ( .A(n5396), .B(n5397), .Z(n5399) );
  ANDN U5780 ( .B(o[0]), .A(n2984), .Z(n5264) );
  NANDN U5781 ( .A(n2995), .B(\stack[1][26] ), .Z(n5263) );
  XNOR U5782 ( .A(n5264), .B(n5263), .Z(n5403) );
  AND U5783 ( .A(\stack[1][26] ), .B(o[1]), .Z(n5404) );
  NANDN U5784 ( .A(n2994), .B(n5404), .Z(n5265) );
  XOR U5785 ( .A(n2996), .B(n5265), .Z(n5266) );
  AND U5786 ( .A(n5266), .B(\stack[1][25] ), .Z(n5402) );
  XOR U5787 ( .A(n5403), .B(n5402), .Z(n5398) );
  XOR U5788 ( .A(n5399), .B(n5398), .Z(n5414) );
  XNOR U5789 ( .A(n5415), .B(n5414), .Z(n5417) );
  AND U5790 ( .A(\stack[1][23] ), .B(o[4]), .Z(n5416) );
  XNOR U5791 ( .A(n5417), .B(n5416), .Z(n5392) );
  AND U5792 ( .A(\stack[1][22] ), .B(o[5]), .Z(n5390) );
  OR U5793 ( .A(n5268), .B(n5267), .Z(n5272) );
  NANDN U5794 ( .A(n5270), .B(n5269), .Z(n5271) );
  NAND U5795 ( .A(n5272), .B(n5271), .Z(n5391) );
  XNOR U5796 ( .A(n5390), .B(n5391), .Z(n5393) );
  XNOR U5797 ( .A(n5392), .B(n5393), .Z(n5385) );
  XOR U5798 ( .A(n5384), .B(n5385), .Z(n5386) );
  AND U5799 ( .A(\stack[1][21] ), .B(o[6]), .Z(n5387) );
  XOR U5800 ( .A(n5386), .B(n5387), .Z(n5380) );
  XOR U5801 ( .A(n5381), .B(n5380), .Z(n5420) );
  XNOR U5802 ( .A(n5421), .B(n5420), .Z(n5422) );
  XNOR U5803 ( .A(n5423), .B(n5422), .Z(n5374) );
  NANDN U5804 ( .A(n16786), .B(o[9]), .Z(n5372) );
  OR U5805 ( .A(n5274), .B(n5273), .Z(n5278) );
  OR U5806 ( .A(n5276), .B(n5275), .Z(n5277) );
  NAND U5807 ( .A(n5278), .B(n5277), .Z(n5373) );
  XOR U5808 ( .A(n5372), .B(n5373), .Z(n5375) );
  XNOR U5809 ( .A(n5374), .B(n5375), .Z(n5426) );
  XNOR U5810 ( .A(n5427), .B(n5426), .Z(n5428) );
  XNOR U5811 ( .A(n5429), .B(n5428), .Z(n5368) );
  NANDN U5812 ( .A(n2977), .B(o[11]), .Z(n5366) );
  OR U5813 ( .A(n5280), .B(n5279), .Z(n5284) );
  OR U5814 ( .A(n5282), .B(n5281), .Z(n5283) );
  NAND U5815 ( .A(n5284), .B(n5283), .Z(n5367) );
  XOR U5816 ( .A(n5366), .B(n5367), .Z(n5369) );
  XNOR U5817 ( .A(n5368), .B(n5369), .Z(n5433) );
  XNOR U5818 ( .A(n5432), .B(n5433), .Z(n5434) );
  XOR U5819 ( .A(n5362), .B(n5363), .Z(n5438) );
  OR U5820 ( .A(n5285), .B(n16983), .Z(n5289) );
  OR U5821 ( .A(n5287), .B(n5286), .Z(n5288) );
  AND U5822 ( .A(n5289), .B(n5288), .Z(n5439) );
  XOR U5823 ( .A(n5438), .B(n5439), .Z(n5441) );
  AND U5824 ( .A(o[14]), .B(\stack[1][13] ), .Z(n5440) );
  XOR U5825 ( .A(n5441), .B(n5440), .Z(n5356) );
  XOR U5826 ( .A(n5357), .B(n5356), .Z(n5445) );
  XOR U5827 ( .A(n5444), .B(n5445), .Z(n5446) );
  XOR U5828 ( .A(n5447), .B(n5446), .Z(n5351) );
  AND U5829 ( .A(o[17]), .B(\stack[1][10] ), .Z(n5348) );
  OR U5830 ( .A(n5291), .B(n5290), .Z(n5295) );
  OR U5831 ( .A(n5293), .B(n5292), .Z(n5294) );
  NAND U5832 ( .A(n5295), .B(n5294), .Z(n5349) );
  XNOR U5833 ( .A(n5348), .B(n5349), .Z(n5350) );
  XOR U5834 ( .A(n5351), .B(n5350), .Z(n5450) );
  XNOR U5835 ( .A(n5451), .B(n5450), .Z(n5452) );
  XNOR U5836 ( .A(n5453), .B(n5452), .Z(n5344) );
  NANDN U5837 ( .A(n3013), .B(\stack[1][8] ), .Z(n5342) );
  OR U5838 ( .A(n5297), .B(n5296), .Z(n5301) );
  OR U5839 ( .A(n5299), .B(n5298), .Z(n5300) );
  NAND U5840 ( .A(n5301), .B(n5300), .Z(n5343) );
  XOR U5841 ( .A(n5342), .B(n5343), .Z(n5345) );
  XNOR U5842 ( .A(n5344), .B(n5345), .Z(n5456) );
  XNOR U5843 ( .A(n5457), .B(n5456), .Z(n5458) );
  XNOR U5844 ( .A(n5459), .B(n5458), .Z(n5338) );
  NANDN U5845 ( .A(n3015), .B(\stack[1][6] ), .Z(n5336) );
  NANDN U5846 ( .A(n5303), .B(n5302), .Z(n5307) );
  NANDN U5847 ( .A(n5305), .B(n5304), .Z(n5306) );
  NAND U5848 ( .A(n5307), .B(n5306), .Z(n5337) );
  XOR U5849 ( .A(n5336), .B(n5337), .Z(n5339) );
  XNOR U5850 ( .A(n5338), .B(n5339), .Z(n5462) );
  XNOR U5851 ( .A(n5463), .B(n5462), .Z(n5464) );
  XNOR U5852 ( .A(n5465), .B(n5464), .Z(n5333) );
  OR U5853 ( .A(n5309), .B(n5308), .Z(n5313) );
  OR U5854 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5855 ( .A(n5313), .B(n5312), .Z(n5325) );
  XNOR U5856 ( .A(n5324), .B(n5325), .Z(n5326) );
  AND U5857 ( .A(o[24]), .B(\stack[1][3] ), .Z(n5327) );
  XOR U5858 ( .A(n5471), .B(n5470), .Z(n5318) );
  XOR U5859 ( .A(n5319), .B(n5318), .Z(n5321) );
  XNOR U5860 ( .A(n5320), .B(n5321), .Z(n16437) );
  XNOR U5861 ( .A(n5315), .B(n5314), .Z(n16438) );
  OR U5862 ( .A(n16437), .B(n16438), .Z(n5316) );
  AND U5863 ( .A(n5317), .B(n5316), .Z(n5475) );
  NANDN U5864 ( .A(n5319), .B(n5318), .Z(n5323) );
  OR U5865 ( .A(n5321), .B(n5320), .Z(n5322) );
  AND U5866 ( .A(n5323), .B(n5322), .Z(n5634) );
  AND U5867 ( .A(o[27]), .B(\stack[1][1] ), .Z(n5635) );
  XNOR U5868 ( .A(n5634), .B(n5635), .Z(n5637) );
  OR U5869 ( .A(n5325), .B(n5324), .Z(n5329) );
  OR U5870 ( .A(n5327), .B(n5326), .Z(n5328) );
  NAND U5871 ( .A(n5329), .B(n5328), .Z(n5485) );
  ANDN U5872 ( .B(\stack[1][3] ), .A(n3019), .Z(n5484) );
  XOR U5873 ( .A(n5485), .B(n5484), .Z(n5486) );
  NANDN U5874 ( .A(n2971), .B(o[24]), .Z(n5631) );
  NANDN U5875 ( .A(n5331), .B(n5330), .Z(n5335) );
  OR U5876 ( .A(n5333), .B(n5332), .Z(n5334) );
  AND U5877 ( .A(n5335), .B(n5334), .Z(n5628) );
  NANDN U5878 ( .A(n17256), .B(o[22]), .Z(n5625) );
  NANDN U5879 ( .A(n5337), .B(n5336), .Z(n5341) );
  NANDN U5880 ( .A(n5339), .B(n5338), .Z(n5340) );
  NAND U5881 ( .A(n5341), .B(n5340), .Z(n5623) );
  NANDN U5882 ( .A(n17179), .B(o[20]), .Z(n5619) );
  NANDN U5883 ( .A(n5343), .B(n5342), .Z(n5347) );
  NANDN U5884 ( .A(n5345), .B(n5344), .Z(n5346) );
  NAND U5885 ( .A(n5347), .B(n5346), .Z(n5617) );
  NANDN U5886 ( .A(n17101), .B(o[18]), .Z(n5613) );
  OR U5887 ( .A(n5349), .B(n5348), .Z(n5353) );
  OR U5888 ( .A(n5351), .B(n5350), .Z(n5352) );
  NAND U5889 ( .A(n5353), .B(n5352), .Z(n5611) );
  NANDN U5890 ( .A(n2973), .B(o[16]), .Z(n5607) );
  OR U5891 ( .A(n5355), .B(n5354), .Z(n5359) );
  NANDN U5892 ( .A(n5357), .B(n5356), .Z(n5358) );
  NAND U5893 ( .A(n5359), .B(n5358), .Z(n5605) );
  NOR U5894 ( .A(n3008), .B(n2975), .Z(n5600) );
  NANDN U5895 ( .A(n5361), .B(n5360), .Z(n5365) );
  NANDN U5896 ( .A(n5363), .B(n5362), .Z(n5364) );
  AND U5897 ( .A(n5365), .B(n5364), .Z(n5598) );
  NANDN U5898 ( .A(n3006), .B(\stack[1][16] ), .Z(n5595) );
  NANDN U5899 ( .A(n5367), .B(n5366), .Z(n5371) );
  NANDN U5900 ( .A(n5369), .B(n5368), .Z(n5370) );
  NAND U5901 ( .A(n5371), .B(n5370), .Z(n5593) );
  NANDN U5902 ( .A(n3004), .B(\stack[1][18] ), .Z(n5589) );
  NANDN U5903 ( .A(n5373), .B(n5372), .Z(n5377) );
  NANDN U5904 ( .A(n5375), .B(n5374), .Z(n5376) );
  NAND U5905 ( .A(n5377), .B(n5376), .Z(n5587) );
  NANDN U5906 ( .A(n3002), .B(\stack[1][20] ), .Z(n5583) );
  OR U5907 ( .A(n5379), .B(n5378), .Z(n5383) );
  OR U5908 ( .A(n5381), .B(n5380), .Z(n5382) );
  NAND U5909 ( .A(n5383), .B(n5382), .Z(n5581) );
  OR U5910 ( .A(n5385), .B(n5384), .Z(n5389) );
  NANDN U5911 ( .A(n5387), .B(n5386), .Z(n5388) );
  AND U5912 ( .A(n5389), .B(n5388), .Z(n5538) );
  AND U5913 ( .A(\stack[1][21] ), .B(o[7]), .Z(n5539) );
  XNOR U5914 ( .A(n5538), .B(n5539), .Z(n5541) );
  OR U5915 ( .A(n5391), .B(n5390), .Z(n5395) );
  OR U5916 ( .A(n5393), .B(n5392), .Z(n5394) );
  AND U5917 ( .A(n5395), .B(n5394), .Z(n5544) );
  OR U5918 ( .A(n5397), .B(n5396), .Z(n5401) );
  OR U5919 ( .A(n5399), .B(n5398), .Z(n5400) );
  NAND U5920 ( .A(n5401), .B(n5400), .Z(n5575) );
  NANDN U5921 ( .A(n5403), .B(n5402), .Z(n5409) );
  ANDN U5922 ( .B(\stack[1][25] ), .A(n2994), .Z(n5405) );
  NAND U5923 ( .A(n5405), .B(n5404), .Z(n5407) );
  NANDN U5924 ( .A(n2982), .B(o[2]), .Z(n5406) );
  AND U5925 ( .A(n5407), .B(n5406), .Z(n5408) );
  ANDN U5926 ( .B(n5409), .A(n5408), .Z(n5556) );
  AND U5927 ( .A(\stack[1][25] ), .B(o[3]), .Z(n5557) );
  XNOR U5928 ( .A(n5556), .B(n5557), .Z(n5559) );
  ANDN U5929 ( .B(o[0]), .A(n2985), .Z(n5411) );
  NANDN U5930 ( .A(n2995), .B(\stack[1][27] ), .Z(n5410) );
  XNOR U5931 ( .A(n5411), .B(n5410), .Z(n5563) );
  AND U5932 ( .A(\stack[1][27] ), .B(o[1]), .Z(n5564) );
  NANDN U5933 ( .A(n2994), .B(n5564), .Z(n5412) );
  XOR U5934 ( .A(n2996), .B(n5412), .Z(n5413) );
  AND U5935 ( .A(n5413), .B(\stack[1][26] ), .Z(n5562) );
  XOR U5936 ( .A(n5563), .B(n5562), .Z(n5558) );
  XOR U5937 ( .A(n5559), .B(n5558), .Z(n5574) );
  XNOR U5938 ( .A(n5575), .B(n5574), .Z(n5577) );
  AND U5939 ( .A(\stack[1][24] ), .B(o[4]), .Z(n5576) );
  XNOR U5940 ( .A(n5577), .B(n5576), .Z(n5552) );
  AND U5941 ( .A(\stack[1][23] ), .B(o[5]), .Z(n5550) );
  OR U5942 ( .A(n5415), .B(n5414), .Z(n5419) );
  NANDN U5943 ( .A(n5417), .B(n5416), .Z(n5418) );
  NAND U5944 ( .A(n5419), .B(n5418), .Z(n5551) );
  XNOR U5945 ( .A(n5550), .B(n5551), .Z(n5553) );
  XNOR U5946 ( .A(n5552), .B(n5553), .Z(n5545) );
  XOR U5947 ( .A(n5544), .B(n5545), .Z(n5546) );
  AND U5948 ( .A(\stack[1][22] ), .B(o[6]), .Z(n5547) );
  XOR U5949 ( .A(n5546), .B(n5547), .Z(n5540) );
  XOR U5950 ( .A(n5541), .B(n5540), .Z(n5580) );
  XNOR U5951 ( .A(n5581), .B(n5580), .Z(n5582) );
  XNOR U5952 ( .A(n5583), .B(n5582), .Z(n5534) );
  NANDN U5953 ( .A(n16746), .B(o[9]), .Z(n5532) );
  OR U5954 ( .A(n5421), .B(n5420), .Z(n5425) );
  OR U5955 ( .A(n5423), .B(n5422), .Z(n5424) );
  NAND U5956 ( .A(n5425), .B(n5424), .Z(n5533) );
  XOR U5957 ( .A(n5532), .B(n5533), .Z(n5535) );
  XNOR U5958 ( .A(n5534), .B(n5535), .Z(n5586) );
  XNOR U5959 ( .A(n5587), .B(n5586), .Z(n5588) );
  XNOR U5960 ( .A(n5589), .B(n5588), .Z(n5528) );
  NANDN U5961 ( .A(n16826), .B(o[11]), .Z(n5526) );
  OR U5962 ( .A(n5427), .B(n5426), .Z(n5431) );
  OR U5963 ( .A(n5429), .B(n5428), .Z(n5430) );
  NAND U5964 ( .A(n5431), .B(n5430), .Z(n5527) );
  XOR U5965 ( .A(n5526), .B(n5527), .Z(n5529) );
  XNOR U5966 ( .A(n5528), .B(n5529), .Z(n5592) );
  XNOR U5967 ( .A(n5593), .B(n5592), .Z(n5594) );
  XOR U5968 ( .A(n5595), .B(n5594), .Z(n5522) );
  AND U5969 ( .A(\stack[1][15] ), .B(o[13]), .Z(n5520) );
  OR U5970 ( .A(n5433), .B(n5432), .Z(n5437) );
  OR U5971 ( .A(n5435), .B(n5434), .Z(n5436) );
  NAND U5972 ( .A(n5437), .B(n5436), .Z(n5521) );
  XNOR U5973 ( .A(n5520), .B(n5521), .Z(n5523) );
  XNOR U5974 ( .A(n5598), .B(n5599), .Z(n5601) );
  XOR U5975 ( .A(n5600), .B(n5601), .Z(n5516) );
  NANDN U5976 ( .A(n5439), .B(n5438), .Z(n5443) );
  OR U5977 ( .A(n5441), .B(n5440), .Z(n5442) );
  AND U5978 ( .A(n5443), .B(n5442), .Z(n5515) );
  NANDN U5979 ( .A(n3009), .B(\stack[1][13] ), .Z(n5514) );
  XOR U5980 ( .A(n5515), .B(n5514), .Z(n5517) );
  XNOR U5981 ( .A(n5516), .B(n5517), .Z(n5604) );
  XNOR U5982 ( .A(n5605), .B(n5604), .Z(n5606) );
  XNOR U5983 ( .A(n5607), .B(n5606), .Z(n5510) );
  OR U5984 ( .A(n5445), .B(n5444), .Z(n5449) );
  NANDN U5985 ( .A(n5447), .B(n5446), .Z(n5448) );
  AND U5986 ( .A(n5449), .B(n5448), .Z(n5509) );
  NANDN U5987 ( .A(n3011), .B(\stack[1][11] ), .Z(n5508) );
  XOR U5988 ( .A(n5509), .B(n5508), .Z(n5511) );
  XNOR U5989 ( .A(n5510), .B(n5511), .Z(n5610) );
  XNOR U5990 ( .A(n5611), .B(n5610), .Z(n5612) );
  XNOR U5991 ( .A(n5613), .B(n5612), .Z(n5504) );
  NANDN U5992 ( .A(n3013), .B(\stack[1][9] ), .Z(n5502) );
  OR U5993 ( .A(n5451), .B(n5450), .Z(n5455) );
  OR U5994 ( .A(n5453), .B(n5452), .Z(n5454) );
  NAND U5995 ( .A(n5455), .B(n5454), .Z(n5503) );
  XOR U5996 ( .A(n5502), .B(n5503), .Z(n5505) );
  XNOR U5997 ( .A(n5504), .B(n5505), .Z(n5616) );
  XNOR U5998 ( .A(n5617), .B(n5616), .Z(n5618) );
  XNOR U5999 ( .A(n5619), .B(n5618), .Z(n5498) );
  NANDN U6000 ( .A(n3015), .B(\stack[1][7] ), .Z(n5496) );
  OR U6001 ( .A(n5457), .B(n5456), .Z(n5461) );
  OR U6002 ( .A(n5459), .B(n5458), .Z(n5460) );
  NAND U6003 ( .A(n5461), .B(n5460), .Z(n5497) );
  XOR U6004 ( .A(n5496), .B(n5497), .Z(n5499) );
  XNOR U6005 ( .A(n5498), .B(n5499), .Z(n5622) );
  XNOR U6006 ( .A(n5623), .B(n5622), .Z(n5624) );
  XOR U6007 ( .A(n5625), .B(n5624), .Z(n5492) );
  AND U6008 ( .A(o[23]), .B(\stack[1][5] ), .Z(n5490) );
  OR U6009 ( .A(n5463), .B(n5462), .Z(n5467) );
  OR U6010 ( .A(n5465), .B(n5464), .Z(n5466) );
  NAND U6011 ( .A(n5467), .B(n5466), .Z(n5491) );
  XNOR U6012 ( .A(n5490), .B(n5491), .Z(n5493) );
  XNOR U6013 ( .A(n5628), .B(n5629), .Z(n5630) );
  XNOR U6014 ( .A(n5631), .B(n5630), .Z(n5487) );
  OR U6015 ( .A(n5469), .B(n5468), .Z(n5473) );
  OR U6016 ( .A(n5471), .B(n5470), .Z(n5472) );
  AND U6017 ( .A(n5473), .B(n5472), .Z(n5479) );
  XNOR U6018 ( .A(n5478), .B(n5479), .Z(n5480) );
  AND U6019 ( .A(o[26]), .B(\stack[1][2] ), .Z(n5481) );
  XOR U6020 ( .A(n5637), .B(n5636), .Z(n5474) );
  NANDN U6021 ( .A(n5475), .B(n5474), .Z(n5477) );
  XOR U6022 ( .A(n5475), .B(n5474), .Z(n16396) );
  AND U6023 ( .A(o[28]), .B(\stack[1][0] ), .Z(n16397) );
  OR U6024 ( .A(n16396), .B(n16397), .Z(n5476) );
  AND U6025 ( .A(n5477), .B(n5476), .Z(n5641) );
  OR U6026 ( .A(n5640), .B(n5641), .Z(n5643) );
  OR U6027 ( .A(n5479), .B(n5478), .Z(n5483) );
  OR U6028 ( .A(n5481), .B(n5480), .Z(n5482) );
  NAND U6029 ( .A(n5483), .B(n5482), .Z(n5645) );
  ANDN U6030 ( .B(o[27]), .A(n2970), .Z(n5644) );
  XOR U6031 ( .A(n5645), .B(n5644), .Z(n5646) );
  NANDN U6032 ( .A(n17375), .B(o[26]), .Z(n5803) );
  NANDN U6033 ( .A(n5485), .B(n5484), .Z(n5489) );
  OR U6034 ( .A(n5487), .B(n5486), .Z(n5488) );
  AND U6035 ( .A(n5489), .B(n5488), .Z(n5800) );
  NANDN U6036 ( .A(n17296), .B(o[24]), .Z(n5797) );
  OR U6037 ( .A(n5491), .B(n5490), .Z(n5495) );
  OR U6038 ( .A(n5493), .B(n5492), .Z(n5494) );
  NAND U6039 ( .A(n5495), .B(n5494), .Z(n5795) );
  NANDN U6040 ( .A(n17219), .B(o[22]), .Z(n5791) );
  NANDN U6041 ( .A(n5497), .B(n5496), .Z(n5501) );
  NANDN U6042 ( .A(n5499), .B(n5498), .Z(n5500) );
  NAND U6043 ( .A(n5501), .B(n5500), .Z(n5789) );
  NANDN U6044 ( .A(n17145), .B(o[20]), .Z(n5785) );
  NANDN U6045 ( .A(n5503), .B(n5502), .Z(n5507) );
  NANDN U6046 ( .A(n5505), .B(n5504), .Z(n5506) );
  NAND U6047 ( .A(n5507), .B(n5506), .Z(n5783) );
  NANDN U6048 ( .A(n2972), .B(o[18]), .Z(n5779) );
  NANDN U6049 ( .A(n5509), .B(n5508), .Z(n5513) );
  NANDN U6050 ( .A(n5511), .B(n5510), .Z(n5512) );
  NAND U6051 ( .A(n5513), .B(n5512), .Z(n5777) );
  NANDN U6052 ( .A(n2974), .B(o[16]), .Z(n5773) );
  NANDN U6053 ( .A(n5515), .B(n5514), .Z(n5519) );
  NANDN U6054 ( .A(n5517), .B(n5516), .Z(n5518) );
  NAND U6055 ( .A(n5519), .B(n5518), .Z(n5771) );
  NANDN U6056 ( .A(n3008), .B(\stack[1][15] ), .Z(n5767) );
  OR U6057 ( .A(n5521), .B(n5520), .Z(n5525) );
  OR U6058 ( .A(n5523), .B(n5522), .Z(n5524) );
  NAND U6059 ( .A(n5525), .B(n5524), .Z(n5765) );
  NANDN U6060 ( .A(n3006), .B(\stack[1][17] ), .Z(n5761) );
  NANDN U6061 ( .A(n5527), .B(n5526), .Z(n5531) );
  NANDN U6062 ( .A(n5529), .B(n5528), .Z(n5530) );
  NAND U6063 ( .A(n5531), .B(n5530), .Z(n5759) );
  NANDN U6064 ( .A(n3004), .B(\stack[1][19] ), .Z(n5755) );
  NANDN U6065 ( .A(n5533), .B(n5532), .Z(n5537) );
  NANDN U6066 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U6067 ( .A(n5537), .B(n5536), .Z(n5753) );
  NANDN U6068 ( .A(n3002), .B(\stack[1][21] ), .Z(n5749) );
  OR U6069 ( .A(n5539), .B(n5538), .Z(n5543) );
  OR U6070 ( .A(n5541), .B(n5540), .Z(n5542) );
  NAND U6071 ( .A(n5543), .B(n5542), .Z(n5747) );
  OR U6072 ( .A(n5545), .B(n5544), .Z(n5549) );
  NANDN U6073 ( .A(n5547), .B(n5546), .Z(n5548) );
  AND U6074 ( .A(n5549), .B(n5548), .Z(n5704) );
  AND U6075 ( .A(\stack[1][22] ), .B(o[7]), .Z(n5705) );
  XNOR U6076 ( .A(n5704), .B(n5705), .Z(n5707) );
  OR U6077 ( .A(n5551), .B(n5550), .Z(n5555) );
  OR U6078 ( .A(n5553), .B(n5552), .Z(n5554) );
  AND U6079 ( .A(n5555), .B(n5554), .Z(n5710) );
  OR U6080 ( .A(n5557), .B(n5556), .Z(n5561) );
  OR U6081 ( .A(n5559), .B(n5558), .Z(n5560) );
  NAND U6082 ( .A(n5561), .B(n5560), .Z(n5741) );
  NANDN U6083 ( .A(n5563), .B(n5562), .Z(n5569) );
  ANDN U6084 ( .B(\stack[1][26] ), .A(n2994), .Z(n5565) );
  NAND U6085 ( .A(n5565), .B(n5564), .Z(n5567) );
  NANDN U6086 ( .A(n2983), .B(o[2]), .Z(n5566) );
  AND U6087 ( .A(n5567), .B(n5566), .Z(n5568) );
  ANDN U6088 ( .B(n5569), .A(n5568), .Z(n5722) );
  AND U6089 ( .A(\stack[1][26] ), .B(o[3]), .Z(n5723) );
  XNOR U6090 ( .A(n5722), .B(n5723), .Z(n5725) );
  ANDN U6091 ( .B(o[0]), .A(n2986), .Z(n5571) );
  NANDN U6092 ( .A(n2995), .B(\stack[1][28] ), .Z(n5570) );
  XNOR U6093 ( .A(n5571), .B(n5570), .Z(n5729) );
  AND U6094 ( .A(\stack[1][28] ), .B(o[1]), .Z(n5730) );
  NANDN U6095 ( .A(n2994), .B(n5730), .Z(n5572) );
  XOR U6096 ( .A(n2996), .B(n5572), .Z(n5573) );
  AND U6097 ( .A(n5573), .B(\stack[1][27] ), .Z(n5728) );
  XOR U6098 ( .A(n5729), .B(n5728), .Z(n5724) );
  XOR U6099 ( .A(n5725), .B(n5724), .Z(n5740) );
  XNOR U6100 ( .A(n5741), .B(n5740), .Z(n5743) );
  AND U6101 ( .A(\stack[1][25] ), .B(o[4]), .Z(n5742) );
  XNOR U6102 ( .A(n5743), .B(n5742), .Z(n5718) );
  AND U6103 ( .A(\stack[1][24] ), .B(o[5]), .Z(n5716) );
  OR U6104 ( .A(n5575), .B(n5574), .Z(n5579) );
  NANDN U6105 ( .A(n5577), .B(n5576), .Z(n5578) );
  NAND U6106 ( .A(n5579), .B(n5578), .Z(n5717) );
  XNOR U6107 ( .A(n5716), .B(n5717), .Z(n5719) );
  XNOR U6108 ( .A(n5718), .B(n5719), .Z(n5711) );
  XOR U6109 ( .A(n5710), .B(n5711), .Z(n5712) );
  AND U6110 ( .A(\stack[1][23] ), .B(o[6]), .Z(n5713) );
  XOR U6111 ( .A(n5712), .B(n5713), .Z(n5706) );
  XOR U6112 ( .A(n5707), .B(n5706), .Z(n5746) );
  XNOR U6113 ( .A(n5747), .B(n5746), .Z(n5748) );
  XNOR U6114 ( .A(n5749), .B(n5748), .Z(n5700) );
  NANDN U6115 ( .A(n16712), .B(o[9]), .Z(n5698) );
  OR U6116 ( .A(n5581), .B(n5580), .Z(n5585) );
  OR U6117 ( .A(n5583), .B(n5582), .Z(n5584) );
  NAND U6118 ( .A(n5585), .B(n5584), .Z(n5699) );
  XOR U6119 ( .A(n5698), .B(n5699), .Z(n5701) );
  XNOR U6120 ( .A(n5700), .B(n5701), .Z(n5752) );
  XNOR U6121 ( .A(n5753), .B(n5752), .Z(n5754) );
  XNOR U6122 ( .A(n5755), .B(n5754), .Z(n5694) );
  NANDN U6123 ( .A(n16786), .B(o[11]), .Z(n5692) );
  OR U6124 ( .A(n5587), .B(n5586), .Z(n5591) );
  OR U6125 ( .A(n5589), .B(n5588), .Z(n5590) );
  NAND U6126 ( .A(n5591), .B(n5590), .Z(n5693) );
  XOR U6127 ( .A(n5692), .B(n5693), .Z(n5695) );
  XNOR U6128 ( .A(n5694), .B(n5695), .Z(n5758) );
  XNOR U6129 ( .A(n5759), .B(n5758), .Z(n5760) );
  XNOR U6130 ( .A(n5761), .B(n5760), .Z(n5688) );
  NANDN U6131 ( .A(n2977), .B(o[13]), .Z(n5686) );
  OR U6132 ( .A(n5593), .B(n5592), .Z(n5597) );
  OR U6133 ( .A(n5595), .B(n5594), .Z(n5596) );
  NAND U6134 ( .A(n5597), .B(n5596), .Z(n5687) );
  XOR U6135 ( .A(n5686), .B(n5687), .Z(n5689) );
  XNOR U6136 ( .A(n5688), .B(n5689), .Z(n5764) );
  XNOR U6137 ( .A(n5765), .B(n5764), .Z(n5766) );
  XNOR U6138 ( .A(n5767), .B(n5766), .Z(n5682) );
  NANDN U6139 ( .A(n3009), .B(\stack[1][14] ), .Z(n5680) );
  OR U6140 ( .A(n5599), .B(n5598), .Z(n5603) );
  IV U6141 ( .A(n5600), .Z(n16944) );
  OR U6142 ( .A(n5601), .B(n16944), .Z(n5602) );
  NAND U6143 ( .A(n5603), .B(n5602), .Z(n5681) );
  XOR U6144 ( .A(n5680), .B(n5681), .Z(n5683) );
  XNOR U6145 ( .A(n5682), .B(n5683), .Z(n5770) );
  XNOR U6146 ( .A(n5771), .B(n5770), .Z(n5772) );
  XNOR U6147 ( .A(n5773), .B(n5772), .Z(n5676) );
  NANDN U6148 ( .A(n3011), .B(\stack[1][12] ), .Z(n5674) );
  OR U6149 ( .A(n5605), .B(n5604), .Z(n5609) );
  OR U6150 ( .A(n5607), .B(n5606), .Z(n5608) );
  NAND U6151 ( .A(n5609), .B(n5608), .Z(n5675) );
  XOR U6152 ( .A(n5674), .B(n5675), .Z(n5677) );
  XNOR U6153 ( .A(n5676), .B(n5677), .Z(n5776) );
  XNOR U6154 ( .A(n5777), .B(n5776), .Z(n5778) );
  XNOR U6155 ( .A(n5779), .B(n5778), .Z(n5670) );
  NANDN U6156 ( .A(n3013), .B(\stack[1][10] ), .Z(n5668) );
  OR U6157 ( .A(n5611), .B(n5610), .Z(n5615) );
  OR U6158 ( .A(n5613), .B(n5612), .Z(n5614) );
  NAND U6159 ( .A(n5615), .B(n5614), .Z(n5669) );
  XOR U6160 ( .A(n5668), .B(n5669), .Z(n5671) );
  XNOR U6161 ( .A(n5670), .B(n5671), .Z(n5782) );
  XNOR U6162 ( .A(n5783), .B(n5782), .Z(n5784) );
  XNOR U6163 ( .A(n5785), .B(n5784), .Z(n5664) );
  NANDN U6164 ( .A(n3015), .B(\stack[1][8] ), .Z(n5662) );
  OR U6165 ( .A(n5617), .B(n5616), .Z(n5621) );
  OR U6166 ( .A(n5619), .B(n5618), .Z(n5620) );
  NAND U6167 ( .A(n5621), .B(n5620), .Z(n5663) );
  XOR U6168 ( .A(n5662), .B(n5663), .Z(n5665) );
  XNOR U6169 ( .A(n5664), .B(n5665), .Z(n5788) );
  XNOR U6170 ( .A(n5789), .B(n5788), .Z(n5790) );
  XNOR U6171 ( .A(n5791), .B(n5790), .Z(n5658) );
  NANDN U6172 ( .A(n3017), .B(\stack[1][6] ), .Z(n5656) );
  OR U6173 ( .A(n5623), .B(n5622), .Z(n5627) );
  OR U6174 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U6175 ( .A(n5627), .B(n5626), .Z(n5657) );
  XOR U6176 ( .A(n5656), .B(n5657), .Z(n5659) );
  XNOR U6177 ( .A(n5658), .B(n5659), .Z(n5794) );
  XNOR U6178 ( .A(n5795), .B(n5794), .Z(n5796) );
  XOR U6179 ( .A(n5797), .B(n5796), .Z(n5652) );
  AND U6180 ( .A(o[25]), .B(\stack[1][4] ), .Z(n5650) );
  OR U6181 ( .A(n5629), .B(n5628), .Z(n5633) );
  OR U6182 ( .A(n5631), .B(n5630), .Z(n5632) );
  NAND U6183 ( .A(n5633), .B(n5632), .Z(n5651) );
  XNOR U6184 ( .A(n5650), .B(n5651), .Z(n5653) );
  XNOR U6185 ( .A(n5800), .B(n5801), .Z(n5802) );
  XNOR U6186 ( .A(n5803), .B(n5802), .Z(n5647) );
  OR U6187 ( .A(n5635), .B(n5634), .Z(n5639) );
  OR U6188 ( .A(n5637), .B(n5636), .Z(n5638) );
  AND U6189 ( .A(n5639), .B(n5638), .Z(n5807) );
  XOR U6190 ( .A(n5806), .B(n5807), .Z(n5808) );
  AND U6191 ( .A(o[28]), .B(\stack[1][1] ), .Z(n5809) );
  XOR U6192 ( .A(n5808), .B(n5809), .Z(n16360) );
  XNOR U6193 ( .A(n5641), .B(n5640), .Z(n16361) );
  OR U6194 ( .A(n16360), .B(n16361), .Z(n5642) );
  AND U6195 ( .A(n5643), .B(n5642), .Z(n5813) );
  NANDN U6196 ( .A(n2970), .B(o[28]), .Z(n5988) );
  NANDN U6197 ( .A(n5645), .B(n5644), .Z(n5649) );
  OR U6198 ( .A(n5647), .B(n5646), .Z(n5648) );
  AND U6199 ( .A(n5649), .B(n5648), .Z(n5985) );
  NANDN U6200 ( .A(n2971), .B(o[26]), .Z(n5982) );
  OR U6201 ( .A(n5651), .B(n5650), .Z(n5655) );
  OR U6202 ( .A(n5653), .B(n5652), .Z(n5654) );
  NAND U6203 ( .A(n5655), .B(n5654), .Z(n5980) );
  NANDN U6204 ( .A(n17256), .B(o[24]), .Z(n5976) );
  NANDN U6205 ( .A(n5657), .B(n5656), .Z(n5661) );
  NANDN U6206 ( .A(n5659), .B(n5658), .Z(n5660) );
  NAND U6207 ( .A(n5661), .B(n5660), .Z(n5974) );
  NANDN U6208 ( .A(n17179), .B(o[22]), .Z(n5970) );
  NANDN U6209 ( .A(n5663), .B(n5662), .Z(n5667) );
  NANDN U6210 ( .A(n5665), .B(n5664), .Z(n5666) );
  NAND U6211 ( .A(n5667), .B(n5666), .Z(n5968) );
  NANDN U6212 ( .A(n17101), .B(o[20]), .Z(n5964) );
  NANDN U6213 ( .A(n5669), .B(n5668), .Z(n5673) );
  NANDN U6214 ( .A(n5671), .B(n5670), .Z(n5672) );
  NAND U6215 ( .A(n5673), .B(n5672), .Z(n5962) );
  NANDN U6216 ( .A(n2973), .B(o[18]), .Z(n5958) );
  NANDN U6217 ( .A(n5675), .B(n5674), .Z(n5679) );
  NANDN U6218 ( .A(n5677), .B(n5676), .Z(n5678) );
  NAND U6219 ( .A(n5679), .B(n5678), .Z(n5956) );
  NANDN U6220 ( .A(n2975), .B(o[16]), .Z(n5952) );
  NANDN U6221 ( .A(n5681), .B(n5680), .Z(n5685) );
  NANDN U6222 ( .A(n5683), .B(n5682), .Z(n5684) );
  NAND U6223 ( .A(n5685), .B(n5684), .Z(n5950) );
  NANDN U6224 ( .A(n3008), .B(\stack[1][16] ), .Z(n5946) );
  NANDN U6225 ( .A(n5687), .B(n5686), .Z(n5691) );
  NANDN U6226 ( .A(n5689), .B(n5688), .Z(n5690) );
  NAND U6227 ( .A(n5691), .B(n5690), .Z(n5944) );
  NANDN U6228 ( .A(n3006), .B(\stack[1][18] ), .Z(n5940) );
  NANDN U6229 ( .A(n5693), .B(n5692), .Z(n5697) );
  NANDN U6230 ( .A(n5695), .B(n5694), .Z(n5696) );
  NAND U6231 ( .A(n5697), .B(n5696), .Z(n5938) );
  NANDN U6232 ( .A(n3004), .B(\stack[1][20] ), .Z(n5934) );
  NANDN U6233 ( .A(n5699), .B(n5698), .Z(n5703) );
  NANDN U6234 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U6235 ( .A(n5703), .B(n5702), .Z(n5932) );
  NANDN U6236 ( .A(n3002), .B(\stack[1][22] ), .Z(n5928) );
  OR U6237 ( .A(n5705), .B(n5704), .Z(n5709) );
  OR U6238 ( .A(n5707), .B(n5706), .Z(n5708) );
  NAND U6239 ( .A(n5709), .B(n5708), .Z(n5926) );
  OR U6240 ( .A(n5711), .B(n5710), .Z(n5715) );
  NANDN U6241 ( .A(n5713), .B(n5712), .Z(n5714) );
  AND U6242 ( .A(n5715), .B(n5714), .Z(n5883) );
  AND U6243 ( .A(\stack[1][23] ), .B(o[7]), .Z(n5884) );
  XNOR U6244 ( .A(n5883), .B(n5884), .Z(n5886) );
  OR U6245 ( .A(n5717), .B(n5716), .Z(n5721) );
  OR U6246 ( .A(n5719), .B(n5718), .Z(n5720) );
  AND U6247 ( .A(n5721), .B(n5720), .Z(n5889) );
  OR U6248 ( .A(n5723), .B(n5722), .Z(n5727) );
  OR U6249 ( .A(n5725), .B(n5724), .Z(n5726) );
  NAND U6250 ( .A(n5727), .B(n5726), .Z(n5920) );
  NANDN U6251 ( .A(n5729), .B(n5728), .Z(n5735) );
  ANDN U6252 ( .B(\stack[1][27] ), .A(n2994), .Z(n5731) );
  NAND U6253 ( .A(n5731), .B(n5730), .Z(n5733) );
  NANDN U6254 ( .A(n2984), .B(o[2]), .Z(n5732) );
  AND U6255 ( .A(n5733), .B(n5732), .Z(n5734) );
  ANDN U6256 ( .B(n5735), .A(n5734), .Z(n5901) );
  AND U6257 ( .A(\stack[1][27] ), .B(o[3]), .Z(n5902) );
  XNOR U6258 ( .A(n5901), .B(n5902), .Z(n5904) );
  ANDN U6259 ( .B(o[0]), .A(n2987), .Z(n5737) );
  NANDN U6260 ( .A(n2995), .B(\stack[1][29] ), .Z(n5736) );
  XNOR U6261 ( .A(n5737), .B(n5736), .Z(n5908) );
  AND U6262 ( .A(\stack[1][29] ), .B(o[1]), .Z(n5909) );
  NANDN U6263 ( .A(n2994), .B(n5909), .Z(n5738) );
  XOR U6264 ( .A(n2996), .B(n5738), .Z(n5739) );
  AND U6265 ( .A(n5739), .B(\stack[1][28] ), .Z(n5907) );
  XOR U6266 ( .A(n5908), .B(n5907), .Z(n5903) );
  XOR U6267 ( .A(n5904), .B(n5903), .Z(n5919) );
  XNOR U6268 ( .A(n5920), .B(n5919), .Z(n5922) );
  AND U6269 ( .A(\stack[1][26] ), .B(o[4]), .Z(n5921) );
  XNOR U6270 ( .A(n5922), .B(n5921), .Z(n5897) );
  AND U6271 ( .A(\stack[1][25] ), .B(o[5]), .Z(n5895) );
  OR U6272 ( .A(n5741), .B(n5740), .Z(n5745) );
  NANDN U6273 ( .A(n5743), .B(n5742), .Z(n5744) );
  NAND U6274 ( .A(n5745), .B(n5744), .Z(n5896) );
  XNOR U6275 ( .A(n5895), .B(n5896), .Z(n5898) );
  XNOR U6276 ( .A(n5897), .B(n5898), .Z(n5890) );
  XOR U6277 ( .A(n5889), .B(n5890), .Z(n5891) );
  AND U6278 ( .A(\stack[1][24] ), .B(o[6]), .Z(n5892) );
  XOR U6279 ( .A(n5891), .B(n5892), .Z(n5885) );
  XOR U6280 ( .A(n5886), .B(n5885), .Z(n5925) );
  XNOR U6281 ( .A(n5926), .B(n5925), .Z(n5927) );
  XNOR U6282 ( .A(n5928), .B(n5927), .Z(n5879) );
  NANDN U6283 ( .A(n2978), .B(o[9]), .Z(n5877) );
  OR U6284 ( .A(n5747), .B(n5746), .Z(n5751) );
  OR U6285 ( .A(n5749), .B(n5748), .Z(n5750) );
  NAND U6286 ( .A(n5751), .B(n5750), .Z(n5878) );
  XOR U6287 ( .A(n5877), .B(n5878), .Z(n5880) );
  XNOR U6288 ( .A(n5879), .B(n5880), .Z(n5931) );
  XNOR U6289 ( .A(n5932), .B(n5931), .Z(n5933) );
  XNOR U6290 ( .A(n5934), .B(n5933), .Z(n5873) );
  NANDN U6291 ( .A(n16746), .B(o[11]), .Z(n5871) );
  OR U6292 ( .A(n5753), .B(n5752), .Z(n5757) );
  OR U6293 ( .A(n5755), .B(n5754), .Z(n5756) );
  NAND U6294 ( .A(n5757), .B(n5756), .Z(n5872) );
  XOR U6295 ( .A(n5871), .B(n5872), .Z(n5874) );
  XNOR U6296 ( .A(n5873), .B(n5874), .Z(n5937) );
  XNOR U6297 ( .A(n5938), .B(n5937), .Z(n5939) );
  XNOR U6298 ( .A(n5940), .B(n5939), .Z(n5867) );
  NANDN U6299 ( .A(n16826), .B(o[13]), .Z(n5865) );
  OR U6300 ( .A(n5759), .B(n5758), .Z(n5763) );
  OR U6301 ( .A(n5761), .B(n5760), .Z(n5762) );
  NAND U6302 ( .A(n5763), .B(n5762), .Z(n5866) );
  XOR U6303 ( .A(n5865), .B(n5866), .Z(n5868) );
  XNOR U6304 ( .A(n5867), .B(n5868), .Z(n5943) );
  XNOR U6305 ( .A(n5944), .B(n5943), .Z(n5945) );
  XNOR U6306 ( .A(n5946), .B(n5945), .Z(n5861) );
  AND U6307 ( .A(o[15]), .B(\stack[1][15] ), .Z(n16905) );
  OR U6308 ( .A(n5765), .B(n5764), .Z(n5769) );
  OR U6309 ( .A(n5767), .B(n5766), .Z(n5768) );
  NAND U6310 ( .A(n5769), .B(n5768), .Z(n5860) );
  XNOR U6311 ( .A(n16905), .B(n5860), .Z(n5862) );
  XNOR U6312 ( .A(n5861), .B(n5862), .Z(n5949) );
  XNOR U6313 ( .A(n5950), .B(n5949), .Z(n5951) );
  XNOR U6314 ( .A(n5952), .B(n5951), .Z(n5856) );
  NANDN U6315 ( .A(n3011), .B(\stack[1][13] ), .Z(n5854) );
  OR U6316 ( .A(n5771), .B(n5770), .Z(n5775) );
  OR U6317 ( .A(n5773), .B(n5772), .Z(n5774) );
  NAND U6318 ( .A(n5775), .B(n5774), .Z(n5855) );
  XOR U6319 ( .A(n5854), .B(n5855), .Z(n5857) );
  XNOR U6320 ( .A(n5856), .B(n5857), .Z(n5955) );
  XNOR U6321 ( .A(n5956), .B(n5955), .Z(n5957) );
  XNOR U6322 ( .A(n5958), .B(n5957), .Z(n5850) );
  NANDN U6323 ( .A(n3013), .B(\stack[1][11] ), .Z(n5848) );
  OR U6324 ( .A(n5777), .B(n5776), .Z(n5781) );
  OR U6325 ( .A(n5779), .B(n5778), .Z(n5780) );
  NAND U6326 ( .A(n5781), .B(n5780), .Z(n5849) );
  XOR U6327 ( .A(n5848), .B(n5849), .Z(n5851) );
  XNOR U6328 ( .A(n5850), .B(n5851), .Z(n5961) );
  XNOR U6329 ( .A(n5962), .B(n5961), .Z(n5963) );
  XNOR U6330 ( .A(n5964), .B(n5963), .Z(n5844) );
  NANDN U6331 ( .A(n3015), .B(\stack[1][9] ), .Z(n5842) );
  OR U6332 ( .A(n5783), .B(n5782), .Z(n5787) );
  OR U6333 ( .A(n5785), .B(n5784), .Z(n5786) );
  NAND U6334 ( .A(n5787), .B(n5786), .Z(n5843) );
  XOR U6335 ( .A(n5842), .B(n5843), .Z(n5845) );
  XNOR U6336 ( .A(n5844), .B(n5845), .Z(n5967) );
  XNOR U6337 ( .A(n5968), .B(n5967), .Z(n5969) );
  XNOR U6338 ( .A(n5970), .B(n5969), .Z(n5838) );
  NANDN U6339 ( .A(n3017), .B(\stack[1][7] ), .Z(n5836) );
  OR U6340 ( .A(n5789), .B(n5788), .Z(n5793) );
  OR U6341 ( .A(n5791), .B(n5790), .Z(n5792) );
  NAND U6342 ( .A(n5793), .B(n5792), .Z(n5837) );
  XOR U6343 ( .A(n5836), .B(n5837), .Z(n5839) );
  XNOR U6344 ( .A(n5838), .B(n5839), .Z(n5973) );
  XNOR U6345 ( .A(n5974), .B(n5973), .Z(n5975) );
  XNOR U6346 ( .A(n5976), .B(n5975), .Z(n5832) );
  NANDN U6347 ( .A(n3019), .B(\stack[1][5] ), .Z(n5830) );
  OR U6348 ( .A(n5795), .B(n5794), .Z(n5799) );
  OR U6349 ( .A(n5797), .B(n5796), .Z(n5798) );
  NAND U6350 ( .A(n5799), .B(n5798), .Z(n5831) );
  XOR U6351 ( .A(n5830), .B(n5831), .Z(n5833) );
  XNOR U6352 ( .A(n5832), .B(n5833), .Z(n5979) );
  XNOR U6353 ( .A(n5980), .B(n5979), .Z(n5981) );
  XNOR U6354 ( .A(n5982), .B(n5981), .Z(n5826) );
  NANDN U6355 ( .A(n17375), .B(o[27]), .Z(n5824) );
  OR U6356 ( .A(n5801), .B(n5800), .Z(n5805) );
  OR U6357 ( .A(n5803), .B(n5802), .Z(n5804) );
  NAND U6358 ( .A(n5805), .B(n5804), .Z(n5825) );
  XOR U6359 ( .A(n5824), .B(n5825), .Z(n5827) );
  XNOR U6360 ( .A(n5826), .B(n5827), .Z(n5986) );
  XNOR U6361 ( .A(n5985), .B(n5986), .Z(n5987) );
  XOR U6362 ( .A(n5988), .B(n5987), .Z(n5820) );
  OR U6363 ( .A(n5807), .B(n5806), .Z(n5811) );
  NANDN U6364 ( .A(n5809), .B(n5808), .Z(n5810) );
  AND U6365 ( .A(n5811), .B(n5810), .Z(n5818) );
  AND U6366 ( .A(o[29]), .B(\stack[1][1] ), .Z(n5819) );
  XNOR U6367 ( .A(n5818), .B(n5819), .Z(n5821) );
  XOR U6368 ( .A(n5820), .B(n5821), .Z(n5812) );
  NANDN U6369 ( .A(n5813), .B(n5812), .Z(n5815) );
  XOR U6370 ( .A(n5813), .B(n5812), .Z(n16320) );
  AND U6371 ( .A(o[30]), .B(\stack[1][0] ), .Z(n16321) );
  OR U6372 ( .A(n16320), .B(n16321), .Z(n5814) );
  AND U6373 ( .A(n5815), .B(n5814), .Z(n5817) );
  OR U6374 ( .A(n5816), .B(n5817), .Z(n5992) );
  XNOR U6375 ( .A(n5817), .B(n5816), .Z(n16280) );
  NANDN U6376 ( .A(n2969), .B(o[30]), .Z(n6170) );
  OR U6377 ( .A(n5819), .B(n5818), .Z(n5823) );
  OR U6378 ( .A(n5821), .B(n5820), .Z(n5822) );
  NAND U6379 ( .A(n5823), .B(n5822), .Z(n6168) );
  NANDN U6380 ( .A(n17375), .B(o[28]), .Z(n6164) );
  NANDN U6381 ( .A(n5825), .B(n5824), .Z(n5829) );
  NANDN U6382 ( .A(n5827), .B(n5826), .Z(n5828) );
  NAND U6383 ( .A(n5829), .B(n5828), .Z(n6162) );
  NANDN U6384 ( .A(n17296), .B(o[26]), .Z(n6158) );
  NANDN U6385 ( .A(n5831), .B(n5830), .Z(n5835) );
  NANDN U6386 ( .A(n5833), .B(n5832), .Z(n5834) );
  NAND U6387 ( .A(n5835), .B(n5834), .Z(n6156) );
  NANDN U6388 ( .A(n17219), .B(o[24]), .Z(n6152) );
  NANDN U6389 ( .A(n5837), .B(n5836), .Z(n5841) );
  NANDN U6390 ( .A(n5839), .B(n5838), .Z(n5840) );
  NAND U6391 ( .A(n5841), .B(n5840), .Z(n6150) );
  NANDN U6392 ( .A(n17145), .B(o[22]), .Z(n6146) );
  NANDN U6393 ( .A(n5843), .B(n5842), .Z(n5847) );
  NANDN U6394 ( .A(n5845), .B(n5844), .Z(n5846) );
  NAND U6395 ( .A(n5847), .B(n5846), .Z(n6144) );
  NANDN U6396 ( .A(n2972), .B(o[20]), .Z(n6140) );
  NANDN U6397 ( .A(n5849), .B(n5848), .Z(n5853) );
  NANDN U6398 ( .A(n5851), .B(n5850), .Z(n5852) );
  NAND U6399 ( .A(n5853), .B(n5852), .Z(n6138) );
  NANDN U6400 ( .A(n2974), .B(o[18]), .Z(n6134) );
  NANDN U6401 ( .A(n5855), .B(n5854), .Z(n5859) );
  NANDN U6402 ( .A(n5857), .B(n5856), .Z(n5858) );
  NAND U6403 ( .A(n5859), .B(n5858), .Z(n6132) );
  NANDN U6404 ( .A(n2976), .B(o[16]), .Z(n6128) );
  OR U6405 ( .A(n5860), .B(n16905), .Z(n5864) );
  NANDN U6406 ( .A(n5862), .B(n5861), .Z(n5863) );
  NAND U6407 ( .A(n5864), .B(n5863), .Z(n6126) );
  NANDN U6408 ( .A(n3008), .B(\stack[1][17] ), .Z(n6122) );
  NANDN U6409 ( .A(n5866), .B(n5865), .Z(n5870) );
  NANDN U6410 ( .A(n5868), .B(n5867), .Z(n5869) );
  NAND U6411 ( .A(n5870), .B(n5869), .Z(n6120) );
  NANDN U6412 ( .A(n3006), .B(\stack[1][19] ), .Z(n6116) );
  NANDN U6413 ( .A(n5872), .B(n5871), .Z(n5876) );
  NANDN U6414 ( .A(n5874), .B(n5873), .Z(n5875) );
  NAND U6415 ( .A(n5876), .B(n5875), .Z(n6114) );
  NANDN U6416 ( .A(n3004), .B(\stack[1][21] ), .Z(n6056) );
  NANDN U6417 ( .A(n5878), .B(n5877), .Z(n5882) );
  NANDN U6418 ( .A(n5880), .B(n5879), .Z(n5881) );
  NAND U6419 ( .A(n5882), .B(n5881), .Z(n6054) );
  NANDN U6420 ( .A(n3002), .B(\stack[1][23] ), .Z(n6110) );
  OR U6421 ( .A(n5884), .B(n5883), .Z(n5888) );
  OR U6422 ( .A(n5886), .B(n5885), .Z(n5887) );
  NAND U6423 ( .A(n5888), .B(n5887), .Z(n6108) );
  OR U6424 ( .A(n5890), .B(n5889), .Z(n5894) );
  NANDN U6425 ( .A(n5892), .B(n5891), .Z(n5893) );
  AND U6426 ( .A(n5894), .B(n5893), .Z(n6065) );
  AND U6427 ( .A(\stack[1][24] ), .B(o[7]), .Z(n6066) );
  XNOR U6428 ( .A(n6065), .B(n6066), .Z(n6068) );
  OR U6429 ( .A(n5896), .B(n5895), .Z(n5900) );
  OR U6430 ( .A(n5898), .B(n5897), .Z(n5899) );
  AND U6431 ( .A(n5900), .B(n5899), .Z(n6071) );
  OR U6432 ( .A(n5902), .B(n5901), .Z(n5906) );
  OR U6433 ( .A(n5904), .B(n5903), .Z(n5905) );
  NAND U6434 ( .A(n5906), .B(n5905), .Z(n6102) );
  NANDN U6435 ( .A(n5908), .B(n5907), .Z(n5914) );
  ANDN U6436 ( .B(\stack[1][28] ), .A(n2994), .Z(n5910) );
  NAND U6437 ( .A(n5910), .B(n5909), .Z(n5912) );
  NANDN U6438 ( .A(n2985), .B(o[2]), .Z(n5911) );
  AND U6439 ( .A(n5912), .B(n5911), .Z(n5913) );
  ANDN U6440 ( .B(n5914), .A(n5913), .Z(n6083) );
  AND U6441 ( .A(\stack[1][28] ), .B(o[3]), .Z(n6084) );
  XNOR U6442 ( .A(n6083), .B(n6084), .Z(n6086) );
  ANDN U6443 ( .B(o[0]), .A(n2988), .Z(n5916) );
  NANDN U6444 ( .A(n2995), .B(\stack[1][30] ), .Z(n5915) );
  XNOR U6445 ( .A(n5916), .B(n5915), .Z(n6090) );
  AND U6446 ( .A(\stack[1][30] ), .B(o[1]), .Z(n6091) );
  NANDN U6447 ( .A(n2994), .B(n6091), .Z(n5917) );
  XOR U6448 ( .A(n2996), .B(n5917), .Z(n5918) );
  AND U6449 ( .A(n5918), .B(\stack[1][29] ), .Z(n6089) );
  XOR U6450 ( .A(n6090), .B(n6089), .Z(n6085) );
  XOR U6451 ( .A(n6086), .B(n6085), .Z(n6101) );
  XNOR U6452 ( .A(n6102), .B(n6101), .Z(n6104) );
  AND U6453 ( .A(\stack[1][27] ), .B(o[4]), .Z(n6103) );
  XNOR U6454 ( .A(n6104), .B(n6103), .Z(n6079) );
  AND U6455 ( .A(\stack[1][26] ), .B(o[5]), .Z(n6077) );
  OR U6456 ( .A(n5920), .B(n5919), .Z(n5924) );
  NANDN U6457 ( .A(n5922), .B(n5921), .Z(n5923) );
  NAND U6458 ( .A(n5924), .B(n5923), .Z(n6078) );
  XNOR U6459 ( .A(n6077), .B(n6078), .Z(n6080) );
  XNOR U6460 ( .A(n6079), .B(n6080), .Z(n6072) );
  XOR U6461 ( .A(n6071), .B(n6072), .Z(n6073) );
  AND U6462 ( .A(\stack[1][25] ), .B(o[6]), .Z(n6074) );
  XOR U6463 ( .A(n6073), .B(n6074), .Z(n6067) );
  XOR U6464 ( .A(n6068), .B(n6067), .Z(n6107) );
  XNOR U6465 ( .A(n6108), .B(n6107), .Z(n6109) );
  XNOR U6466 ( .A(n6110), .B(n6109), .Z(n6061) );
  NANDN U6467 ( .A(n2979), .B(o[9]), .Z(n6059) );
  OR U6468 ( .A(n5926), .B(n5925), .Z(n5930) );
  OR U6469 ( .A(n5928), .B(n5927), .Z(n5929) );
  NAND U6470 ( .A(n5930), .B(n5929), .Z(n6060) );
  XOR U6471 ( .A(n6059), .B(n6060), .Z(n6062) );
  XNOR U6472 ( .A(n6061), .B(n6062), .Z(n6053) );
  XNOR U6473 ( .A(n6054), .B(n6053), .Z(n6055) );
  XNOR U6474 ( .A(n6056), .B(n6055), .Z(n6049) );
  NANDN U6475 ( .A(n16712), .B(o[11]), .Z(n6047) );
  OR U6476 ( .A(n5932), .B(n5931), .Z(n5936) );
  OR U6477 ( .A(n5934), .B(n5933), .Z(n5935) );
  NAND U6478 ( .A(n5936), .B(n5935), .Z(n6048) );
  XOR U6479 ( .A(n6047), .B(n6048), .Z(n6050) );
  XNOR U6480 ( .A(n6049), .B(n6050), .Z(n6113) );
  XNOR U6481 ( .A(n6114), .B(n6113), .Z(n6115) );
  XNOR U6482 ( .A(n6116), .B(n6115), .Z(n6043) );
  NANDN U6483 ( .A(n16786), .B(o[13]), .Z(n6041) );
  OR U6484 ( .A(n5938), .B(n5937), .Z(n5942) );
  OR U6485 ( .A(n5940), .B(n5939), .Z(n5941) );
  NAND U6486 ( .A(n5942), .B(n5941), .Z(n6042) );
  XOR U6487 ( .A(n6041), .B(n6042), .Z(n6044) );
  XNOR U6488 ( .A(n6043), .B(n6044), .Z(n6119) );
  XNOR U6489 ( .A(n6120), .B(n6119), .Z(n6121) );
  XNOR U6490 ( .A(n6122), .B(n6121), .Z(n6037) );
  NANDN U6491 ( .A(n2977), .B(o[15]), .Z(n6035) );
  OR U6492 ( .A(n5944), .B(n5943), .Z(n5948) );
  OR U6493 ( .A(n5946), .B(n5945), .Z(n5947) );
  NAND U6494 ( .A(n5948), .B(n5947), .Z(n6036) );
  XOR U6495 ( .A(n6035), .B(n6036), .Z(n6038) );
  XNOR U6496 ( .A(n6037), .B(n6038), .Z(n6125) );
  XNOR U6497 ( .A(n6126), .B(n6125), .Z(n6127) );
  XNOR U6498 ( .A(n6128), .B(n6127), .Z(n6031) );
  NANDN U6499 ( .A(n3011), .B(\stack[1][14] ), .Z(n6029) );
  OR U6500 ( .A(n5950), .B(n5949), .Z(n5954) );
  OR U6501 ( .A(n5952), .B(n5951), .Z(n5953) );
  NAND U6502 ( .A(n5954), .B(n5953), .Z(n6030) );
  XOR U6503 ( .A(n6029), .B(n6030), .Z(n6032) );
  XNOR U6504 ( .A(n6031), .B(n6032), .Z(n6131) );
  XNOR U6505 ( .A(n6132), .B(n6131), .Z(n6133) );
  XNOR U6506 ( .A(n6134), .B(n6133), .Z(n6025) );
  NANDN U6507 ( .A(n3013), .B(\stack[1][12] ), .Z(n6023) );
  OR U6508 ( .A(n5956), .B(n5955), .Z(n5960) );
  OR U6509 ( .A(n5958), .B(n5957), .Z(n5959) );
  NAND U6510 ( .A(n5960), .B(n5959), .Z(n6024) );
  XOR U6511 ( .A(n6023), .B(n6024), .Z(n6026) );
  XNOR U6512 ( .A(n6025), .B(n6026), .Z(n6137) );
  XNOR U6513 ( .A(n6138), .B(n6137), .Z(n6139) );
  XNOR U6514 ( .A(n6140), .B(n6139), .Z(n6019) );
  NANDN U6515 ( .A(n3015), .B(\stack[1][10] ), .Z(n6017) );
  OR U6516 ( .A(n5962), .B(n5961), .Z(n5966) );
  OR U6517 ( .A(n5964), .B(n5963), .Z(n5965) );
  NAND U6518 ( .A(n5966), .B(n5965), .Z(n6018) );
  XOR U6519 ( .A(n6017), .B(n6018), .Z(n6020) );
  XNOR U6520 ( .A(n6019), .B(n6020), .Z(n6143) );
  XNOR U6521 ( .A(n6144), .B(n6143), .Z(n6145) );
  XNOR U6522 ( .A(n6146), .B(n6145), .Z(n6013) );
  NANDN U6523 ( .A(n3017), .B(\stack[1][8] ), .Z(n6011) );
  OR U6524 ( .A(n5968), .B(n5967), .Z(n5972) );
  OR U6525 ( .A(n5970), .B(n5969), .Z(n5971) );
  NAND U6526 ( .A(n5972), .B(n5971), .Z(n6012) );
  XOR U6527 ( .A(n6011), .B(n6012), .Z(n6014) );
  XNOR U6528 ( .A(n6013), .B(n6014), .Z(n6149) );
  XNOR U6529 ( .A(n6150), .B(n6149), .Z(n6151) );
  XNOR U6530 ( .A(n6152), .B(n6151), .Z(n6007) );
  NANDN U6531 ( .A(n3019), .B(\stack[1][6] ), .Z(n6005) );
  OR U6532 ( .A(n5974), .B(n5973), .Z(n5978) );
  OR U6533 ( .A(n5976), .B(n5975), .Z(n5977) );
  NAND U6534 ( .A(n5978), .B(n5977), .Z(n6006) );
  XOR U6535 ( .A(n6005), .B(n6006), .Z(n6008) );
  XNOR U6536 ( .A(n6007), .B(n6008), .Z(n6155) );
  XNOR U6537 ( .A(n6156), .B(n6155), .Z(n6157) );
  XNOR U6538 ( .A(n6158), .B(n6157), .Z(n6001) );
  AND U6539 ( .A(o[27]), .B(\stack[1][4] ), .Z(n5999) );
  OR U6540 ( .A(n5980), .B(n5979), .Z(n5984) );
  OR U6541 ( .A(n5982), .B(n5981), .Z(n5983) );
  NAND U6542 ( .A(n5984), .B(n5983), .Z(n6000) );
  XNOR U6543 ( .A(n5999), .B(n6000), .Z(n6002) );
  XNOR U6544 ( .A(n6001), .B(n6002), .Z(n6161) );
  XNOR U6545 ( .A(n6162), .B(n6161), .Z(n6163) );
  XOR U6546 ( .A(n6164), .B(n6163), .Z(n5996) );
  AND U6547 ( .A(o[29]), .B(\stack[1][2] ), .Z(n5993) );
  OR U6548 ( .A(n5986), .B(n5985), .Z(n5990) );
  OR U6549 ( .A(n5988), .B(n5987), .Z(n5989) );
  NAND U6550 ( .A(n5990), .B(n5989), .Z(n5994) );
  XOR U6551 ( .A(n5993), .B(n5994), .Z(n5995) );
  XNOR U6552 ( .A(n5996), .B(n5995), .Z(n6167) );
  XNOR U6553 ( .A(n6168), .B(n6167), .Z(n6169) );
  XOR U6554 ( .A(n6170), .B(n6169), .Z(n16281) );
  OR U6555 ( .A(n16280), .B(n16281), .Z(n5991) );
  AND U6556 ( .A(n5992), .B(n5991), .Z(n6174) );
  NANDN U6557 ( .A(n2970), .B(o[30]), .Z(n6362) );
  OR U6558 ( .A(n5994), .B(n5993), .Z(n5998) );
  NANDN U6559 ( .A(n5996), .B(n5995), .Z(n5997) );
  NAND U6560 ( .A(n5998), .B(n5997), .Z(n6360) );
  NANDN U6561 ( .A(n2971), .B(o[28]), .Z(n6356) );
  OR U6562 ( .A(n6000), .B(n5999), .Z(n6004) );
  NANDN U6563 ( .A(n6002), .B(n6001), .Z(n6003) );
  NAND U6564 ( .A(n6004), .B(n6003), .Z(n6354) );
  NANDN U6565 ( .A(n17256), .B(o[26]), .Z(n6350) );
  NANDN U6566 ( .A(n6006), .B(n6005), .Z(n6010) );
  NANDN U6567 ( .A(n6008), .B(n6007), .Z(n6009) );
  NAND U6568 ( .A(n6010), .B(n6009), .Z(n6348) );
  NANDN U6569 ( .A(n17179), .B(o[24]), .Z(n6344) );
  NANDN U6570 ( .A(n6012), .B(n6011), .Z(n6016) );
  NANDN U6571 ( .A(n6014), .B(n6013), .Z(n6015) );
  NAND U6572 ( .A(n6016), .B(n6015), .Z(n6342) );
  NANDN U6573 ( .A(n17101), .B(o[22]), .Z(n6338) );
  NANDN U6574 ( .A(n6018), .B(n6017), .Z(n6022) );
  NANDN U6575 ( .A(n6020), .B(n6019), .Z(n6021) );
  NAND U6576 ( .A(n6022), .B(n6021), .Z(n6336) );
  NANDN U6577 ( .A(n2973), .B(o[20]), .Z(n6332) );
  NANDN U6578 ( .A(n6024), .B(n6023), .Z(n6028) );
  NANDN U6579 ( .A(n6026), .B(n6025), .Z(n6027) );
  NAND U6580 ( .A(n6028), .B(n6027), .Z(n6330) );
  NANDN U6581 ( .A(n2975), .B(o[18]), .Z(n6326) );
  NANDN U6582 ( .A(n6030), .B(n6029), .Z(n6034) );
  NANDN U6583 ( .A(n6032), .B(n6031), .Z(n6033) );
  NAND U6584 ( .A(n6034), .B(n6033), .Z(n6324) );
  NOR U6585 ( .A(n3010), .B(n2977), .Z(n6319) );
  NANDN U6586 ( .A(n6036), .B(n6035), .Z(n6040) );
  NANDN U6587 ( .A(n6038), .B(n6037), .Z(n6039) );
  NAND U6588 ( .A(n6040), .B(n6039), .Z(n6318) );
  NANDN U6589 ( .A(n3008), .B(\stack[1][18] ), .Z(n6314) );
  NANDN U6590 ( .A(n6042), .B(n6041), .Z(n6046) );
  NANDN U6591 ( .A(n6044), .B(n6043), .Z(n6045) );
  NAND U6592 ( .A(n6046), .B(n6045), .Z(n6312) );
  AND U6593 ( .A(\stack[1][20] ), .B(o[12]), .Z(n6308) );
  NANDN U6594 ( .A(n6048), .B(n6047), .Z(n6052) );
  NANDN U6595 ( .A(n6050), .B(n6049), .Z(n6051) );
  AND U6596 ( .A(n6052), .B(n6051), .Z(n6305) );
  AND U6597 ( .A(\stack[1][21] ), .B(o[11]), .Z(n6239) );
  OR U6598 ( .A(n6054), .B(n6053), .Z(n6058) );
  OR U6599 ( .A(n6056), .B(n6055), .Z(n6057) );
  NAND U6600 ( .A(n6058), .B(n6057), .Z(n6240) );
  XNOR U6601 ( .A(n6239), .B(n6240), .Z(n6242) );
  NANDN U6602 ( .A(n6060), .B(n6059), .Z(n6064) );
  NANDN U6603 ( .A(n6062), .B(n6061), .Z(n6063) );
  AND U6604 ( .A(n6064), .B(n6063), .Z(n6245) );
  OR U6605 ( .A(n6066), .B(n6065), .Z(n6070) );
  OR U6606 ( .A(n6068), .B(n6067), .Z(n6069) );
  NAND U6607 ( .A(n6070), .B(n6069), .Z(n6300) );
  OR U6608 ( .A(n6072), .B(n6071), .Z(n6076) );
  NANDN U6609 ( .A(n6074), .B(n6073), .Z(n6075) );
  AND U6610 ( .A(n6076), .B(n6075), .Z(n6257) );
  AND U6611 ( .A(\stack[1][25] ), .B(o[7]), .Z(n6258) );
  XNOR U6612 ( .A(n6257), .B(n6258), .Z(n6260) );
  OR U6613 ( .A(n6078), .B(n6077), .Z(n6082) );
  OR U6614 ( .A(n6080), .B(n6079), .Z(n6081) );
  AND U6615 ( .A(n6082), .B(n6081), .Z(n6263) );
  OR U6616 ( .A(n6084), .B(n6083), .Z(n6088) );
  OR U6617 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U6618 ( .A(n6088), .B(n6087), .Z(n6294) );
  NANDN U6619 ( .A(n6090), .B(n6089), .Z(n6096) );
  ANDN U6620 ( .B(\stack[1][29] ), .A(n2994), .Z(n6092) );
  NAND U6621 ( .A(n6092), .B(n6091), .Z(n6094) );
  NANDN U6622 ( .A(n2986), .B(o[2]), .Z(n6093) );
  AND U6623 ( .A(n6094), .B(n6093), .Z(n6095) );
  ANDN U6624 ( .B(n6096), .A(n6095), .Z(n6275) );
  AND U6625 ( .A(\stack[1][29] ), .B(o[3]), .Z(n6276) );
  XNOR U6626 ( .A(n6275), .B(n6276), .Z(n6278) );
  ANDN U6627 ( .B(o[0]), .A(n2989), .Z(n6098) );
  NANDN U6628 ( .A(n2995), .B(\stack[1][31] ), .Z(n6097) );
  XNOR U6629 ( .A(n6098), .B(n6097), .Z(n6282) );
  AND U6630 ( .A(\stack[1][31] ), .B(o[1]), .Z(n6283) );
  NANDN U6631 ( .A(n2994), .B(n6283), .Z(n6099) );
  XOR U6632 ( .A(n2996), .B(n6099), .Z(n6100) );
  AND U6633 ( .A(n6100), .B(\stack[1][30] ), .Z(n6281) );
  XOR U6634 ( .A(n6282), .B(n6281), .Z(n6277) );
  XOR U6635 ( .A(n6278), .B(n6277), .Z(n6293) );
  XNOR U6636 ( .A(n6294), .B(n6293), .Z(n6296) );
  AND U6637 ( .A(\stack[1][28] ), .B(o[4]), .Z(n6295) );
  XNOR U6638 ( .A(n6296), .B(n6295), .Z(n6271) );
  AND U6639 ( .A(\stack[1][27] ), .B(o[5]), .Z(n6269) );
  OR U6640 ( .A(n6102), .B(n6101), .Z(n6106) );
  NANDN U6641 ( .A(n6104), .B(n6103), .Z(n6105) );
  NAND U6642 ( .A(n6106), .B(n6105), .Z(n6270) );
  XNOR U6643 ( .A(n6269), .B(n6270), .Z(n6272) );
  XNOR U6644 ( .A(n6271), .B(n6272), .Z(n6264) );
  XNOR U6645 ( .A(n6263), .B(n6264), .Z(n6265) );
  AND U6646 ( .A(\stack[1][26] ), .B(o[6]), .Z(n6266) );
  XNOR U6647 ( .A(n6260), .B(n6259), .Z(n6299) );
  XOR U6648 ( .A(n6300), .B(n6299), .Z(n6302) );
  AND U6649 ( .A(\stack[1][24] ), .B(o[8]), .Z(n6301) );
  XNOR U6650 ( .A(n6302), .B(n6301), .Z(n6253) );
  AND U6651 ( .A(\stack[1][23] ), .B(o[9]), .Z(n6251) );
  OR U6652 ( .A(n6108), .B(n6107), .Z(n6112) );
  OR U6653 ( .A(n6110), .B(n6109), .Z(n6111) );
  NAND U6654 ( .A(n6112), .B(n6111), .Z(n6252) );
  XNOR U6655 ( .A(n6251), .B(n6252), .Z(n6254) );
  XNOR U6656 ( .A(n6253), .B(n6254), .Z(n6246) );
  XNOR U6657 ( .A(n6245), .B(n6246), .Z(n6247) );
  AND U6658 ( .A(\stack[1][22] ), .B(o[10]), .Z(n6248) );
  XNOR U6659 ( .A(n6242), .B(n6241), .Z(n6306) );
  XOR U6660 ( .A(n6305), .B(n6306), .Z(n6307) );
  XOR U6661 ( .A(n6308), .B(n6307), .Z(n6236) );
  AND U6662 ( .A(\stack[1][19] ), .B(o[13]), .Z(n6233) );
  OR U6663 ( .A(n6114), .B(n6113), .Z(n6118) );
  OR U6664 ( .A(n6116), .B(n6115), .Z(n6117) );
  NAND U6665 ( .A(n6118), .B(n6117), .Z(n6234) );
  XNOR U6666 ( .A(n6233), .B(n6234), .Z(n6235) );
  XOR U6667 ( .A(n6236), .B(n6235), .Z(n6311) );
  XNOR U6668 ( .A(n6312), .B(n6311), .Z(n6313) );
  XNOR U6669 ( .A(n6314), .B(n6313), .Z(n6229) );
  NANDN U6670 ( .A(n16826), .B(o[15]), .Z(n6227) );
  OR U6671 ( .A(n6120), .B(n6119), .Z(n6124) );
  OR U6672 ( .A(n6122), .B(n6121), .Z(n6123) );
  NAND U6673 ( .A(n6124), .B(n6123), .Z(n6228) );
  XOR U6674 ( .A(n6227), .B(n6228), .Z(n6230) );
  XNOR U6675 ( .A(n6229), .B(n6230), .Z(n6317) );
  XNOR U6676 ( .A(n6318), .B(n6317), .Z(n6320) );
  XOR U6677 ( .A(n6319), .B(n6320), .Z(n6223) );
  NANDN U6678 ( .A(n3011), .B(\stack[1][15] ), .Z(n6221) );
  OR U6679 ( .A(n6126), .B(n6125), .Z(n6130) );
  OR U6680 ( .A(n6128), .B(n6127), .Z(n6129) );
  NAND U6681 ( .A(n6130), .B(n6129), .Z(n6222) );
  XOR U6682 ( .A(n6221), .B(n6222), .Z(n6224) );
  XNOR U6683 ( .A(n6223), .B(n6224), .Z(n6323) );
  XNOR U6684 ( .A(n6324), .B(n6323), .Z(n6325) );
  XNOR U6685 ( .A(n6326), .B(n6325), .Z(n6217) );
  NANDN U6686 ( .A(n3013), .B(\stack[1][13] ), .Z(n6215) );
  OR U6687 ( .A(n6132), .B(n6131), .Z(n6136) );
  OR U6688 ( .A(n6134), .B(n6133), .Z(n6135) );
  NAND U6689 ( .A(n6136), .B(n6135), .Z(n6216) );
  XOR U6690 ( .A(n6215), .B(n6216), .Z(n6218) );
  XNOR U6691 ( .A(n6217), .B(n6218), .Z(n6329) );
  XNOR U6692 ( .A(n6330), .B(n6329), .Z(n6331) );
  XNOR U6693 ( .A(n6332), .B(n6331), .Z(n6211) );
  NANDN U6694 ( .A(n3015), .B(\stack[1][11] ), .Z(n6209) );
  OR U6695 ( .A(n6138), .B(n6137), .Z(n6142) );
  OR U6696 ( .A(n6140), .B(n6139), .Z(n6141) );
  NAND U6697 ( .A(n6142), .B(n6141), .Z(n6210) );
  XOR U6698 ( .A(n6209), .B(n6210), .Z(n6212) );
  XNOR U6699 ( .A(n6211), .B(n6212), .Z(n6335) );
  XNOR U6700 ( .A(n6336), .B(n6335), .Z(n6337) );
  XNOR U6701 ( .A(n6338), .B(n6337), .Z(n6205) );
  NANDN U6702 ( .A(n3017), .B(\stack[1][9] ), .Z(n6203) );
  OR U6703 ( .A(n6144), .B(n6143), .Z(n6148) );
  OR U6704 ( .A(n6146), .B(n6145), .Z(n6147) );
  NAND U6705 ( .A(n6148), .B(n6147), .Z(n6204) );
  XOR U6706 ( .A(n6203), .B(n6204), .Z(n6206) );
  XNOR U6707 ( .A(n6205), .B(n6206), .Z(n6341) );
  XNOR U6708 ( .A(n6342), .B(n6341), .Z(n6343) );
  XNOR U6709 ( .A(n6344), .B(n6343), .Z(n6199) );
  NANDN U6710 ( .A(n3019), .B(\stack[1][7] ), .Z(n6197) );
  OR U6711 ( .A(n6150), .B(n6149), .Z(n6154) );
  OR U6712 ( .A(n6152), .B(n6151), .Z(n6153) );
  NAND U6713 ( .A(n6154), .B(n6153), .Z(n6198) );
  XOR U6714 ( .A(n6197), .B(n6198), .Z(n6200) );
  XNOR U6715 ( .A(n6199), .B(n6200), .Z(n6347) );
  XNOR U6716 ( .A(n6348), .B(n6347), .Z(n6349) );
  XNOR U6717 ( .A(n6350), .B(n6349), .Z(n6193) );
  NANDN U6718 ( .A(n17296), .B(o[27]), .Z(n6191) );
  OR U6719 ( .A(n6156), .B(n6155), .Z(n6160) );
  OR U6720 ( .A(n6158), .B(n6157), .Z(n6159) );
  NAND U6721 ( .A(n6160), .B(n6159), .Z(n6192) );
  XOR U6722 ( .A(n6191), .B(n6192), .Z(n6194) );
  XNOR U6723 ( .A(n6193), .B(n6194), .Z(n6353) );
  XNOR U6724 ( .A(n6354), .B(n6353), .Z(n6355) );
  XNOR U6725 ( .A(n6356), .B(n6355), .Z(n6187) );
  NANDN U6726 ( .A(n17375), .B(o[29]), .Z(n6185) );
  OR U6727 ( .A(n6162), .B(n6161), .Z(n6166) );
  OR U6728 ( .A(n6164), .B(n6163), .Z(n6165) );
  NAND U6729 ( .A(n6166), .B(n6165), .Z(n6186) );
  XOR U6730 ( .A(n6185), .B(n6186), .Z(n6188) );
  XNOR U6731 ( .A(n6187), .B(n6188), .Z(n6359) );
  XNOR U6732 ( .A(n6360), .B(n6359), .Z(n6361) );
  AND U6733 ( .A(o[31]), .B(\stack[1][1] ), .Z(n6179) );
  OR U6734 ( .A(n6168), .B(n6167), .Z(n6172) );
  OR U6735 ( .A(n6170), .B(n6169), .Z(n6171) );
  NAND U6736 ( .A(n6172), .B(n6171), .Z(n6180) );
  XNOR U6737 ( .A(n6179), .B(n6180), .Z(n6182) );
  XOR U6738 ( .A(n6181), .B(n6182), .Z(n6173) );
  NANDN U6739 ( .A(n6174), .B(n6173), .Z(n6176) );
  XOR U6740 ( .A(n6174), .B(n6173), .Z(n16242) );
  AND U6741 ( .A(o[32]), .B(\stack[1][0] ), .Z(n16243) );
  OR U6742 ( .A(n16242), .B(n16243), .Z(n6175) );
  AND U6743 ( .A(n6176), .B(n6175), .Z(n6178) );
  OR U6744 ( .A(n6177), .B(n6178), .Z(n6366) );
  XNOR U6745 ( .A(n6178), .B(n6177), .Z(n16204) );
  NANDN U6746 ( .A(n2969), .B(o[32]), .Z(n6556) );
  OR U6747 ( .A(n6180), .B(n6179), .Z(n6184) );
  OR U6748 ( .A(n6182), .B(n6181), .Z(n6183) );
  NAND U6749 ( .A(n6184), .B(n6183), .Z(n6554) );
  NANDN U6750 ( .A(n17375), .B(o[30]), .Z(n6550) );
  NANDN U6751 ( .A(n6186), .B(n6185), .Z(n6190) );
  NANDN U6752 ( .A(n6188), .B(n6187), .Z(n6189) );
  NAND U6753 ( .A(n6190), .B(n6189), .Z(n6548) );
  NANDN U6754 ( .A(n17296), .B(o[28]), .Z(n6544) );
  NANDN U6755 ( .A(n6192), .B(n6191), .Z(n6196) );
  NANDN U6756 ( .A(n6194), .B(n6193), .Z(n6195) );
  NAND U6757 ( .A(n6196), .B(n6195), .Z(n6542) );
  NANDN U6758 ( .A(n17219), .B(o[26]), .Z(n6538) );
  NANDN U6759 ( .A(n6198), .B(n6197), .Z(n6202) );
  NANDN U6760 ( .A(n6200), .B(n6199), .Z(n6201) );
  NAND U6761 ( .A(n6202), .B(n6201), .Z(n6536) );
  NANDN U6762 ( .A(n17145), .B(o[24]), .Z(n6532) );
  NANDN U6763 ( .A(n6204), .B(n6203), .Z(n6208) );
  NANDN U6764 ( .A(n6206), .B(n6205), .Z(n6207) );
  NAND U6765 ( .A(n6208), .B(n6207), .Z(n6530) );
  NANDN U6766 ( .A(n2972), .B(o[22]), .Z(n6526) );
  NANDN U6767 ( .A(n6210), .B(n6209), .Z(n6214) );
  NANDN U6768 ( .A(n6212), .B(n6211), .Z(n6213) );
  NAND U6769 ( .A(n6214), .B(n6213), .Z(n6524) );
  NANDN U6770 ( .A(n2974), .B(o[20]), .Z(n6520) );
  NANDN U6771 ( .A(n6216), .B(n6215), .Z(n6220) );
  NANDN U6772 ( .A(n6218), .B(n6217), .Z(n6219) );
  NAND U6773 ( .A(n6220), .B(n6219), .Z(n6518) );
  NANDN U6774 ( .A(n2976), .B(o[18]), .Z(n6514) );
  NANDN U6775 ( .A(n6222), .B(n6221), .Z(n6226) );
  NANDN U6776 ( .A(n6224), .B(n6223), .Z(n6225) );
  NAND U6777 ( .A(n6226), .B(n6225), .Z(n6512) );
  NANDN U6778 ( .A(n3010), .B(\stack[1][17] ), .Z(n6508) );
  NANDN U6779 ( .A(n6228), .B(n6227), .Z(n6232) );
  NANDN U6780 ( .A(n6230), .B(n6229), .Z(n6231) );
  NAND U6781 ( .A(n6232), .B(n6231), .Z(n6506) );
  NANDN U6782 ( .A(n3008), .B(\stack[1][19] ), .Z(n6502) );
  OR U6783 ( .A(n6234), .B(n6233), .Z(n6238) );
  OR U6784 ( .A(n6236), .B(n6235), .Z(n6237) );
  NAND U6785 ( .A(n6238), .B(n6237), .Z(n6500) );
  NANDN U6786 ( .A(n3006), .B(\stack[1][21] ), .Z(n6430) );
  OR U6787 ( .A(n6240), .B(n6239), .Z(n6244) );
  OR U6788 ( .A(n6242), .B(n6241), .Z(n6243) );
  NAND U6789 ( .A(n6244), .B(n6243), .Z(n6428) );
  OR U6790 ( .A(n6246), .B(n6245), .Z(n6250) );
  OR U6791 ( .A(n6248), .B(n6247), .Z(n6249) );
  AND U6792 ( .A(n6250), .B(n6249), .Z(n6493) );
  AND U6793 ( .A(\stack[1][22] ), .B(o[11]), .Z(n6494) );
  XNOR U6794 ( .A(n6493), .B(n6494), .Z(n6496) );
  OR U6795 ( .A(n6252), .B(n6251), .Z(n6256) );
  OR U6796 ( .A(n6254), .B(n6253), .Z(n6255) );
  AND U6797 ( .A(n6256), .B(n6255), .Z(n6433) );
  OR U6798 ( .A(n6258), .B(n6257), .Z(n6262) );
  OR U6799 ( .A(n6260), .B(n6259), .Z(n6261) );
  NAND U6800 ( .A(n6262), .B(n6261), .Z(n6488) );
  OR U6801 ( .A(n6264), .B(n6263), .Z(n6268) );
  OR U6802 ( .A(n6266), .B(n6265), .Z(n6267) );
  AND U6803 ( .A(n6268), .B(n6267), .Z(n6445) );
  AND U6804 ( .A(\stack[1][26] ), .B(o[7]), .Z(n6446) );
  XNOR U6805 ( .A(n6445), .B(n6446), .Z(n6448) );
  OR U6806 ( .A(n6270), .B(n6269), .Z(n6274) );
  OR U6807 ( .A(n6272), .B(n6271), .Z(n6273) );
  AND U6808 ( .A(n6274), .B(n6273), .Z(n6451) );
  OR U6809 ( .A(n6276), .B(n6275), .Z(n6280) );
  OR U6810 ( .A(n6278), .B(n6277), .Z(n6279) );
  NAND U6811 ( .A(n6280), .B(n6279), .Z(n6482) );
  NANDN U6812 ( .A(n6282), .B(n6281), .Z(n6288) );
  ANDN U6813 ( .B(\stack[1][30] ), .A(n2994), .Z(n6284) );
  NAND U6814 ( .A(n6284), .B(n6283), .Z(n6286) );
  NANDN U6815 ( .A(n2987), .B(o[2]), .Z(n6285) );
  AND U6816 ( .A(n6286), .B(n6285), .Z(n6287) );
  ANDN U6817 ( .B(n6288), .A(n6287), .Z(n6463) );
  AND U6818 ( .A(\stack[1][30] ), .B(o[3]), .Z(n6464) );
  XNOR U6819 ( .A(n6463), .B(n6464), .Z(n6466) );
  ANDN U6820 ( .B(o[0]), .A(n2990), .Z(n6290) );
  NANDN U6821 ( .A(n2995), .B(\stack[1][32] ), .Z(n6289) );
  XNOR U6822 ( .A(n6290), .B(n6289), .Z(n6470) );
  AND U6823 ( .A(\stack[1][32] ), .B(o[1]), .Z(n6471) );
  NANDN U6824 ( .A(n2994), .B(n6471), .Z(n6291) );
  XOR U6825 ( .A(n2996), .B(n6291), .Z(n6292) );
  AND U6826 ( .A(n6292), .B(\stack[1][31] ), .Z(n6469) );
  XOR U6827 ( .A(n6470), .B(n6469), .Z(n6465) );
  XOR U6828 ( .A(n6466), .B(n6465), .Z(n6481) );
  XNOR U6829 ( .A(n6482), .B(n6481), .Z(n6484) );
  AND U6830 ( .A(\stack[1][29] ), .B(o[4]), .Z(n6483) );
  XNOR U6831 ( .A(n6484), .B(n6483), .Z(n6459) );
  AND U6832 ( .A(\stack[1][28] ), .B(o[5]), .Z(n6457) );
  OR U6833 ( .A(n6294), .B(n6293), .Z(n6298) );
  NANDN U6834 ( .A(n6296), .B(n6295), .Z(n6297) );
  NAND U6835 ( .A(n6298), .B(n6297), .Z(n6458) );
  XNOR U6836 ( .A(n6457), .B(n6458), .Z(n6460) );
  XNOR U6837 ( .A(n6459), .B(n6460), .Z(n6452) );
  XNOR U6838 ( .A(n6451), .B(n6452), .Z(n6453) );
  AND U6839 ( .A(\stack[1][27] ), .B(o[6]), .Z(n6454) );
  XNOR U6840 ( .A(n6448), .B(n6447), .Z(n6487) );
  XOR U6841 ( .A(n6488), .B(n6487), .Z(n6490) );
  AND U6842 ( .A(\stack[1][25] ), .B(o[8]), .Z(n6489) );
  XNOR U6843 ( .A(n6490), .B(n6489), .Z(n6441) );
  AND U6844 ( .A(\stack[1][24] ), .B(o[9]), .Z(n6439) );
  NANDN U6845 ( .A(n6300), .B(n6299), .Z(n6304) );
  NANDN U6846 ( .A(n6302), .B(n6301), .Z(n6303) );
  NAND U6847 ( .A(n6304), .B(n6303), .Z(n6440) );
  XNOR U6848 ( .A(n6439), .B(n6440), .Z(n6442) );
  XNOR U6849 ( .A(n6441), .B(n6442), .Z(n6434) );
  XOR U6850 ( .A(n6433), .B(n6434), .Z(n6435) );
  AND U6851 ( .A(\stack[1][23] ), .B(o[10]), .Z(n6436) );
  XOR U6852 ( .A(n6435), .B(n6436), .Z(n6495) );
  XOR U6853 ( .A(n6496), .B(n6495), .Z(n6427) );
  XNOR U6854 ( .A(n6428), .B(n6427), .Z(n6429) );
  XNOR U6855 ( .A(n6430), .B(n6429), .Z(n6423) );
  OR U6856 ( .A(n6306), .B(n6305), .Z(n6310) );
  NANDN U6857 ( .A(n6308), .B(n6307), .Z(n6309) );
  AND U6858 ( .A(n6310), .B(n6309), .Z(n6422) );
  NANDN U6859 ( .A(n16712), .B(o[13]), .Z(n6421) );
  XOR U6860 ( .A(n6422), .B(n6421), .Z(n6424) );
  XNOR U6861 ( .A(n6423), .B(n6424), .Z(n6499) );
  XNOR U6862 ( .A(n6500), .B(n6499), .Z(n6501) );
  XNOR U6863 ( .A(n6502), .B(n6501), .Z(n6417) );
  NANDN U6864 ( .A(n16786), .B(o[15]), .Z(n6415) );
  OR U6865 ( .A(n6312), .B(n6311), .Z(n6316) );
  OR U6866 ( .A(n6314), .B(n6313), .Z(n6315) );
  NAND U6867 ( .A(n6316), .B(n6315), .Z(n6416) );
  XOR U6868 ( .A(n6415), .B(n6416), .Z(n6418) );
  XNOR U6869 ( .A(n6417), .B(n6418), .Z(n6505) );
  XNOR U6870 ( .A(n6506), .B(n6505), .Z(n6507) );
  XNOR U6871 ( .A(n6508), .B(n6507), .Z(n6411) );
  NANDN U6872 ( .A(n3011), .B(\stack[1][16] ), .Z(n6409) );
  OR U6873 ( .A(n6318), .B(n6317), .Z(n6322) );
  IV U6874 ( .A(n6319), .Z(n16869) );
  OR U6875 ( .A(n6320), .B(n16869), .Z(n6321) );
  NAND U6876 ( .A(n6322), .B(n6321), .Z(n6410) );
  XOR U6877 ( .A(n6409), .B(n6410), .Z(n6412) );
  XNOR U6878 ( .A(n6411), .B(n6412), .Z(n6511) );
  XNOR U6879 ( .A(n6512), .B(n6511), .Z(n6513) );
  XNOR U6880 ( .A(n6514), .B(n6513), .Z(n6405) );
  NANDN U6881 ( .A(n3013), .B(\stack[1][14] ), .Z(n6403) );
  OR U6882 ( .A(n6324), .B(n6323), .Z(n6328) );
  OR U6883 ( .A(n6326), .B(n6325), .Z(n6327) );
  NAND U6884 ( .A(n6328), .B(n6327), .Z(n6404) );
  XOR U6885 ( .A(n6403), .B(n6404), .Z(n6406) );
  XNOR U6886 ( .A(n6405), .B(n6406), .Z(n6517) );
  XNOR U6887 ( .A(n6518), .B(n6517), .Z(n6519) );
  XNOR U6888 ( .A(n6520), .B(n6519), .Z(n6399) );
  NANDN U6889 ( .A(n3015), .B(\stack[1][12] ), .Z(n6397) );
  OR U6890 ( .A(n6330), .B(n6329), .Z(n6334) );
  OR U6891 ( .A(n6332), .B(n6331), .Z(n6333) );
  NAND U6892 ( .A(n6334), .B(n6333), .Z(n6398) );
  XOR U6893 ( .A(n6397), .B(n6398), .Z(n6400) );
  XNOR U6894 ( .A(n6399), .B(n6400), .Z(n6523) );
  XNOR U6895 ( .A(n6524), .B(n6523), .Z(n6525) );
  XNOR U6896 ( .A(n6526), .B(n6525), .Z(n6393) );
  NANDN U6897 ( .A(n3017), .B(\stack[1][10] ), .Z(n6391) );
  OR U6898 ( .A(n6336), .B(n6335), .Z(n6340) );
  OR U6899 ( .A(n6338), .B(n6337), .Z(n6339) );
  NAND U6900 ( .A(n6340), .B(n6339), .Z(n6392) );
  XOR U6901 ( .A(n6391), .B(n6392), .Z(n6394) );
  XNOR U6902 ( .A(n6393), .B(n6394), .Z(n6529) );
  XNOR U6903 ( .A(n6530), .B(n6529), .Z(n6531) );
  XNOR U6904 ( .A(n6532), .B(n6531), .Z(n6387) );
  NANDN U6905 ( .A(n3019), .B(\stack[1][8] ), .Z(n6385) );
  OR U6906 ( .A(n6342), .B(n6341), .Z(n6346) );
  OR U6907 ( .A(n6344), .B(n6343), .Z(n6345) );
  NAND U6908 ( .A(n6346), .B(n6345), .Z(n6386) );
  XOR U6909 ( .A(n6385), .B(n6386), .Z(n6388) );
  XNOR U6910 ( .A(n6387), .B(n6388), .Z(n6535) );
  XNOR U6911 ( .A(n6536), .B(n6535), .Z(n6537) );
  XNOR U6912 ( .A(n6538), .B(n6537), .Z(n6381) );
  NANDN U6913 ( .A(n17256), .B(o[27]), .Z(n6379) );
  OR U6914 ( .A(n6348), .B(n6347), .Z(n6352) );
  OR U6915 ( .A(n6350), .B(n6349), .Z(n6351) );
  NAND U6916 ( .A(n6352), .B(n6351), .Z(n6380) );
  XOR U6917 ( .A(n6379), .B(n6380), .Z(n6382) );
  XNOR U6918 ( .A(n6381), .B(n6382), .Z(n6541) );
  XNOR U6919 ( .A(n6542), .B(n6541), .Z(n6543) );
  XNOR U6920 ( .A(n6544), .B(n6543), .Z(n6375) );
  AND U6921 ( .A(o[29]), .B(\stack[1][4] ), .Z(n6373) );
  OR U6922 ( .A(n6354), .B(n6353), .Z(n6358) );
  OR U6923 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U6924 ( .A(n6358), .B(n6357), .Z(n6374) );
  XNOR U6925 ( .A(n6373), .B(n6374), .Z(n6376) );
  XNOR U6926 ( .A(n6375), .B(n6376), .Z(n6547) );
  XNOR U6927 ( .A(n6548), .B(n6547), .Z(n6549) );
  XOR U6928 ( .A(n6550), .B(n6549), .Z(n6370) );
  AND U6929 ( .A(o[31]), .B(\stack[1][2] ), .Z(n6367) );
  OR U6930 ( .A(n6360), .B(n6359), .Z(n6364) );
  OR U6931 ( .A(n6362), .B(n6361), .Z(n6363) );
  NAND U6932 ( .A(n6364), .B(n6363), .Z(n6368) );
  XOR U6933 ( .A(n6367), .B(n6368), .Z(n6369) );
  XNOR U6934 ( .A(n6370), .B(n6369), .Z(n6553) );
  XNOR U6935 ( .A(n6554), .B(n6553), .Z(n6555) );
  XOR U6936 ( .A(n6556), .B(n6555), .Z(n16205) );
  OR U6937 ( .A(n16204), .B(n16205), .Z(n6365) );
  AND U6938 ( .A(n6366), .B(n6365), .Z(n6560) );
  NANDN U6939 ( .A(n2970), .B(o[32]), .Z(n6759) );
  OR U6940 ( .A(n6368), .B(n6367), .Z(n6372) );
  NANDN U6941 ( .A(n6370), .B(n6369), .Z(n6371) );
  NAND U6942 ( .A(n6372), .B(n6371), .Z(n6757) );
  NANDN U6943 ( .A(n2971), .B(o[30]), .Z(n6753) );
  OR U6944 ( .A(n6374), .B(n6373), .Z(n6378) );
  NANDN U6945 ( .A(n6376), .B(n6375), .Z(n6377) );
  NAND U6946 ( .A(n6378), .B(n6377), .Z(n6751) );
  NANDN U6947 ( .A(n17256), .B(o[28]), .Z(n6747) );
  NANDN U6948 ( .A(n6380), .B(n6379), .Z(n6384) );
  NANDN U6949 ( .A(n6382), .B(n6381), .Z(n6383) );
  NAND U6950 ( .A(n6384), .B(n6383), .Z(n6745) );
  NANDN U6951 ( .A(n17179), .B(o[26]), .Z(n6741) );
  NANDN U6952 ( .A(n6386), .B(n6385), .Z(n6390) );
  NANDN U6953 ( .A(n6388), .B(n6387), .Z(n6389) );
  NAND U6954 ( .A(n6390), .B(n6389), .Z(n6739) );
  NANDN U6955 ( .A(n17101), .B(o[24]), .Z(n6735) );
  NANDN U6956 ( .A(n6392), .B(n6391), .Z(n6396) );
  NANDN U6957 ( .A(n6394), .B(n6393), .Z(n6395) );
  NAND U6958 ( .A(n6396), .B(n6395), .Z(n6733) );
  NANDN U6959 ( .A(n2973), .B(o[22]), .Z(n6729) );
  NANDN U6960 ( .A(n6398), .B(n6397), .Z(n6402) );
  NANDN U6961 ( .A(n6400), .B(n6399), .Z(n6401) );
  NAND U6962 ( .A(n6402), .B(n6401), .Z(n6727) );
  NANDN U6963 ( .A(n2975), .B(o[20]), .Z(n6723) );
  NANDN U6964 ( .A(n6404), .B(n6403), .Z(n6408) );
  NANDN U6965 ( .A(n6406), .B(n6405), .Z(n6407) );
  NAND U6966 ( .A(n6408), .B(n6407), .Z(n6721) );
  NANDN U6967 ( .A(n2977), .B(o[18]), .Z(n6717) );
  NANDN U6968 ( .A(n6410), .B(n6409), .Z(n6414) );
  NANDN U6969 ( .A(n6412), .B(n6411), .Z(n6413) );
  NAND U6970 ( .A(n6414), .B(n6413), .Z(n6715) );
  NANDN U6971 ( .A(n3010), .B(\stack[1][18] ), .Z(n6711) );
  NANDN U6972 ( .A(n6416), .B(n6415), .Z(n6420) );
  NANDN U6973 ( .A(n6418), .B(n6417), .Z(n6419) );
  NAND U6974 ( .A(n6420), .B(n6419), .Z(n6709) );
  NANDN U6975 ( .A(n3008), .B(\stack[1][20] ), .Z(n6705) );
  NANDN U6976 ( .A(n6422), .B(n6421), .Z(n6426) );
  NANDN U6977 ( .A(n6424), .B(n6423), .Z(n6425) );
  NAND U6978 ( .A(n6426), .B(n6425), .Z(n6703) );
  AND U6979 ( .A(\stack[1][21] ), .B(o[13]), .Z(n6624) );
  OR U6980 ( .A(n6428), .B(n6427), .Z(n6432) );
  OR U6981 ( .A(n6430), .B(n6429), .Z(n6431) );
  NAND U6982 ( .A(n6432), .B(n6431), .Z(n6625) );
  XNOR U6983 ( .A(n6624), .B(n6625), .Z(n6627) );
  OR U6984 ( .A(n6434), .B(n6433), .Z(n6438) );
  NANDN U6985 ( .A(n6436), .B(n6435), .Z(n6437) );
  NAND U6986 ( .A(n6438), .B(n6437), .Z(n6631) );
  ANDN U6987 ( .B(o[11]), .A(n2980), .Z(n6630) );
  XOR U6988 ( .A(n6631), .B(n6630), .Z(n6632) );
  NANDN U6989 ( .A(n3004), .B(\stack[1][24] ), .Z(n6639) );
  OR U6990 ( .A(n6440), .B(n6439), .Z(n6444) );
  OR U6991 ( .A(n6442), .B(n6441), .Z(n6443) );
  NAND U6992 ( .A(n6444), .B(n6443), .Z(n6637) );
  NANDN U6993 ( .A(n3002), .B(\stack[1][26] ), .Z(n6693) );
  OR U6994 ( .A(n6446), .B(n6445), .Z(n6450) );
  OR U6995 ( .A(n6448), .B(n6447), .Z(n6449) );
  NAND U6996 ( .A(n6450), .B(n6449), .Z(n6691) );
  OR U6997 ( .A(n6452), .B(n6451), .Z(n6456) );
  OR U6998 ( .A(n6454), .B(n6453), .Z(n6455) );
  AND U6999 ( .A(n6456), .B(n6455), .Z(n6648) );
  AND U7000 ( .A(\stack[1][27] ), .B(o[7]), .Z(n6649) );
  XNOR U7001 ( .A(n6648), .B(n6649), .Z(n6651) );
  OR U7002 ( .A(n6458), .B(n6457), .Z(n6462) );
  OR U7003 ( .A(n6460), .B(n6459), .Z(n6461) );
  AND U7004 ( .A(n6462), .B(n6461), .Z(n6654) );
  OR U7005 ( .A(n6464), .B(n6463), .Z(n6468) );
  OR U7006 ( .A(n6466), .B(n6465), .Z(n6467) );
  NAND U7007 ( .A(n6468), .B(n6467), .Z(n6685) );
  NANDN U7008 ( .A(n6470), .B(n6469), .Z(n6476) );
  ANDN U7009 ( .B(\stack[1][31] ), .A(n2994), .Z(n6472) );
  NAND U7010 ( .A(n6472), .B(n6471), .Z(n6474) );
  NANDN U7011 ( .A(n2988), .B(o[2]), .Z(n6473) );
  AND U7012 ( .A(n6474), .B(n6473), .Z(n6475) );
  ANDN U7013 ( .B(n6476), .A(n6475), .Z(n6666) );
  AND U7014 ( .A(\stack[1][31] ), .B(o[3]), .Z(n6667) );
  XNOR U7015 ( .A(n6666), .B(n6667), .Z(n6669) );
  ANDN U7016 ( .B(o[0]), .A(n2991), .Z(n6478) );
  NANDN U7017 ( .A(n2995), .B(\stack[1][33] ), .Z(n6477) );
  XNOR U7018 ( .A(n6478), .B(n6477), .Z(n6673) );
  AND U7019 ( .A(\stack[1][33] ), .B(o[1]), .Z(n6674) );
  NANDN U7020 ( .A(n2994), .B(n6674), .Z(n6479) );
  XOR U7021 ( .A(n2996), .B(n6479), .Z(n6480) );
  AND U7022 ( .A(n6480), .B(\stack[1][32] ), .Z(n6672) );
  XOR U7023 ( .A(n6673), .B(n6672), .Z(n6668) );
  XOR U7024 ( .A(n6669), .B(n6668), .Z(n6684) );
  XNOR U7025 ( .A(n6685), .B(n6684), .Z(n6687) );
  AND U7026 ( .A(\stack[1][30] ), .B(o[4]), .Z(n6686) );
  XNOR U7027 ( .A(n6687), .B(n6686), .Z(n6662) );
  AND U7028 ( .A(\stack[1][29] ), .B(o[5]), .Z(n6660) );
  OR U7029 ( .A(n6482), .B(n6481), .Z(n6486) );
  NANDN U7030 ( .A(n6484), .B(n6483), .Z(n6485) );
  NAND U7031 ( .A(n6486), .B(n6485), .Z(n6661) );
  XNOR U7032 ( .A(n6660), .B(n6661), .Z(n6663) );
  XNOR U7033 ( .A(n6662), .B(n6663), .Z(n6655) );
  XOR U7034 ( .A(n6654), .B(n6655), .Z(n6656) );
  AND U7035 ( .A(\stack[1][28] ), .B(o[6]), .Z(n6657) );
  XOR U7036 ( .A(n6656), .B(n6657), .Z(n6650) );
  XOR U7037 ( .A(n6651), .B(n6650), .Z(n6690) );
  XNOR U7038 ( .A(n6691), .B(n6690), .Z(n6692) );
  XNOR U7039 ( .A(n6693), .B(n6692), .Z(n6644) );
  AND U7040 ( .A(\stack[1][25] ), .B(o[9]), .Z(n6642) );
  NANDN U7041 ( .A(n6488), .B(n6487), .Z(n6492) );
  NANDN U7042 ( .A(n6490), .B(n6489), .Z(n6491) );
  NAND U7043 ( .A(n6492), .B(n6491), .Z(n6643) );
  XNOR U7044 ( .A(n6642), .B(n6643), .Z(n6645) );
  XNOR U7045 ( .A(n6644), .B(n6645), .Z(n6636) );
  XNOR U7046 ( .A(n6637), .B(n6636), .Z(n6638) );
  XNOR U7047 ( .A(n6639), .B(n6638), .Z(n6633) );
  OR U7048 ( .A(n6494), .B(n6493), .Z(n6498) );
  OR U7049 ( .A(n6496), .B(n6495), .Z(n6497) );
  AND U7050 ( .A(n6498), .B(n6497), .Z(n6697) );
  XNOR U7051 ( .A(n6696), .B(n6697), .Z(n6699) );
  AND U7052 ( .A(\stack[1][22] ), .B(o[12]), .Z(n6698) );
  XNOR U7053 ( .A(n6699), .B(n6698), .Z(n6626) );
  XOR U7054 ( .A(n6627), .B(n6626), .Z(n6702) );
  XNOR U7055 ( .A(n6703), .B(n6702), .Z(n6704) );
  XNOR U7056 ( .A(n6705), .B(n6704), .Z(n6620) );
  NANDN U7057 ( .A(n16746), .B(o[15]), .Z(n6618) );
  OR U7058 ( .A(n6500), .B(n6499), .Z(n6504) );
  OR U7059 ( .A(n6502), .B(n6501), .Z(n6503) );
  NAND U7060 ( .A(n6504), .B(n6503), .Z(n6619) );
  XOR U7061 ( .A(n6618), .B(n6619), .Z(n6621) );
  XNOR U7062 ( .A(n6620), .B(n6621), .Z(n6708) );
  XNOR U7063 ( .A(n6709), .B(n6708), .Z(n6710) );
  XNOR U7064 ( .A(n6711), .B(n6710), .Z(n6614) );
  AND U7065 ( .A(o[17]), .B(\stack[1][17] ), .Z(n16827) );
  OR U7066 ( .A(n6506), .B(n6505), .Z(n6510) );
  OR U7067 ( .A(n6508), .B(n6507), .Z(n6509) );
  NAND U7068 ( .A(n6510), .B(n6509), .Z(n6613) );
  XNOR U7069 ( .A(n16827), .B(n6613), .Z(n6615) );
  XNOR U7070 ( .A(n6614), .B(n6615), .Z(n6714) );
  XNOR U7071 ( .A(n6715), .B(n6714), .Z(n6716) );
  XNOR U7072 ( .A(n6717), .B(n6716), .Z(n6609) );
  NANDN U7073 ( .A(n3013), .B(\stack[1][15] ), .Z(n6607) );
  OR U7074 ( .A(n6512), .B(n6511), .Z(n6516) );
  OR U7075 ( .A(n6514), .B(n6513), .Z(n6515) );
  NAND U7076 ( .A(n6516), .B(n6515), .Z(n6608) );
  XOR U7077 ( .A(n6607), .B(n6608), .Z(n6610) );
  XNOR U7078 ( .A(n6609), .B(n6610), .Z(n6720) );
  XNOR U7079 ( .A(n6721), .B(n6720), .Z(n6722) );
  XNOR U7080 ( .A(n6723), .B(n6722), .Z(n6603) );
  NANDN U7081 ( .A(n3015), .B(\stack[1][13] ), .Z(n6601) );
  OR U7082 ( .A(n6518), .B(n6517), .Z(n6522) );
  OR U7083 ( .A(n6520), .B(n6519), .Z(n6521) );
  NAND U7084 ( .A(n6522), .B(n6521), .Z(n6602) );
  XOR U7085 ( .A(n6601), .B(n6602), .Z(n6604) );
  XNOR U7086 ( .A(n6603), .B(n6604), .Z(n6726) );
  XNOR U7087 ( .A(n6727), .B(n6726), .Z(n6728) );
  XNOR U7088 ( .A(n6729), .B(n6728), .Z(n6597) );
  NANDN U7089 ( .A(n3017), .B(\stack[1][11] ), .Z(n6595) );
  OR U7090 ( .A(n6524), .B(n6523), .Z(n6528) );
  OR U7091 ( .A(n6526), .B(n6525), .Z(n6527) );
  NAND U7092 ( .A(n6528), .B(n6527), .Z(n6596) );
  XOR U7093 ( .A(n6595), .B(n6596), .Z(n6598) );
  XNOR U7094 ( .A(n6597), .B(n6598), .Z(n6732) );
  XNOR U7095 ( .A(n6733), .B(n6732), .Z(n6734) );
  XNOR U7096 ( .A(n6735), .B(n6734), .Z(n6591) );
  NANDN U7097 ( .A(n3019), .B(\stack[1][9] ), .Z(n6589) );
  OR U7098 ( .A(n6530), .B(n6529), .Z(n6534) );
  OR U7099 ( .A(n6532), .B(n6531), .Z(n6533) );
  NAND U7100 ( .A(n6534), .B(n6533), .Z(n6590) );
  XOR U7101 ( .A(n6589), .B(n6590), .Z(n6592) );
  XNOR U7102 ( .A(n6591), .B(n6592), .Z(n6738) );
  XNOR U7103 ( .A(n6739), .B(n6738), .Z(n6740) );
  XNOR U7104 ( .A(n6741), .B(n6740), .Z(n6585) );
  NANDN U7105 ( .A(n17219), .B(o[27]), .Z(n6583) );
  OR U7106 ( .A(n6536), .B(n6535), .Z(n6540) );
  OR U7107 ( .A(n6538), .B(n6537), .Z(n6539) );
  NAND U7108 ( .A(n6540), .B(n6539), .Z(n6584) );
  XOR U7109 ( .A(n6583), .B(n6584), .Z(n6586) );
  XNOR U7110 ( .A(n6585), .B(n6586), .Z(n6744) );
  XNOR U7111 ( .A(n6745), .B(n6744), .Z(n6746) );
  XNOR U7112 ( .A(n6747), .B(n6746), .Z(n6579) );
  NANDN U7113 ( .A(n17296), .B(o[29]), .Z(n6577) );
  OR U7114 ( .A(n6542), .B(n6541), .Z(n6546) );
  OR U7115 ( .A(n6544), .B(n6543), .Z(n6545) );
  NAND U7116 ( .A(n6546), .B(n6545), .Z(n6578) );
  XOR U7117 ( .A(n6577), .B(n6578), .Z(n6580) );
  XNOR U7118 ( .A(n6579), .B(n6580), .Z(n6750) );
  XNOR U7119 ( .A(n6751), .B(n6750), .Z(n6752) );
  XNOR U7120 ( .A(n6753), .B(n6752), .Z(n6573) );
  NANDN U7121 ( .A(n17375), .B(o[31]), .Z(n6571) );
  OR U7122 ( .A(n6548), .B(n6547), .Z(n6552) );
  OR U7123 ( .A(n6550), .B(n6549), .Z(n6551) );
  NAND U7124 ( .A(n6552), .B(n6551), .Z(n6572) );
  XOR U7125 ( .A(n6571), .B(n6572), .Z(n6574) );
  XNOR U7126 ( .A(n6573), .B(n6574), .Z(n6756) );
  XNOR U7127 ( .A(n6757), .B(n6756), .Z(n6758) );
  AND U7128 ( .A(o[33]), .B(\stack[1][1] ), .Z(n6565) );
  OR U7129 ( .A(n6554), .B(n6553), .Z(n6558) );
  OR U7130 ( .A(n6556), .B(n6555), .Z(n6557) );
  NAND U7131 ( .A(n6558), .B(n6557), .Z(n6566) );
  XNOR U7132 ( .A(n6565), .B(n6566), .Z(n6568) );
  XOR U7133 ( .A(n6567), .B(n6568), .Z(n6559) );
  NANDN U7134 ( .A(n6560), .B(n6559), .Z(n6562) );
  XOR U7135 ( .A(n6560), .B(n6559), .Z(n16166) );
  AND U7136 ( .A(o[34]), .B(\stack[1][0] ), .Z(n16167) );
  OR U7137 ( .A(n16166), .B(n16167), .Z(n6561) );
  AND U7138 ( .A(n6562), .B(n6561), .Z(n6564) );
  OR U7139 ( .A(n6563), .B(n6564), .Z(n6763) );
  XNOR U7140 ( .A(n6564), .B(n6563), .Z(n16128) );
  NANDN U7141 ( .A(n2969), .B(o[34]), .Z(n6965) );
  OR U7142 ( .A(n6566), .B(n6565), .Z(n6570) );
  OR U7143 ( .A(n6568), .B(n6567), .Z(n6569) );
  NAND U7144 ( .A(n6570), .B(n6569), .Z(n6963) );
  NANDN U7145 ( .A(n17375), .B(o[32]), .Z(n6959) );
  NANDN U7146 ( .A(n6572), .B(n6571), .Z(n6576) );
  NANDN U7147 ( .A(n6574), .B(n6573), .Z(n6575) );
  NAND U7148 ( .A(n6576), .B(n6575), .Z(n6957) );
  NANDN U7149 ( .A(n17296), .B(o[30]), .Z(n6953) );
  NANDN U7150 ( .A(n6578), .B(n6577), .Z(n6582) );
  NANDN U7151 ( .A(n6580), .B(n6579), .Z(n6581) );
  NAND U7152 ( .A(n6582), .B(n6581), .Z(n6951) );
  NANDN U7153 ( .A(n17219), .B(o[28]), .Z(n6947) );
  NANDN U7154 ( .A(n6584), .B(n6583), .Z(n6588) );
  NANDN U7155 ( .A(n6586), .B(n6585), .Z(n6587) );
  NAND U7156 ( .A(n6588), .B(n6587), .Z(n6945) );
  NANDN U7157 ( .A(n17145), .B(o[26]), .Z(n6941) );
  NANDN U7158 ( .A(n6590), .B(n6589), .Z(n6594) );
  NANDN U7159 ( .A(n6592), .B(n6591), .Z(n6593) );
  NAND U7160 ( .A(n6594), .B(n6593), .Z(n6939) );
  NANDN U7161 ( .A(n2972), .B(o[24]), .Z(n6935) );
  NANDN U7162 ( .A(n6596), .B(n6595), .Z(n6600) );
  NANDN U7163 ( .A(n6598), .B(n6597), .Z(n6599) );
  NAND U7164 ( .A(n6600), .B(n6599), .Z(n6933) );
  NANDN U7165 ( .A(n2974), .B(o[22]), .Z(n6929) );
  NANDN U7166 ( .A(n6602), .B(n6601), .Z(n6606) );
  NANDN U7167 ( .A(n6604), .B(n6603), .Z(n6605) );
  NAND U7168 ( .A(n6606), .B(n6605), .Z(n6927) );
  NANDN U7169 ( .A(n2976), .B(o[20]), .Z(n6923) );
  NANDN U7170 ( .A(n6608), .B(n6607), .Z(n6612) );
  NANDN U7171 ( .A(n6610), .B(n6609), .Z(n6611) );
  NAND U7172 ( .A(n6612), .B(n6611), .Z(n6921) );
  NANDN U7173 ( .A(n16826), .B(o[18]), .Z(n6917) );
  OR U7174 ( .A(n6613), .B(n16827), .Z(n6617) );
  NANDN U7175 ( .A(n6615), .B(n6614), .Z(n6616) );
  NAND U7176 ( .A(n6617), .B(n6616), .Z(n6915) );
  NANDN U7177 ( .A(n3010), .B(\stack[1][19] ), .Z(n6911) );
  NANDN U7178 ( .A(n6619), .B(n6618), .Z(n6623) );
  NANDN U7179 ( .A(n6621), .B(n6620), .Z(n6622) );
  NAND U7180 ( .A(n6623), .B(n6622), .Z(n6909) );
  NANDN U7181 ( .A(n3008), .B(\stack[1][21] ), .Z(n6905) );
  OR U7182 ( .A(n6625), .B(n6624), .Z(n6629) );
  OR U7183 ( .A(n6627), .B(n6626), .Z(n6628) );
  NAND U7184 ( .A(n6629), .B(n6628), .Z(n6903) );
  NANDN U7185 ( .A(n3006), .B(\stack[1][23] ), .Z(n6833) );
  NANDN U7186 ( .A(n6631), .B(n6630), .Z(n6635) );
  OR U7187 ( .A(n6633), .B(n6632), .Z(n6634) );
  AND U7188 ( .A(n6635), .B(n6634), .Z(n6830) );
  AND U7189 ( .A(\stack[1][24] ), .B(o[11]), .Z(n6896) );
  OR U7190 ( .A(n6637), .B(n6636), .Z(n6641) );
  OR U7191 ( .A(n6639), .B(n6638), .Z(n6640) );
  NAND U7192 ( .A(n6641), .B(n6640), .Z(n6897) );
  XNOR U7193 ( .A(n6896), .B(n6897), .Z(n6899) );
  OR U7194 ( .A(n6643), .B(n6642), .Z(n6647) );
  NANDN U7195 ( .A(n6645), .B(n6644), .Z(n6646) );
  AND U7196 ( .A(n6647), .B(n6646), .Z(n6836) );
  OR U7197 ( .A(n6649), .B(n6648), .Z(n6653) );
  OR U7198 ( .A(n6651), .B(n6650), .Z(n6652) );
  NAND U7199 ( .A(n6653), .B(n6652), .Z(n6891) );
  OR U7200 ( .A(n6655), .B(n6654), .Z(n6659) );
  NANDN U7201 ( .A(n6657), .B(n6656), .Z(n6658) );
  AND U7202 ( .A(n6659), .B(n6658), .Z(n6848) );
  AND U7203 ( .A(\stack[1][28] ), .B(o[7]), .Z(n6849) );
  XNOR U7204 ( .A(n6848), .B(n6849), .Z(n6851) );
  OR U7205 ( .A(n6661), .B(n6660), .Z(n6665) );
  OR U7206 ( .A(n6663), .B(n6662), .Z(n6664) );
  AND U7207 ( .A(n6665), .B(n6664), .Z(n6854) );
  OR U7208 ( .A(n6667), .B(n6666), .Z(n6671) );
  OR U7209 ( .A(n6669), .B(n6668), .Z(n6670) );
  NAND U7210 ( .A(n6671), .B(n6670), .Z(n6885) );
  NANDN U7211 ( .A(n6673), .B(n6672), .Z(n6679) );
  ANDN U7212 ( .B(\stack[1][32] ), .A(n2994), .Z(n6675) );
  NAND U7213 ( .A(n6675), .B(n6674), .Z(n6677) );
  NANDN U7214 ( .A(n2989), .B(o[2]), .Z(n6676) );
  AND U7215 ( .A(n6677), .B(n6676), .Z(n6678) );
  ANDN U7216 ( .B(n6679), .A(n6678), .Z(n6866) );
  AND U7217 ( .A(\stack[1][32] ), .B(o[3]), .Z(n6867) );
  XNOR U7218 ( .A(n6866), .B(n6867), .Z(n6869) );
  ANDN U7219 ( .B(o[0]), .A(n2992), .Z(n6681) );
  NANDN U7220 ( .A(n2995), .B(\stack[1][34] ), .Z(n6680) );
  XNOR U7221 ( .A(n6681), .B(n6680), .Z(n6873) );
  AND U7222 ( .A(\stack[1][34] ), .B(o[1]), .Z(n6874) );
  NANDN U7223 ( .A(n2994), .B(n6874), .Z(n6682) );
  XOR U7224 ( .A(n2996), .B(n6682), .Z(n6683) );
  AND U7225 ( .A(n6683), .B(\stack[1][33] ), .Z(n6872) );
  XOR U7226 ( .A(n6873), .B(n6872), .Z(n6868) );
  XOR U7227 ( .A(n6869), .B(n6868), .Z(n6884) );
  XNOR U7228 ( .A(n6885), .B(n6884), .Z(n6887) );
  AND U7229 ( .A(\stack[1][31] ), .B(o[4]), .Z(n6886) );
  XNOR U7230 ( .A(n6887), .B(n6886), .Z(n6862) );
  AND U7231 ( .A(\stack[1][30] ), .B(o[5]), .Z(n6860) );
  OR U7232 ( .A(n6685), .B(n6684), .Z(n6689) );
  NANDN U7233 ( .A(n6687), .B(n6686), .Z(n6688) );
  NAND U7234 ( .A(n6689), .B(n6688), .Z(n6861) );
  XNOR U7235 ( .A(n6860), .B(n6861), .Z(n6863) );
  XNOR U7236 ( .A(n6862), .B(n6863), .Z(n6855) );
  XNOR U7237 ( .A(n6854), .B(n6855), .Z(n6856) );
  AND U7238 ( .A(\stack[1][29] ), .B(o[6]), .Z(n6857) );
  XNOR U7239 ( .A(n6851), .B(n6850), .Z(n6890) );
  XOR U7240 ( .A(n6891), .B(n6890), .Z(n6893) );
  AND U7241 ( .A(\stack[1][27] ), .B(o[8]), .Z(n6892) );
  XNOR U7242 ( .A(n6893), .B(n6892), .Z(n6844) );
  AND U7243 ( .A(\stack[1][26] ), .B(o[9]), .Z(n6842) );
  OR U7244 ( .A(n6691), .B(n6690), .Z(n6695) );
  OR U7245 ( .A(n6693), .B(n6692), .Z(n6694) );
  NAND U7246 ( .A(n6695), .B(n6694), .Z(n6843) );
  XNOR U7247 ( .A(n6842), .B(n6843), .Z(n6845) );
  XNOR U7248 ( .A(n6844), .B(n6845), .Z(n6837) );
  XNOR U7249 ( .A(n6836), .B(n6837), .Z(n6838) );
  AND U7250 ( .A(\stack[1][25] ), .B(o[10]), .Z(n6839) );
  XOR U7251 ( .A(n6899), .B(n6898), .Z(n6831) );
  XNOR U7252 ( .A(n6830), .B(n6831), .Z(n6832) );
  XNOR U7253 ( .A(n6833), .B(n6832), .Z(n6826) );
  OR U7254 ( .A(n6697), .B(n6696), .Z(n6701) );
  OR U7255 ( .A(n6699), .B(n6698), .Z(n6700) );
  AND U7256 ( .A(n6701), .B(n6700), .Z(n6825) );
  NANDN U7257 ( .A(n2979), .B(o[13]), .Z(n6824) );
  XOR U7258 ( .A(n6825), .B(n6824), .Z(n6827) );
  XNOR U7259 ( .A(n6826), .B(n6827), .Z(n6902) );
  XNOR U7260 ( .A(n6903), .B(n6902), .Z(n6904) );
  XNOR U7261 ( .A(n6905), .B(n6904), .Z(n6820) );
  NANDN U7262 ( .A(n16712), .B(o[15]), .Z(n6818) );
  OR U7263 ( .A(n6703), .B(n6702), .Z(n6707) );
  OR U7264 ( .A(n6705), .B(n6704), .Z(n6706) );
  NAND U7265 ( .A(n6707), .B(n6706), .Z(n6819) );
  XOR U7266 ( .A(n6818), .B(n6819), .Z(n6821) );
  XNOR U7267 ( .A(n6820), .B(n6821), .Z(n6908) );
  XNOR U7268 ( .A(n6909), .B(n6908), .Z(n6910) );
  XNOR U7269 ( .A(n6911), .B(n6910), .Z(n6814) );
  NANDN U7270 ( .A(n16786), .B(o[17]), .Z(n6812) );
  OR U7271 ( .A(n6709), .B(n6708), .Z(n6713) );
  OR U7272 ( .A(n6711), .B(n6710), .Z(n6712) );
  NAND U7273 ( .A(n6713), .B(n6712), .Z(n6813) );
  XOR U7274 ( .A(n6812), .B(n6813), .Z(n6815) );
  XNOR U7275 ( .A(n6814), .B(n6815), .Z(n6914) );
  XNOR U7276 ( .A(n6915), .B(n6914), .Z(n6916) );
  XNOR U7277 ( .A(n6917), .B(n6916), .Z(n6808) );
  NANDN U7278 ( .A(n3013), .B(\stack[1][16] ), .Z(n6806) );
  OR U7279 ( .A(n6715), .B(n6714), .Z(n6719) );
  OR U7280 ( .A(n6717), .B(n6716), .Z(n6718) );
  NAND U7281 ( .A(n6719), .B(n6718), .Z(n6807) );
  XOR U7282 ( .A(n6806), .B(n6807), .Z(n6809) );
  XNOR U7283 ( .A(n6808), .B(n6809), .Z(n6920) );
  XNOR U7284 ( .A(n6921), .B(n6920), .Z(n6922) );
  XNOR U7285 ( .A(n6923), .B(n6922), .Z(n6802) );
  NANDN U7286 ( .A(n3015), .B(\stack[1][14] ), .Z(n6800) );
  OR U7287 ( .A(n6721), .B(n6720), .Z(n6725) );
  OR U7288 ( .A(n6723), .B(n6722), .Z(n6724) );
  NAND U7289 ( .A(n6725), .B(n6724), .Z(n6801) );
  XOR U7290 ( .A(n6800), .B(n6801), .Z(n6803) );
  XNOR U7291 ( .A(n6802), .B(n6803), .Z(n6926) );
  XNOR U7292 ( .A(n6927), .B(n6926), .Z(n6928) );
  XNOR U7293 ( .A(n6929), .B(n6928), .Z(n6796) );
  NANDN U7294 ( .A(n3017), .B(\stack[1][12] ), .Z(n6794) );
  OR U7295 ( .A(n6727), .B(n6726), .Z(n6731) );
  OR U7296 ( .A(n6729), .B(n6728), .Z(n6730) );
  NAND U7297 ( .A(n6731), .B(n6730), .Z(n6795) );
  XOR U7298 ( .A(n6794), .B(n6795), .Z(n6797) );
  XNOR U7299 ( .A(n6796), .B(n6797), .Z(n6932) );
  XNOR U7300 ( .A(n6933), .B(n6932), .Z(n6934) );
  XNOR U7301 ( .A(n6935), .B(n6934), .Z(n6790) );
  NANDN U7302 ( .A(n3019), .B(\stack[1][10] ), .Z(n6788) );
  OR U7303 ( .A(n6733), .B(n6732), .Z(n6737) );
  OR U7304 ( .A(n6735), .B(n6734), .Z(n6736) );
  NAND U7305 ( .A(n6737), .B(n6736), .Z(n6789) );
  XOR U7306 ( .A(n6788), .B(n6789), .Z(n6791) );
  XNOR U7307 ( .A(n6790), .B(n6791), .Z(n6938) );
  XNOR U7308 ( .A(n6939), .B(n6938), .Z(n6940) );
  XNOR U7309 ( .A(n6941), .B(n6940), .Z(n6784) );
  NANDN U7310 ( .A(n17179), .B(o[27]), .Z(n6782) );
  OR U7311 ( .A(n6739), .B(n6738), .Z(n6743) );
  OR U7312 ( .A(n6741), .B(n6740), .Z(n6742) );
  NAND U7313 ( .A(n6743), .B(n6742), .Z(n6783) );
  XOR U7314 ( .A(n6782), .B(n6783), .Z(n6785) );
  XNOR U7315 ( .A(n6784), .B(n6785), .Z(n6944) );
  XNOR U7316 ( .A(n6945), .B(n6944), .Z(n6946) );
  XNOR U7317 ( .A(n6947), .B(n6946), .Z(n6778) );
  NANDN U7318 ( .A(n17256), .B(o[29]), .Z(n6776) );
  OR U7319 ( .A(n6745), .B(n6744), .Z(n6749) );
  OR U7320 ( .A(n6747), .B(n6746), .Z(n6748) );
  NAND U7321 ( .A(n6749), .B(n6748), .Z(n6777) );
  XOR U7322 ( .A(n6776), .B(n6777), .Z(n6779) );
  XNOR U7323 ( .A(n6778), .B(n6779), .Z(n6950) );
  XNOR U7324 ( .A(n6951), .B(n6950), .Z(n6952) );
  XNOR U7325 ( .A(n6953), .B(n6952), .Z(n6772) );
  AND U7326 ( .A(o[31]), .B(\stack[1][4] ), .Z(n6770) );
  OR U7327 ( .A(n6751), .B(n6750), .Z(n6755) );
  OR U7328 ( .A(n6753), .B(n6752), .Z(n6754) );
  NAND U7329 ( .A(n6755), .B(n6754), .Z(n6771) );
  XNOR U7330 ( .A(n6770), .B(n6771), .Z(n6773) );
  XNOR U7331 ( .A(n6772), .B(n6773), .Z(n6956) );
  XNOR U7332 ( .A(n6957), .B(n6956), .Z(n6958) );
  XOR U7333 ( .A(n6959), .B(n6958), .Z(n6767) );
  AND U7334 ( .A(o[33]), .B(\stack[1][2] ), .Z(n6764) );
  OR U7335 ( .A(n6757), .B(n6756), .Z(n6761) );
  OR U7336 ( .A(n6759), .B(n6758), .Z(n6760) );
  NAND U7337 ( .A(n6761), .B(n6760), .Z(n6765) );
  XOR U7338 ( .A(n6764), .B(n6765), .Z(n6766) );
  XNOR U7339 ( .A(n6767), .B(n6766), .Z(n6962) );
  XNOR U7340 ( .A(n6963), .B(n6962), .Z(n6964) );
  XOR U7341 ( .A(n6965), .B(n6964), .Z(n16129) );
  OR U7342 ( .A(n16128), .B(n16129), .Z(n6762) );
  AND U7343 ( .A(n6763), .B(n6762), .Z(n6969) );
  NANDN U7344 ( .A(n2970), .B(o[34]), .Z(n7180) );
  OR U7345 ( .A(n6765), .B(n6764), .Z(n6769) );
  NANDN U7346 ( .A(n6767), .B(n6766), .Z(n6768) );
  NAND U7347 ( .A(n6769), .B(n6768), .Z(n7178) );
  NANDN U7348 ( .A(n2971), .B(o[32]), .Z(n7174) );
  OR U7349 ( .A(n6771), .B(n6770), .Z(n6775) );
  NANDN U7350 ( .A(n6773), .B(n6772), .Z(n6774) );
  NAND U7351 ( .A(n6775), .B(n6774), .Z(n7172) );
  NANDN U7352 ( .A(n17256), .B(o[30]), .Z(n7168) );
  NANDN U7353 ( .A(n6777), .B(n6776), .Z(n6781) );
  NANDN U7354 ( .A(n6779), .B(n6778), .Z(n6780) );
  NAND U7355 ( .A(n6781), .B(n6780), .Z(n7166) );
  NANDN U7356 ( .A(n17179), .B(o[28]), .Z(n7162) );
  NANDN U7357 ( .A(n6783), .B(n6782), .Z(n6787) );
  NANDN U7358 ( .A(n6785), .B(n6784), .Z(n6786) );
  NAND U7359 ( .A(n6787), .B(n6786), .Z(n7160) );
  NANDN U7360 ( .A(n17101), .B(o[26]), .Z(n7156) );
  NANDN U7361 ( .A(n6789), .B(n6788), .Z(n6793) );
  NANDN U7362 ( .A(n6791), .B(n6790), .Z(n6792) );
  NAND U7363 ( .A(n6793), .B(n6792), .Z(n7154) );
  NANDN U7364 ( .A(n2973), .B(o[24]), .Z(n7150) );
  NANDN U7365 ( .A(n6795), .B(n6794), .Z(n6799) );
  NANDN U7366 ( .A(n6797), .B(n6796), .Z(n6798) );
  NAND U7367 ( .A(n6799), .B(n6798), .Z(n7148) );
  NANDN U7368 ( .A(n2975), .B(o[22]), .Z(n7144) );
  NANDN U7369 ( .A(n6801), .B(n6800), .Z(n6805) );
  NANDN U7370 ( .A(n6803), .B(n6802), .Z(n6804) );
  NAND U7371 ( .A(n6805), .B(n6804), .Z(n7142) );
  NANDN U7372 ( .A(n2977), .B(o[20]), .Z(n7138) );
  NANDN U7373 ( .A(n6807), .B(n6806), .Z(n6811) );
  NANDN U7374 ( .A(n6809), .B(n6808), .Z(n6810) );
  NAND U7375 ( .A(n6811), .B(n6810), .Z(n7136) );
  NOR U7376 ( .A(n3012), .B(n16786), .Z(n7131) );
  NANDN U7377 ( .A(n6813), .B(n6812), .Z(n6817) );
  NANDN U7378 ( .A(n6815), .B(n6814), .Z(n6816) );
  NAND U7379 ( .A(n6817), .B(n6816), .Z(n7130) );
  NANDN U7380 ( .A(n3010), .B(\stack[1][20] ), .Z(n7126) );
  NANDN U7381 ( .A(n6819), .B(n6818), .Z(n6823) );
  NANDN U7382 ( .A(n6821), .B(n6820), .Z(n6822) );
  NAND U7383 ( .A(n6823), .B(n6822), .Z(n7124) );
  NANDN U7384 ( .A(n3008), .B(\stack[1][22] ), .Z(n7043) );
  NANDN U7385 ( .A(n6825), .B(n6824), .Z(n6829) );
  NANDN U7386 ( .A(n6827), .B(n6826), .Z(n6828) );
  NAND U7387 ( .A(n6829), .B(n6828), .Z(n7041) );
  AND U7388 ( .A(\stack[1][23] ), .B(o[13]), .Z(n7117) );
  OR U7389 ( .A(n6831), .B(n6830), .Z(n6835) );
  OR U7390 ( .A(n6833), .B(n6832), .Z(n6834) );
  NAND U7391 ( .A(n6835), .B(n6834), .Z(n7118) );
  XNOR U7392 ( .A(n7117), .B(n7118), .Z(n7120) );
  OR U7393 ( .A(n6837), .B(n6836), .Z(n6841) );
  OR U7394 ( .A(n6839), .B(n6838), .Z(n6840) );
  NAND U7395 ( .A(n6841), .B(n6840), .Z(n7053) );
  ANDN U7396 ( .B(o[11]), .A(n2982), .Z(n7052) );
  XOR U7397 ( .A(n7053), .B(n7052), .Z(n7054) );
  NANDN U7398 ( .A(n3004), .B(\stack[1][26] ), .Z(n7114) );
  OR U7399 ( .A(n6843), .B(n6842), .Z(n6847) );
  OR U7400 ( .A(n6845), .B(n6844), .Z(n6846) );
  NAND U7401 ( .A(n6847), .B(n6846), .Z(n7112) );
  NANDN U7402 ( .A(n3002), .B(\stack[1][28] ), .Z(n7108) );
  OR U7403 ( .A(n6849), .B(n6848), .Z(n6853) );
  OR U7404 ( .A(n6851), .B(n6850), .Z(n6852) );
  NAND U7405 ( .A(n6853), .B(n6852), .Z(n7106) );
  OR U7406 ( .A(n6855), .B(n6854), .Z(n6859) );
  OR U7407 ( .A(n6857), .B(n6856), .Z(n6858) );
  AND U7408 ( .A(n6859), .B(n6858), .Z(n7064) );
  AND U7409 ( .A(\stack[1][29] ), .B(o[7]), .Z(n7065) );
  XNOR U7410 ( .A(n7064), .B(n7065), .Z(n7067) );
  OR U7411 ( .A(n6861), .B(n6860), .Z(n6865) );
  OR U7412 ( .A(n6863), .B(n6862), .Z(n6864) );
  AND U7413 ( .A(n6865), .B(n6864), .Z(n7070) );
  OR U7414 ( .A(n6867), .B(n6866), .Z(n6871) );
  OR U7415 ( .A(n6869), .B(n6868), .Z(n6870) );
  NAND U7416 ( .A(n6871), .B(n6870), .Z(n7100) );
  NANDN U7417 ( .A(n6873), .B(n6872), .Z(n6879) );
  ANDN U7418 ( .B(\stack[1][33] ), .A(n2994), .Z(n6875) );
  NAND U7419 ( .A(n6875), .B(n6874), .Z(n6877) );
  NANDN U7420 ( .A(n2990), .B(o[2]), .Z(n6876) );
  AND U7421 ( .A(n6877), .B(n6876), .Z(n6878) );
  ANDN U7422 ( .B(n6879), .A(n6878), .Z(n7082) );
  AND U7423 ( .A(\stack[1][33] ), .B(o[3]), .Z(n7083) );
  XNOR U7424 ( .A(n7082), .B(n7083), .Z(n7085) );
  ANDN U7425 ( .B(o[0]), .A(n2993), .Z(n6881) );
  NANDN U7426 ( .A(n2995), .B(\stack[1][35] ), .Z(n6880) );
  XNOR U7427 ( .A(n6881), .B(n6880), .Z(n7089) );
  AND U7428 ( .A(\stack[1][35] ), .B(o[1]), .Z(n7090) );
  NANDN U7429 ( .A(n2994), .B(n7090), .Z(n6882) );
  XOR U7430 ( .A(n2996), .B(n6882), .Z(n6883) );
  AND U7431 ( .A(n6883), .B(\stack[1][34] ), .Z(n7088) );
  XOR U7432 ( .A(n7089), .B(n7088), .Z(n7084) );
  XOR U7433 ( .A(n7085), .B(n7084), .Z(n7099) );
  XNOR U7434 ( .A(n7100), .B(n7099), .Z(n7102) );
  AND U7435 ( .A(\stack[1][32] ), .B(o[4]), .Z(n7101) );
  XNOR U7436 ( .A(n7102), .B(n7101), .Z(n7078) );
  AND U7437 ( .A(\stack[1][31] ), .B(o[5]), .Z(n7076) );
  OR U7438 ( .A(n6885), .B(n6884), .Z(n6889) );
  NANDN U7439 ( .A(n6887), .B(n6886), .Z(n6888) );
  NAND U7440 ( .A(n6889), .B(n6888), .Z(n7077) );
  XNOR U7441 ( .A(n7076), .B(n7077), .Z(n7079) );
  XNOR U7442 ( .A(n7078), .B(n7079), .Z(n7071) );
  XOR U7443 ( .A(n7070), .B(n7071), .Z(n7072) );
  AND U7444 ( .A(\stack[1][30] ), .B(o[6]), .Z(n7073) );
  XOR U7445 ( .A(n7072), .B(n7073), .Z(n7066) );
  XOR U7446 ( .A(n7067), .B(n7066), .Z(n7105) );
  XNOR U7447 ( .A(n7106), .B(n7105), .Z(n7107) );
  XNOR U7448 ( .A(n7108), .B(n7107), .Z(n7060) );
  AND U7449 ( .A(\stack[1][27] ), .B(o[9]), .Z(n7058) );
  NANDN U7450 ( .A(n6891), .B(n6890), .Z(n6895) );
  NANDN U7451 ( .A(n6893), .B(n6892), .Z(n6894) );
  NAND U7452 ( .A(n6895), .B(n6894), .Z(n7059) );
  XNOR U7453 ( .A(n7058), .B(n7059), .Z(n7061) );
  XNOR U7454 ( .A(n7060), .B(n7061), .Z(n7111) );
  XNOR U7455 ( .A(n7112), .B(n7111), .Z(n7113) );
  XNOR U7456 ( .A(n7114), .B(n7113), .Z(n7055) );
  OR U7457 ( .A(n6897), .B(n6896), .Z(n6901) );
  OR U7458 ( .A(n6899), .B(n6898), .Z(n6900) );
  AND U7459 ( .A(n6901), .B(n6900), .Z(n7047) );
  XNOR U7460 ( .A(n7046), .B(n7047), .Z(n7049) );
  AND U7461 ( .A(\stack[1][24] ), .B(o[12]), .Z(n7048) );
  XNOR U7462 ( .A(n7049), .B(n7048), .Z(n7119) );
  XOR U7463 ( .A(n7120), .B(n7119), .Z(n7040) );
  XNOR U7464 ( .A(n7041), .B(n7040), .Z(n7042) );
  XNOR U7465 ( .A(n7043), .B(n7042), .Z(n7036) );
  NANDN U7466 ( .A(n2978), .B(o[15]), .Z(n7034) );
  OR U7467 ( .A(n6903), .B(n6902), .Z(n6907) );
  OR U7468 ( .A(n6905), .B(n6904), .Z(n6906) );
  NAND U7469 ( .A(n6907), .B(n6906), .Z(n7035) );
  XOR U7470 ( .A(n7034), .B(n7035), .Z(n7037) );
  XNOR U7471 ( .A(n7036), .B(n7037), .Z(n7123) );
  XNOR U7472 ( .A(n7124), .B(n7123), .Z(n7125) );
  XNOR U7473 ( .A(n7126), .B(n7125), .Z(n7030) );
  NANDN U7474 ( .A(n16746), .B(o[17]), .Z(n7028) );
  OR U7475 ( .A(n6909), .B(n6908), .Z(n6913) );
  OR U7476 ( .A(n6911), .B(n6910), .Z(n6912) );
  NAND U7477 ( .A(n6913), .B(n6912), .Z(n7029) );
  XOR U7478 ( .A(n7028), .B(n7029), .Z(n7031) );
  XNOR U7479 ( .A(n7030), .B(n7031), .Z(n7129) );
  XNOR U7480 ( .A(n7130), .B(n7129), .Z(n7132) );
  XOR U7481 ( .A(n7131), .B(n7132), .Z(n7024) );
  NANDN U7482 ( .A(n3013), .B(\stack[1][17] ), .Z(n7022) );
  OR U7483 ( .A(n6915), .B(n6914), .Z(n6919) );
  OR U7484 ( .A(n6917), .B(n6916), .Z(n6918) );
  NAND U7485 ( .A(n6919), .B(n6918), .Z(n7023) );
  XOR U7486 ( .A(n7022), .B(n7023), .Z(n7025) );
  XNOR U7487 ( .A(n7024), .B(n7025), .Z(n7135) );
  XNOR U7488 ( .A(n7136), .B(n7135), .Z(n7137) );
  XNOR U7489 ( .A(n7138), .B(n7137), .Z(n7018) );
  NANDN U7490 ( .A(n3015), .B(\stack[1][15] ), .Z(n7016) );
  OR U7491 ( .A(n6921), .B(n6920), .Z(n6925) );
  OR U7492 ( .A(n6923), .B(n6922), .Z(n6924) );
  NAND U7493 ( .A(n6925), .B(n6924), .Z(n7017) );
  XOR U7494 ( .A(n7016), .B(n7017), .Z(n7019) );
  XNOR U7495 ( .A(n7018), .B(n7019), .Z(n7141) );
  XNOR U7496 ( .A(n7142), .B(n7141), .Z(n7143) );
  XNOR U7497 ( .A(n7144), .B(n7143), .Z(n7012) );
  NANDN U7498 ( .A(n3017), .B(\stack[1][13] ), .Z(n7010) );
  OR U7499 ( .A(n6927), .B(n6926), .Z(n6931) );
  OR U7500 ( .A(n6929), .B(n6928), .Z(n6930) );
  NAND U7501 ( .A(n6931), .B(n6930), .Z(n7011) );
  XOR U7502 ( .A(n7010), .B(n7011), .Z(n7013) );
  XNOR U7503 ( .A(n7012), .B(n7013), .Z(n7147) );
  XNOR U7504 ( .A(n7148), .B(n7147), .Z(n7149) );
  XNOR U7505 ( .A(n7150), .B(n7149), .Z(n7006) );
  NANDN U7506 ( .A(n3019), .B(\stack[1][11] ), .Z(n7004) );
  OR U7507 ( .A(n6933), .B(n6932), .Z(n6937) );
  OR U7508 ( .A(n6935), .B(n6934), .Z(n6936) );
  NAND U7509 ( .A(n6937), .B(n6936), .Z(n7005) );
  XOR U7510 ( .A(n7004), .B(n7005), .Z(n7007) );
  XNOR U7511 ( .A(n7006), .B(n7007), .Z(n7153) );
  XNOR U7512 ( .A(n7154), .B(n7153), .Z(n7155) );
  XNOR U7513 ( .A(n7156), .B(n7155), .Z(n7000) );
  NANDN U7514 ( .A(n17145), .B(o[27]), .Z(n6998) );
  OR U7515 ( .A(n6939), .B(n6938), .Z(n6943) );
  OR U7516 ( .A(n6941), .B(n6940), .Z(n6942) );
  NAND U7517 ( .A(n6943), .B(n6942), .Z(n6999) );
  XOR U7518 ( .A(n6998), .B(n6999), .Z(n7001) );
  XNOR U7519 ( .A(n7000), .B(n7001), .Z(n7159) );
  XNOR U7520 ( .A(n7160), .B(n7159), .Z(n7161) );
  XNOR U7521 ( .A(n7162), .B(n7161), .Z(n6994) );
  NANDN U7522 ( .A(n17219), .B(o[29]), .Z(n6992) );
  OR U7523 ( .A(n6945), .B(n6944), .Z(n6949) );
  OR U7524 ( .A(n6947), .B(n6946), .Z(n6948) );
  NAND U7525 ( .A(n6949), .B(n6948), .Z(n6993) );
  XOR U7526 ( .A(n6992), .B(n6993), .Z(n6995) );
  XNOR U7527 ( .A(n6994), .B(n6995), .Z(n7165) );
  XNOR U7528 ( .A(n7166), .B(n7165), .Z(n7167) );
  XNOR U7529 ( .A(n7168), .B(n7167), .Z(n6988) );
  NANDN U7530 ( .A(n17296), .B(o[31]), .Z(n6986) );
  OR U7531 ( .A(n6951), .B(n6950), .Z(n6955) );
  OR U7532 ( .A(n6953), .B(n6952), .Z(n6954) );
  NAND U7533 ( .A(n6955), .B(n6954), .Z(n6987) );
  XOR U7534 ( .A(n6986), .B(n6987), .Z(n6989) );
  XNOR U7535 ( .A(n6988), .B(n6989), .Z(n7171) );
  XNOR U7536 ( .A(n7172), .B(n7171), .Z(n7173) );
  XNOR U7537 ( .A(n7174), .B(n7173), .Z(n6982) );
  NANDN U7538 ( .A(n17375), .B(o[33]), .Z(n6980) );
  OR U7539 ( .A(n6957), .B(n6956), .Z(n6961) );
  OR U7540 ( .A(n6959), .B(n6958), .Z(n6960) );
  NAND U7541 ( .A(n6961), .B(n6960), .Z(n6981) );
  XOR U7542 ( .A(n6980), .B(n6981), .Z(n6983) );
  XNOR U7543 ( .A(n6982), .B(n6983), .Z(n7177) );
  XNOR U7544 ( .A(n7178), .B(n7177), .Z(n7179) );
  AND U7545 ( .A(o[35]), .B(\stack[1][1] ), .Z(n6974) );
  OR U7546 ( .A(n6963), .B(n6962), .Z(n6967) );
  OR U7547 ( .A(n6965), .B(n6964), .Z(n6966) );
  NAND U7548 ( .A(n6967), .B(n6966), .Z(n6975) );
  XNOR U7549 ( .A(n6974), .B(n6975), .Z(n6977) );
  XOR U7550 ( .A(n6976), .B(n6977), .Z(n6968) );
  NANDN U7551 ( .A(n6969), .B(n6968), .Z(n6971) );
  XOR U7552 ( .A(n6969), .B(n6968), .Z(n16090) );
  AND U7553 ( .A(o[36]), .B(\stack[1][0] ), .Z(n16091) );
  OR U7554 ( .A(n16090), .B(n16091), .Z(n6970) );
  AND U7555 ( .A(n6971), .B(n6970), .Z(n6973) );
  OR U7556 ( .A(n6972), .B(n6973), .Z(n7184) );
  XNOR U7557 ( .A(n6973), .B(n6972), .Z(n16052) );
  NANDN U7558 ( .A(n2969), .B(o[36]), .Z(n7397) );
  OR U7559 ( .A(n6975), .B(n6974), .Z(n6979) );
  OR U7560 ( .A(n6977), .B(n6976), .Z(n6978) );
  NAND U7561 ( .A(n6979), .B(n6978), .Z(n7395) );
  NANDN U7562 ( .A(n17375), .B(o[34]), .Z(n7391) );
  NANDN U7563 ( .A(n6981), .B(n6980), .Z(n6985) );
  NANDN U7564 ( .A(n6983), .B(n6982), .Z(n6984) );
  NAND U7565 ( .A(n6985), .B(n6984), .Z(n7389) );
  NANDN U7566 ( .A(n17296), .B(o[32]), .Z(n7385) );
  NANDN U7567 ( .A(n6987), .B(n6986), .Z(n6991) );
  NANDN U7568 ( .A(n6989), .B(n6988), .Z(n6990) );
  NAND U7569 ( .A(n6991), .B(n6990), .Z(n7383) );
  NANDN U7570 ( .A(n17219), .B(o[30]), .Z(n7379) );
  NANDN U7571 ( .A(n6993), .B(n6992), .Z(n6997) );
  NANDN U7572 ( .A(n6995), .B(n6994), .Z(n6996) );
  NAND U7573 ( .A(n6997), .B(n6996), .Z(n7377) );
  NANDN U7574 ( .A(n17145), .B(o[28]), .Z(n7373) );
  NANDN U7575 ( .A(n6999), .B(n6998), .Z(n7003) );
  NANDN U7576 ( .A(n7001), .B(n7000), .Z(n7002) );
  NAND U7577 ( .A(n7003), .B(n7002), .Z(n7371) );
  NANDN U7578 ( .A(n2972), .B(o[26]), .Z(n7367) );
  NANDN U7579 ( .A(n7005), .B(n7004), .Z(n7009) );
  NANDN U7580 ( .A(n7007), .B(n7006), .Z(n7008) );
  NAND U7581 ( .A(n7009), .B(n7008), .Z(n7365) );
  NANDN U7582 ( .A(n2974), .B(o[24]), .Z(n7361) );
  NANDN U7583 ( .A(n7011), .B(n7010), .Z(n7015) );
  NANDN U7584 ( .A(n7013), .B(n7012), .Z(n7014) );
  NAND U7585 ( .A(n7015), .B(n7014), .Z(n7359) );
  NANDN U7586 ( .A(n2976), .B(o[22]), .Z(n7230) );
  NANDN U7587 ( .A(n7017), .B(n7016), .Z(n7021) );
  NANDN U7588 ( .A(n7019), .B(n7018), .Z(n7020) );
  NAND U7589 ( .A(n7021), .B(n7020), .Z(n7228) );
  NANDN U7590 ( .A(n16826), .B(o[20]), .Z(n7355) );
  NANDN U7591 ( .A(n7023), .B(n7022), .Z(n7027) );
  NANDN U7592 ( .A(n7025), .B(n7024), .Z(n7026) );
  NAND U7593 ( .A(n7027), .B(n7026), .Z(n7353) );
  NANDN U7594 ( .A(n3012), .B(\stack[1][19] ), .Z(n7349) );
  NANDN U7595 ( .A(n7029), .B(n7028), .Z(n7033) );
  NANDN U7596 ( .A(n7031), .B(n7030), .Z(n7032) );
  NAND U7597 ( .A(n7033), .B(n7032), .Z(n7347) );
  AND U7598 ( .A(\stack[1][21] ), .B(o[16]), .Z(n7254) );
  NANDN U7599 ( .A(n7035), .B(n7034), .Z(n7039) );
  NANDN U7600 ( .A(n7037), .B(n7036), .Z(n7038) );
  AND U7601 ( .A(n7039), .B(n7038), .Z(n7251) );
  AND U7602 ( .A(\stack[1][22] ), .B(o[15]), .Z(n7340) );
  OR U7603 ( .A(n7041), .B(n7040), .Z(n7045) );
  OR U7604 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U7605 ( .A(n7045), .B(n7044), .Z(n7341) );
  XNOR U7606 ( .A(n7340), .B(n7341), .Z(n7343) );
  OR U7607 ( .A(n7047), .B(n7046), .Z(n7051) );
  OR U7608 ( .A(n7049), .B(n7048), .Z(n7050) );
  NAND U7609 ( .A(n7051), .B(n7050), .Z(n7264) );
  ANDN U7610 ( .B(o[13]), .A(n2981), .Z(n7263) );
  XNOR U7611 ( .A(n7264), .B(n7263), .Z(n7265) );
  NANDN U7612 ( .A(n3006), .B(\stack[1][25] ), .Z(n7337) );
  NANDN U7613 ( .A(n7053), .B(n7052), .Z(n7057) );
  OR U7614 ( .A(n7055), .B(n7054), .Z(n7056) );
  AND U7615 ( .A(n7057), .B(n7056), .Z(n7334) );
  NANDN U7616 ( .A(n3004), .B(\stack[1][27] ), .Z(n7331) );
  OR U7617 ( .A(n7059), .B(n7058), .Z(n7063) );
  NANDN U7618 ( .A(n7061), .B(n7060), .Z(n7062) );
  NAND U7619 ( .A(n7063), .B(n7062), .Z(n7329) );
  NANDN U7620 ( .A(n3002), .B(\stack[1][29] ), .Z(n7325) );
  OR U7621 ( .A(n7065), .B(n7064), .Z(n7069) );
  OR U7622 ( .A(n7067), .B(n7066), .Z(n7068) );
  NAND U7623 ( .A(n7069), .B(n7068), .Z(n7323) );
  OR U7624 ( .A(n7071), .B(n7070), .Z(n7075) );
  NANDN U7625 ( .A(n7073), .B(n7072), .Z(n7074) );
  AND U7626 ( .A(n7075), .B(n7074), .Z(n7281) );
  AND U7627 ( .A(\stack[1][30] ), .B(o[7]), .Z(n7282) );
  XNOR U7628 ( .A(n7281), .B(n7282), .Z(n7284) );
  OR U7629 ( .A(n7077), .B(n7076), .Z(n7081) );
  OR U7630 ( .A(n7079), .B(n7078), .Z(n7080) );
  AND U7631 ( .A(n7081), .B(n7080), .Z(n7287) );
  OR U7632 ( .A(n7083), .B(n7082), .Z(n7087) );
  OR U7633 ( .A(n7085), .B(n7084), .Z(n7086) );
  NAND U7634 ( .A(n7087), .B(n7086), .Z(n7317) );
  NANDN U7635 ( .A(n7089), .B(n7088), .Z(n7095) );
  ANDN U7636 ( .B(\stack[1][34] ), .A(n2994), .Z(n7091) );
  NAND U7637 ( .A(n7091), .B(n7090), .Z(n7093) );
  NANDN U7638 ( .A(n2991), .B(o[2]), .Z(n7092) );
  AND U7639 ( .A(n7093), .B(n7092), .Z(n7094) );
  ANDN U7640 ( .B(n7095), .A(n7094), .Z(n7299) );
  AND U7641 ( .A(\stack[1][34] ), .B(o[3]), .Z(n7300) );
  XNOR U7642 ( .A(n7299), .B(n7300), .Z(n7302) );
  ANDN U7643 ( .B(\stack[1][37] ), .A(n2994), .Z(n7540) );
  NANDN U7644 ( .A(n2995), .B(\stack[1][36] ), .Z(n7096) );
  XNOR U7645 ( .A(n7540), .B(n7096), .Z(n7306) );
  AND U7646 ( .A(\stack[1][36] ), .B(o[1]), .Z(n7307) );
  NANDN U7647 ( .A(n2994), .B(n7307), .Z(n7097) );
  XOR U7648 ( .A(n2996), .B(n7097), .Z(n7098) );
  AND U7649 ( .A(n7098), .B(\stack[1][35] ), .Z(n7305) );
  XOR U7650 ( .A(n7306), .B(n7305), .Z(n7301) );
  XOR U7651 ( .A(n7302), .B(n7301), .Z(n7316) );
  XNOR U7652 ( .A(n7317), .B(n7316), .Z(n7319) );
  AND U7653 ( .A(\stack[1][33] ), .B(o[4]), .Z(n7318) );
  XNOR U7654 ( .A(n7319), .B(n7318), .Z(n7295) );
  AND U7655 ( .A(\stack[1][32] ), .B(o[5]), .Z(n7293) );
  OR U7656 ( .A(n7100), .B(n7099), .Z(n7104) );
  NANDN U7657 ( .A(n7102), .B(n7101), .Z(n7103) );
  NAND U7658 ( .A(n7104), .B(n7103), .Z(n7294) );
  XNOR U7659 ( .A(n7293), .B(n7294), .Z(n7296) );
  XNOR U7660 ( .A(n7295), .B(n7296), .Z(n7288) );
  XOR U7661 ( .A(n7287), .B(n7288), .Z(n7289) );
  AND U7662 ( .A(\stack[1][31] ), .B(o[6]), .Z(n7290) );
  XOR U7663 ( .A(n7289), .B(n7290), .Z(n7283) );
  XOR U7664 ( .A(n7284), .B(n7283), .Z(n7322) );
  XNOR U7665 ( .A(n7323), .B(n7322), .Z(n7324) );
  XNOR U7666 ( .A(n7325), .B(n7324), .Z(n7277) );
  NANDN U7667 ( .A(n2985), .B(o[9]), .Z(n7275) );
  OR U7668 ( .A(n7106), .B(n7105), .Z(n7110) );
  OR U7669 ( .A(n7108), .B(n7107), .Z(n7109) );
  NAND U7670 ( .A(n7110), .B(n7109), .Z(n7276) );
  XOR U7671 ( .A(n7275), .B(n7276), .Z(n7278) );
  XNOR U7672 ( .A(n7277), .B(n7278), .Z(n7328) );
  XNOR U7673 ( .A(n7329), .B(n7328), .Z(n7330) );
  XNOR U7674 ( .A(n7331), .B(n7330), .Z(n7271) );
  NANDN U7675 ( .A(n2983), .B(o[11]), .Z(n7269) );
  OR U7676 ( .A(n7112), .B(n7111), .Z(n7116) );
  OR U7677 ( .A(n7114), .B(n7113), .Z(n7115) );
  NAND U7678 ( .A(n7116), .B(n7115), .Z(n7270) );
  XOR U7679 ( .A(n7269), .B(n7270), .Z(n7272) );
  XNOR U7680 ( .A(n7271), .B(n7272), .Z(n7335) );
  XNOR U7681 ( .A(n7334), .B(n7335), .Z(n7336) );
  XOR U7682 ( .A(n7265), .B(n7266), .Z(n7257) );
  OR U7683 ( .A(n7118), .B(n7117), .Z(n7122) );
  OR U7684 ( .A(n7120), .B(n7119), .Z(n7121) );
  AND U7685 ( .A(n7122), .B(n7121), .Z(n7258) );
  XOR U7686 ( .A(n7257), .B(n7258), .Z(n7260) );
  AND U7687 ( .A(\stack[1][23] ), .B(o[14]), .Z(n7259) );
  XOR U7688 ( .A(n7260), .B(n7259), .Z(n7342) );
  XOR U7689 ( .A(n7343), .B(n7342), .Z(n7252) );
  XOR U7690 ( .A(n7251), .B(n7252), .Z(n7253) );
  XOR U7691 ( .A(n7254), .B(n7253), .Z(n7248) );
  AND U7692 ( .A(\stack[1][20] ), .B(o[17]), .Z(n7245) );
  OR U7693 ( .A(n7124), .B(n7123), .Z(n7128) );
  OR U7694 ( .A(n7126), .B(n7125), .Z(n7127) );
  NAND U7695 ( .A(n7128), .B(n7127), .Z(n7246) );
  XNOR U7696 ( .A(n7245), .B(n7246), .Z(n7247) );
  XOR U7697 ( .A(n7248), .B(n7247), .Z(n7346) );
  XNOR U7698 ( .A(n7347), .B(n7346), .Z(n7348) );
  XNOR U7699 ( .A(n7349), .B(n7348), .Z(n7241) );
  NANDN U7700 ( .A(n3013), .B(\stack[1][18] ), .Z(n7239) );
  OR U7701 ( .A(n7130), .B(n7129), .Z(n7134) );
  IV U7702 ( .A(n7131), .Z(n16787) );
  OR U7703 ( .A(n7132), .B(n16787), .Z(n7133) );
  NAND U7704 ( .A(n7134), .B(n7133), .Z(n7240) );
  XOR U7705 ( .A(n7239), .B(n7240), .Z(n7242) );
  XNOR U7706 ( .A(n7241), .B(n7242), .Z(n7352) );
  XNOR U7707 ( .A(n7353), .B(n7352), .Z(n7354) );
  XNOR U7708 ( .A(n7355), .B(n7354), .Z(n7235) );
  NANDN U7709 ( .A(n3015), .B(\stack[1][16] ), .Z(n7233) );
  OR U7710 ( .A(n7136), .B(n7135), .Z(n7140) );
  OR U7711 ( .A(n7138), .B(n7137), .Z(n7139) );
  NAND U7712 ( .A(n7140), .B(n7139), .Z(n7234) );
  XOR U7713 ( .A(n7233), .B(n7234), .Z(n7236) );
  XNOR U7714 ( .A(n7235), .B(n7236), .Z(n7227) );
  XNOR U7715 ( .A(n7228), .B(n7227), .Z(n7229) );
  XNOR U7716 ( .A(n7230), .B(n7229), .Z(n7223) );
  NANDN U7717 ( .A(n3017), .B(\stack[1][14] ), .Z(n7221) );
  OR U7718 ( .A(n7142), .B(n7141), .Z(n7146) );
  OR U7719 ( .A(n7144), .B(n7143), .Z(n7145) );
  NAND U7720 ( .A(n7146), .B(n7145), .Z(n7222) );
  XOR U7721 ( .A(n7221), .B(n7222), .Z(n7224) );
  XNOR U7722 ( .A(n7223), .B(n7224), .Z(n7358) );
  XNOR U7723 ( .A(n7359), .B(n7358), .Z(n7360) );
  XNOR U7724 ( .A(n7361), .B(n7360), .Z(n7217) );
  NANDN U7725 ( .A(n3019), .B(\stack[1][12] ), .Z(n7215) );
  OR U7726 ( .A(n7148), .B(n7147), .Z(n7152) );
  OR U7727 ( .A(n7150), .B(n7149), .Z(n7151) );
  NAND U7728 ( .A(n7152), .B(n7151), .Z(n7216) );
  XOR U7729 ( .A(n7215), .B(n7216), .Z(n7218) );
  XNOR U7730 ( .A(n7217), .B(n7218), .Z(n7364) );
  XNOR U7731 ( .A(n7365), .B(n7364), .Z(n7366) );
  XNOR U7732 ( .A(n7367), .B(n7366), .Z(n7211) );
  NANDN U7733 ( .A(n17101), .B(o[27]), .Z(n7209) );
  OR U7734 ( .A(n7154), .B(n7153), .Z(n7158) );
  OR U7735 ( .A(n7156), .B(n7155), .Z(n7157) );
  NAND U7736 ( .A(n7158), .B(n7157), .Z(n7210) );
  XOR U7737 ( .A(n7209), .B(n7210), .Z(n7212) );
  XNOR U7738 ( .A(n7211), .B(n7212), .Z(n7370) );
  XNOR U7739 ( .A(n7371), .B(n7370), .Z(n7372) );
  XNOR U7740 ( .A(n7373), .B(n7372), .Z(n7205) );
  NANDN U7741 ( .A(n17179), .B(o[29]), .Z(n7203) );
  OR U7742 ( .A(n7160), .B(n7159), .Z(n7164) );
  OR U7743 ( .A(n7162), .B(n7161), .Z(n7163) );
  NAND U7744 ( .A(n7164), .B(n7163), .Z(n7204) );
  XOR U7745 ( .A(n7203), .B(n7204), .Z(n7206) );
  XNOR U7746 ( .A(n7205), .B(n7206), .Z(n7376) );
  XNOR U7747 ( .A(n7377), .B(n7376), .Z(n7378) );
  XNOR U7748 ( .A(n7379), .B(n7378), .Z(n7199) );
  NANDN U7749 ( .A(n17256), .B(o[31]), .Z(n7197) );
  OR U7750 ( .A(n7166), .B(n7165), .Z(n7170) );
  OR U7751 ( .A(n7168), .B(n7167), .Z(n7169) );
  NAND U7752 ( .A(n7170), .B(n7169), .Z(n7198) );
  XOR U7753 ( .A(n7197), .B(n7198), .Z(n7200) );
  XNOR U7754 ( .A(n7199), .B(n7200), .Z(n7382) );
  XNOR U7755 ( .A(n7383), .B(n7382), .Z(n7384) );
  XNOR U7756 ( .A(n7385), .B(n7384), .Z(n7193) );
  AND U7757 ( .A(o[33]), .B(\stack[1][4] ), .Z(n7191) );
  OR U7758 ( .A(n7172), .B(n7171), .Z(n7176) );
  OR U7759 ( .A(n7174), .B(n7173), .Z(n7175) );
  NAND U7760 ( .A(n7176), .B(n7175), .Z(n7192) );
  XNOR U7761 ( .A(n7191), .B(n7192), .Z(n7194) );
  XNOR U7762 ( .A(n7193), .B(n7194), .Z(n7388) );
  XNOR U7763 ( .A(n7389), .B(n7388), .Z(n7390) );
  XOR U7764 ( .A(n7391), .B(n7390), .Z(n7188) );
  AND U7765 ( .A(o[35]), .B(\stack[1][2] ), .Z(n7185) );
  OR U7766 ( .A(n7178), .B(n7177), .Z(n7182) );
  OR U7767 ( .A(n7180), .B(n7179), .Z(n7181) );
  NAND U7768 ( .A(n7182), .B(n7181), .Z(n7186) );
  XOR U7769 ( .A(n7185), .B(n7186), .Z(n7187) );
  XNOR U7770 ( .A(n7188), .B(n7187), .Z(n7394) );
  XNOR U7771 ( .A(n7395), .B(n7394), .Z(n7396) );
  XOR U7772 ( .A(n7397), .B(n7396), .Z(n16053) );
  OR U7773 ( .A(n16052), .B(n16053), .Z(n7183) );
  AND U7774 ( .A(n7184), .B(n7183), .Z(n7401) );
  NANDN U7775 ( .A(n2970), .B(o[36]), .Z(n7626) );
  OR U7776 ( .A(n7186), .B(n7185), .Z(n7190) );
  NANDN U7777 ( .A(n7188), .B(n7187), .Z(n7189) );
  NAND U7778 ( .A(n7190), .B(n7189), .Z(n7624) );
  NANDN U7779 ( .A(n2971), .B(o[34]), .Z(n7620) );
  OR U7780 ( .A(n7192), .B(n7191), .Z(n7196) );
  NANDN U7781 ( .A(n7194), .B(n7193), .Z(n7195) );
  NAND U7782 ( .A(n7196), .B(n7195), .Z(n7618) );
  NANDN U7783 ( .A(n17256), .B(o[32]), .Z(n7614) );
  NANDN U7784 ( .A(n7198), .B(n7197), .Z(n7202) );
  NANDN U7785 ( .A(n7200), .B(n7199), .Z(n7201) );
  NAND U7786 ( .A(n7202), .B(n7201), .Z(n7612) );
  NANDN U7787 ( .A(n17179), .B(o[30]), .Z(n7608) );
  NANDN U7788 ( .A(n7204), .B(n7203), .Z(n7208) );
  NANDN U7789 ( .A(n7206), .B(n7205), .Z(n7207) );
  NAND U7790 ( .A(n7208), .B(n7207), .Z(n7606) );
  NANDN U7791 ( .A(n17101), .B(o[28]), .Z(n7602) );
  NANDN U7792 ( .A(n7210), .B(n7209), .Z(n7214) );
  NANDN U7793 ( .A(n7212), .B(n7211), .Z(n7213) );
  NAND U7794 ( .A(n7214), .B(n7213), .Z(n7600) );
  NANDN U7795 ( .A(n2973), .B(o[26]), .Z(n7596) );
  NANDN U7796 ( .A(n7216), .B(n7215), .Z(n7220) );
  NANDN U7797 ( .A(n7218), .B(n7217), .Z(n7219) );
  NAND U7798 ( .A(n7220), .B(n7219), .Z(n7594) );
  AND U7799 ( .A(o[24]), .B(\stack[1][14] ), .Z(n7451) );
  NANDN U7800 ( .A(n7222), .B(n7221), .Z(n7226) );
  NANDN U7801 ( .A(n7224), .B(n7223), .Z(n7225) );
  AND U7802 ( .A(n7226), .B(n7225), .Z(n7448) );
  AND U7803 ( .A(o[23]), .B(\stack[1][15] ), .Z(n7587) );
  OR U7804 ( .A(n7228), .B(n7227), .Z(n7232) );
  OR U7805 ( .A(n7230), .B(n7229), .Z(n7231) );
  NAND U7806 ( .A(n7232), .B(n7231), .Z(n7588) );
  XNOR U7807 ( .A(n7587), .B(n7588), .Z(n7590) );
  NANDN U7808 ( .A(n7234), .B(n7233), .Z(n7238) );
  NANDN U7809 ( .A(n7236), .B(n7235), .Z(n7237) );
  AND U7810 ( .A(n7238), .B(n7237), .Z(n7454) );
  NANDN U7811 ( .A(n7240), .B(n7239), .Z(n7244) );
  NANDN U7812 ( .A(n7242), .B(n7241), .Z(n7243) );
  NAND U7813 ( .A(n7244), .B(n7243), .Z(n7582) );
  AND U7814 ( .A(\stack[1][20] ), .B(o[18]), .Z(n7474) );
  OR U7815 ( .A(n7246), .B(n7245), .Z(n7250) );
  OR U7816 ( .A(n7248), .B(n7247), .Z(n7249) );
  AND U7817 ( .A(n7250), .B(n7249), .Z(n7471) );
  OR U7818 ( .A(n7252), .B(n7251), .Z(n7256) );
  NANDN U7819 ( .A(n7254), .B(n7253), .Z(n7255) );
  AND U7820 ( .A(n7256), .B(n7255), .Z(n7575) );
  AND U7821 ( .A(\stack[1][21] ), .B(o[17]), .Z(n7576) );
  XNOR U7822 ( .A(n7575), .B(n7576), .Z(n7578) );
  NANDN U7823 ( .A(n7258), .B(n7257), .Z(n7262) );
  OR U7824 ( .A(n7260), .B(n7259), .Z(n7261) );
  NAND U7825 ( .A(n7262), .B(n7261), .Z(n7484) );
  ANDN U7826 ( .B(o[15]), .A(n2980), .Z(n7483) );
  XNOR U7827 ( .A(n7484), .B(n7483), .Z(n7485) );
  NANDN U7828 ( .A(n3008), .B(\stack[1][24] ), .Z(n7572) );
  NANDN U7829 ( .A(n7264), .B(n7263), .Z(n7268) );
  NANDN U7830 ( .A(n7266), .B(n7265), .Z(n7267) );
  AND U7831 ( .A(n7268), .B(n7267), .Z(n7569) );
  NANDN U7832 ( .A(n3006), .B(\stack[1][26] ), .Z(n7566) );
  NANDN U7833 ( .A(n7270), .B(n7269), .Z(n7274) );
  NANDN U7834 ( .A(n7272), .B(n7271), .Z(n7273) );
  NAND U7835 ( .A(n7274), .B(n7273), .Z(n7564) );
  NANDN U7836 ( .A(n3004), .B(\stack[1][28] ), .Z(n7560) );
  NANDN U7837 ( .A(n7276), .B(n7275), .Z(n7280) );
  NANDN U7838 ( .A(n7278), .B(n7277), .Z(n7279) );
  NAND U7839 ( .A(n7280), .B(n7279), .Z(n7558) );
  NANDN U7840 ( .A(n3002), .B(\stack[1][30] ), .Z(n7554) );
  OR U7841 ( .A(n7282), .B(n7281), .Z(n7286) );
  OR U7842 ( .A(n7284), .B(n7283), .Z(n7285) );
  NAND U7843 ( .A(n7286), .B(n7285), .Z(n7552) );
  OR U7844 ( .A(n7288), .B(n7287), .Z(n7292) );
  NANDN U7845 ( .A(n7290), .B(n7289), .Z(n7291) );
  AND U7846 ( .A(n7292), .B(n7291), .Z(n7507) );
  AND U7847 ( .A(\stack[1][31] ), .B(o[7]), .Z(n7508) );
  XNOR U7848 ( .A(n7507), .B(n7508), .Z(n7510) );
  OR U7849 ( .A(n7294), .B(n7293), .Z(n7298) );
  OR U7850 ( .A(n7296), .B(n7295), .Z(n7297) );
  AND U7851 ( .A(n7298), .B(n7297), .Z(n7513) );
  OR U7852 ( .A(n7300), .B(n7299), .Z(n7304) );
  OR U7853 ( .A(n7302), .B(n7301), .Z(n7303) );
  NAND U7854 ( .A(n7304), .B(n7303), .Z(n7546) );
  NANDN U7855 ( .A(n7306), .B(n7305), .Z(n7312) );
  ANDN U7856 ( .B(\stack[1][35] ), .A(n2994), .Z(n7308) );
  NAND U7857 ( .A(n7308), .B(n7307), .Z(n7310) );
  NANDN U7858 ( .A(n2992), .B(o[2]), .Z(n7309) );
  AND U7859 ( .A(n7310), .B(n7309), .Z(n7311) );
  ANDN U7860 ( .B(n7312), .A(n7311), .Z(n7525) );
  AND U7861 ( .A(\stack[1][35] ), .B(o[3]), .Z(n7526) );
  XNOR U7862 ( .A(n7525), .B(n7526), .Z(n7528) );
  ANDN U7863 ( .B(\stack[1][38] ), .A(n2994), .Z(n7542) );
  NANDN U7864 ( .A(n2995), .B(\stack[1][37] ), .Z(n7313) );
  XNOR U7865 ( .A(n7542), .B(n7313), .Z(n7532) );
  AND U7866 ( .A(\stack[1][37] ), .B(o[1]), .Z(n7533) );
  NANDN U7867 ( .A(n2994), .B(n7533), .Z(n7314) );
  XOR U7868 ( .A(n2996), .B(n7314), .Z(n7315) );
  AND U7869 ( .A(n7315), .B(\stack[1][36] ), .Z(n7531) );
  XOR U7870 ( .A(n7532), .B(n7531), .Z(n7527) );
  XOR U7871 ( .A(n7528), .B(n7527), .Z(n7545) );
  XNOR U7872 ( .A(n7546), .B(n7545), .Z(n7548) );
  AND U7873 ( .A(\stack[1][34] ), .B(o[4]), .Z(n7547) );
  XNOR U7874 ( .A(n7548), .B(n7547), .Z(n7521) );
  AND U7875 ( .A(\stack[1][33] ), .B(o[5]), .Z(n7519) );
  OR U7876 ( .A(n7317), .B(n7316), .Z(n7321) );
  NANDN U7877 ( .A(n7319), .B(n7318), .Z(n7320) );
  NAND U7878 ( .A(n7321), .B(n7320), .Z(n7520) );
  XNOR U7879 ( .A(n7519), .B(n7520), .Z(n7522) );
  XNOR U7880 ( .A(n7521), .B(n7522), .Z(n7514) );
  XOR U7881 ( .A(n7513), .B(n7514), .Z(n7515) );
  AND U7882 ( .A(\stack[1][32] ), .B(o[6]), .Z(n7516) );
  XOR U7883 ( .A(n7515), .B(n7516), .Z(n7509) );
  XOR U7884 ( .A(n7510), .B(n7509), .Z(n7551) );
  XNOR U7885 ( .A(n7552), .B(n7551), .Z(n7553) );
  XNOR U7886 ( .A(n7554), .B(n7553), .Z(n7503) );
  NANDN U7887 ( .A(n2986), .B(o[9]), .Z(n7501) );
  OR U7888 ( .A(n7323), .B(n7322), .Z(n7327) );
  OR U7889 ( .A(n7325), .B(n7324), .Z(n7326) );
  NAND U7890 ( .A(n7327), .B(n7326), .Z(n7502) );
  XOR U7891 ( .A(n7501), .B(n7502), .Z(n7504) );
  XNOR U7892 ( .A(n7503), .B(n7504), .Z(n7557) );
  XNOR U7893 ( .A(n7558), .B(n7557), .Z(n7559) );
  XNOR U7894 ( .A(n7560), .B(n7559), .Z(n7497) );
  NANDN U7895 ( .A(n2984), .B(o[11]), .Z(n7495) );
  OR U7896 ( .A(n7329), .B(n7328), .Z(n7333) );
  OR U7897 ( .A(n7331), .B(n7330), .Z(n7332) );
  NAND U7898 ( .A(n7333), .B(n7332), .Z(n7496) );
  XOR U7899 ( .A(n7495), .B(n7496), .Z(n7498) );
  XNOR U7900 ( .A(n7497), .B(n7498), .Z(n7563) );
  XNOR U7901 ( .A(n7564), .B(n7563), .Z(n7565) );
  XNOR U7902 ( .A(n7566), .B(n7565), .Z(n7491) );
  NANDN U7903 ( .A(n2982), .B(o[13]), .Z(n7489) );
  OR U7904 ( .A(n7335), .B(n7334), .Z(n7339) );
  OR U7905 ( .A(n7337), .B(n7336), .Z(n7338) );
  NAND U7906 ( .A(n7339), .B(n7338), .Z(n7490) );
  XOR U7907 ( .A(n7489), .B(n7490), .Z(n7492) );
  XNOR U7908 ( .A(n7491), .B(n7492), .Z(n7570) );
  XNOR U7909 ( .A(n7569), .B(n7570), .Z(n7571) );
  XOR U7910 ( .A(n7485), .B(n7486), .Z(n7477) );
  OR U7911 ( .A(n7341), .B(n7340), .Z(n7345) );
  NANDN U7912 ( .A(n7343), .B(n7342), .Z(n7344) );
  AND U7913 ( .A(n7345), .B(n7344), .Z(n7478) );
  XOR U7914 ( .A(n7477), .B(n7478), .Z(n7480) );
  AND U7915 ( .A(\stack[1][22] ), .B(o[16]), .Z(n7479) );
  XOR U7916 ( .A(n7480), .B(n7479), .Z(n7577) );
  XOR U7917 ( .A(n7578), .B(n7577), .Z(n7472) );
  XOR U7918 ( .A(n7471), .B(n7472), .Z(n7473) );
  XOR U7919 ( .A(n7474), .B(n7473), .Z(n7468) );
  AND U7920 ( .A(o[19]), .B(\stack[1][19] ), .Z(n16747) );
  OR U7921 ( .A(n7347), .B(n7346), .Z(n7351) );
  OR U7922 ( .A(n7349), .B(n7348), .Z(n7350) );
  NAND U7923 ( .A(n7351), .B(n7350), .Z(n7466) );
  XNOR U7924 ( .A(n16747), .B(n7466), .Z(n7467) );
  XNOR U7925 ( .A(n7468), .B(n7467), .Z(n7581) );
  XOR U7926 ( .A(n7582), .B(n7581), .Z(n7584) );
  AND U7927 ( .A(o[20]), .B(\stack[1][18] ), .Z(n7583) );
  XNOR U7928 ( .A(n7584), .B(n7583), .Z(n7462) );
  AND U7929 ( .A(o[21]), .B(\stack[1][17] ), .Z(n7460) );
  OR U7930 ( .A(n7353), .B(n7352), .Z(n7357) );
  OR U7931 ( .A(n7355), .B(n7354), .Z(n7356) );
  NAND U7932 ( .A(n7357), .B(n7356), .Z(n7461) );
  XNOR U7933 ( .A(n7460), .B(n7461), .Z(n7463) );
  XNOR U7934 ( .A(n7462), .B(n7463), .Z(n7455) );
  XNOR U7935 ( .A(n7454), .B(n7455), .Z(n7456) );
  AND U7936 ( .A(o[22]), .B(\stack[1][16] ), .Z(n7457) );
  XNOR U7937 ( .A(n7590), .B(n7589), .Z(n7449) );
  XOR U7938 ( .A(n7448), .B(n7449), .Z(n7450) );
  XOR U7939 ( .A(n7451), .B(n7450), .Z(n7445) );
  AND U7940 ( .A(o[25]), .B(\stack[1][13] ), .Z(n7442) );
  OR U7941 ( .A(n7359), .B(n7358), .Z(n7363) );
  OR U7942 ( .A(n7361), .B(n7360), .Z(n7362) );
  NAND U7943 ( .A(n7363), .B(n7362), .Z(n7443) );
  XNOR U7944 ( .A(n7442), .B(n7443), .Z(n7444) );
  XOR U7945 ( .A(n7445), .B(n7444), .Z(n7593) );
  XNOR U7946 ( .A(n7594), .B(n7593), .Z(n7595) );
  XNOR U7947 ( .A(n7596), .B(n7595), .Z(n7438) );
  NANDN U7948 ( .A(n2972), .B(o[27]), .Z(n7436) );
  OR U7949 ( .A(n7365), .B(n7364), .Z(n7369) );
  OR U7950 ( .A(n7367), .B(n7366), .Z(n7368) );
  NAND U7951 ( .A(n7369), .B(n7368), .Z(n7437) );
  XOR U7952 ( .A(n7436), .B(n7437), .Z(n7439) );
  XNOR U7953 ( .A(n7438), .B(n7439), .Z(n7599) );
  XNOR U7954 ( .A(n7600), .B(n7599), .Z(n7601) );
  XNOR U7955 ( .A(n7602), .B(n7601), .Z(n7432) );
  NANDN U7956 ( .A(n17145), .B(o[29]), .Z(n7430) );
  OR U7957 ( .A(n7371), .B(n7370), .Z(n7375) );
  OR U7958 ( .A(n7373), .B(n7372), .Z(n7374) );
  NAND U7959 ( .A(n7375), .B(n7374), .Z(n7431) );
  XOR U7960 ( .A(n7430), .B(n7431), .Z(n7433) );
  XNOR U7961 ( .A(n7432), .B(n7433), .Z(n7605) );
  XNOR U7962 ( .A(n7606), .B(n7605), .Z(n7607) );
  XNOR U7963 ( .A(n7608), .B(n7607), .Z(n7426) );
  NANDN U7964 ( .A(n17219), .B(o[31]), .Z(n7424) );
  OR U7965 ( .A(n7377), .B(n7376), .Z(n7381) );
  OR U7966 ( .A(n7379), .B(n7378), .Z(n7380) );
  NAND U7967 ( .A(n7381), .B(n7380), .Z(n7425) );
  XOR U7968 ( .A(n7424), .B(n7425), .Z(n7427) );
  XNOR U7969 ( .A(n7426), .B(n7427), .Z(n7611) );
  XNOR U7970 ( .A(n7612), .B(n7611), .Z(n7613) );
  XNOR U7971 ( .A(n7614), .B(n7613), .Z(n7420) );
  NANDN U7972 ( .A(n17296), .B(o[33]), .Z(n7418) );
  OR U7973 ( .A(n7383), .B(n7382), .Z(n7387) );
  OR U7974 ( .A(n7385), .B(n7384), .Z(n7386) );
  NAND U7975 ( .A(n7387), .B(n7386), .Z(n7419) );
  XOR U7976 ( .A(n7418), .B(n7419), .Z(n7421) );
  XNOR U7977 ( .A(n7420), .B(n7421), .Z(n7617) );
  XNOR U7978 ( .A(n7618), .B(n7617), .Z(n7619) );
  XNOR U7979 ( .A(n7620), .B(n7619), .Z(n7414) );
  NANDN U7980 ( .A(n17375), .B(o[35]), .Z(n7412) );
  OR U7981 ( .A(n7389), .B(n7388), .Z(n7393) );
  OR U7982 ( .A(n7391), .B(n7390), .Z(n7392) );
  NAND U7983 ( .A(n7393), .B(n7392), .Z(n7413) );
  XOR U7984 ( .A(n7412), .B(n7413), .Z(n7415) );
  XNOR U7985 ( .A(n7414), .B(n7415), .Z(n7623) );
  XNOR U7986 ( .A(n7624), .B(n7623), .Z(n7625) );
  AND U7987 ( .A(o[37]), .B(\stack[1][1] ), .Z(n7406) );
  OR U7988 ( .A(n7395), .B(n7394), .Z(n7399) );
  OR U7989 ( .A(n7397), .B(n7396), .Z(n7398) );
  NAND U7990 ( .A(n7399), .B(n7398), .Z(n7407) );
  XNOR U7991 ( .A(n7406), .B(n7407), .Z(n7409) );
  XOR U7992 ( .A(n7408), .B(n7409), .Z(n7400) );
  NANDN U7993 ( .A(n7401), .B(n7400), .Z(n7403) );
  XOR U7994 ( .A(n7401), .B(n7400), .Z(n16014) );
  AND U7995 ( .A(o[38]), .B(\stack[1][0] ), .Z(n16015) );
  OR U7996 ( .A(n16014), .B(n16015), .Z(n7402) );
  AND U7997 ( .A(n7403), .B(n7402), .Z(n7405) );
  OR U7998 ( .A(n7404), .B(n7405), .Z(n7630) );
  XNOR U7999 ( .A(n7405), .B(n7404), .Z(n15976) );
  NANDN U8000 ( .A(n2969), .B(o[38]), .Z(n7851) );
  OR U8001 ( .A(n7407), .B(n7406), .Z(n7411) );
  OR U8002 ( .A(n7409), .B(n7408), .Z(n7410) );
  NAND U8003 ( .A(n7411), .B(n7410), .Z(n7849) );
  NANDN U8004 ( .A(n17375), .B(o[36]), .Z(n7845) );
  NANDN U8005 ( .A(n7413), .B(n7412), .Z(n7417) );
  NANDN U8006 ( .A(n7415), .B(n7414), .Z(n7416) );
  NAND U8007 ( .A(n7417), .B(n7416), .Z(n7843) );
  NANDN U8008 ( .A(n17296), .B(o[34]), .Z(n7839) );
  NANDN U8009 ( .A(n7419), .B(n7418), .Z(n7423) );
  NANDN U8010 ( .A(n7421), .B(n7420), .Z(n7422) );
  NAND U8011 ( .A(n7423), .B(n7422), .Z(n7837) );
  NANDN U8012 ( .A(n17219), .B(o[32]), .Z(n7833) );
  NANDN U8013 ( .A(n7425), .B(n7424), .Z(n7429) );
  NANDN U8014 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U8015 ( .A(n7429), .B(n7428), .Z(n7831) );
  NANDN U8016 ( .A(n17145), .B(o[30]), .Z(n7827) );
  NANDN U8017 ( .A(n7431), .B(n7430), .Z(n7435) );
  NANDN U8018 ( .A(n7433), .B(n7432), .Z(n7434) );
  NAND U8019 ( .A(n7435), .B(n7434), .Z(n7825) );
  NANDN U8020 ( .A(n2972), .B(o[28]), .Z(n7821) );
  NANDN U8021 ( .A(n7437), .B(n7436), .Z(n7441) );
  NANDN U8022 ( .A(n7439), .B(n7438), .Z(n7440) );
  NAND U8023 ( .A(n7441), .B(n7440), .Z(n7819) );
  AND U8024 ( .A(o[26]), .B(\stack[1][13] ), .Z(n7670) );
  OR U8025 ( .A(n7443), .B(n7442), .Z(n7447) );
  OR U8026 ( .A(n7445), .B(n7444), .Z(n7446) );
  AND U8027 ( .A(n7447), .B(n7446), .Z(n7667) );
  OR U8028 ( .A(n7449), .B(n7448), .Z(n7453) );
  NANDN U8029 ( .A(n7451), .B(n7450), .Z(n7452) );
  AND U8030 ( .A(n7453), .B(n7452), .Z(n7812) );
  AND U8031 ( .A(o[25]), .B(\stack[1][14] ), .Z(n7813) );
  XNOR U8032 ( .A(n7812), .B(n7813), .Z(n7815) );
  OR U8033 ( .A(n7455), .B(n7454), .Z(n7459) );
  OR U8034 ( .A(n7457), .B(n7456), .Z(n7458) );
  NAND U8035 ( .A(n7459), .B(n7458), .Z(n7680) );
  ANDN U8036 ( .B(\stack[1][16] ), .A(n3017), .Z(n7679) );
  XOR U8037 ( .A(n7680), .B(n7679), .Z(n7681) );
  NANDN U8038 ( .A(n16826), .B(o[22]), .Z(n7809) );
  OR U8039 ( .A(n7461), .B(n7460), .Z(n7465) );
  OR U8040 ( .A(n7463), .B(n7462), .Z(n7464) );
  NAND U8041 ( .A(n7465), .B(n7464), .Z(n7807) );
  AND U8042 ( .A(o[20]), .B(\stack[1][19] ), .Z(n7803) );
  OR U8043 ( .A(n7466), .B(n16747), .Z(n7470) );
  OR U8044 ( .A(n7468), .B(n7467), .Z(n7469) );
  AND U8045 ( .A(n7470), .B(n7469), .Z(n7800) );
  OR U8046 ( .A(n7472), .B(n7471), .Z(n7476) );
  NANDN U8047 ( .A(n7474), .B(n7473), .Z(n7475) );
  AND U8048 ( .A(n7476), .B(n7475), .Z(n7691) );
  AND U8049 ( .A(\stack[1][20] ), .B(o[19]), .Z(n7692) );
  XNOR U8050 ( .A(n7691), .B(n7692), .Z(n7694) );
  NANDN U8051 ( .A(n7478), .B(n7477), .Z(n7482) );
  OR U8052 ( .A(n7480), .B(n7479), .Z(n7481) );
  NAND U8053 ( .A(n7482), .B(n7481), .Z(n7698) );
  ANDN U8054 ( .B(o[17]), .A(n2979), .Z(n7697) );
  XNOR U8055 ( .A(n7698), .B(n7697), .Z(n7699) );
  NANDN U8056 ( .A(n3010), .B(\stack[1][23] ), .Z(n7791) );
  NANDN U8057 ( .A(n7484), .B(n7483), .Z(n7488) );
  NANDN U8058 ( .A(n7486), .B(n7485), .Z(n7487) );
  AND U8059 ( .A(n7488), .B(n7487), .Z(n7788) );
  NANDN U8060 ( .A(n3008), .B(\stack[1][25] ), .Z(n7785) );
  NANDN U8061 ( .A(n7490), .B(n7489), .Z(n7494) );
  NANDN U8062 ( .A(n7492), .B(n7491), .Z(n7493) );
  NAND U8063 ( .A(n7494), .B(n7493), .Z(n7783) );
  NANDN U8064 ( .A(n3006), .B(\stack[1][27] ), .Z(n7779) );
  NANDN U8065 ( .A(n7496), .B(n7495), .Z(n7500) );
  NANDN U8066 ( .A(n7498), .B(n7497), .Z(n7499) );
  NAND U8067 ( .A(n7500), .B(n7499), .Z(n7777) );
  NANDN U8068 ( .A(n3004), .B(\stack[1][29] ), .Z(n7724) );
  NANDN U8069 ( .A(n7502), .B(n7501), .Z(n7506) );
  NANDN U8070 ( .A(n7504), .B(n7503), .Z(n7505) );
  NAND U8071 ( .A(n7506), .B(n7505), .Z(n7722) );
  NANDN U8072 ( .A(n3002), .B(\stack[1][31] ), .Z(n7773) );
  OR U8073 ( .A(n7508), .B(n7507), .Z(n7512) );
  OR U8074 ( .A(n7510), .B(n7509), .Z(n7511) );
  NAND U8075 ( .A(n7512), .B(n7511), .Z(n7771) );
  OR U8076 ( .A(n7514), .B(n7513), .Z(n7518) );
  NANDN U8077 ( .A(n7516), .B(n7515), .Z(n7517) );
  AND U8078 ( .A(n7518), .B(n7517), .Z(n7733) );
  AND U8079 ( .A(\stack[1][32] ), .B(o[7]), .Z(n7734) );
  XNOR U8080 ( .A(n7733), .B(n7734), .Z(n7736) );
  OR U8081 ( .A(n7520), .B(n7519), .Z(n7524) );
  OR U8082 ( .A(n7522), .B(n7521), .Z(n7523) );
  AND U8083 ( .A(n7524), .B(n7523), .Z(n7739) );
  OR U8084 ( .A(n7526), .B(n7525), .Z(n7530) );
  OR U8085 ( .A(n7528), .B(n7527), .Z(n7529) );
  NAND U8086 ( .A(n7530), .B(n7529), .Z(n7746) );
  NANDN U8087 ( .A(n7532), .B(n7531), .Z(n7538) );
  ANDN U8088 ( .B(\stack[1][36] ), .A(n2994), .Z(n7534) );
  NAND U8089 ( .A(n7534), .B(n7533), .Z(n7536) );
  NANDN U8090 ( .A(n2993), .B(o[2]), .Z(n7535) );
  AND U8091 ( .A(n7536), .B(n7535), .Z(n7537) );
  ANDN U8092 ( .B(n7538), .A(n7537), .Z(n7751) );
  AND U8093 ( .A(\stack[1][36] ), .B(o[3]), .Z(n7752) );
  XNOR U8094 ( .A(n7751), .B(n7752), .Z(n7754) );
  ANDN U8095 ( .B(\stack[1][39] ), .A(n2994), .Z(n7761) );
  ANDN U8096 ( .B(\stack[1][38] ), .A(n2995), .Z(n7539) );
  XNOR U8097 ( .A(n7761), .B(n7539), .Z(n7541) );
  AND U8098 ( .A(n7540), .B(n7539), .Z(n7543) );
  ANDN U8099 ( .B(n7541), .A(n7543), .Z(n7759) );
  AND U8100 ( .A(\stack[1][39] ), .B(o[1]), .Z(n7762) );
  NAND U8101 ( .A(n7542), .B(n7762), .Z(n7983) );
  NAND U8102 ( .A(n7543), .B(n7983), .Z(n7544) );
  NANDN U8103 ( .A(n7759), .B(n7544), .Z(n7758) );
  AND U8104 ( .A(\stack[1][37] ), .B(o[2]), .Z(n7757) );
  XNOR U8105 ( .A(n7758), .B(n7757), .Z(n7753) );
  XOR U8106 ( .A(n7746), .B(n7745), .Z(n7748) );
  AND U8107 ( .A(\stack[1][35] ), .B(o[4]), .Z(n7747) );
  XNOR U8108 ( .A(n7748), .B(n7747), .Z(n7766) );
  AND U8109 ( .A(\stack[1][34] ), .B(o[5]), .Z(n7764) );
  OR U8110 ( .A(n7546), .B(n7545), .Z(n7550) );
  NANDN U8111 ( .A(n7548), .B(n7547), .Z(n7549) );
  NAND U8112 ( .A(n7550), .B(n7549), .Z(n7765) );
  XNOR U8113 ( .A(n7764), .B(n7765), .Z(n7767) );
  XNOR U8114 ( .A(n7766), .B(n7767), .Z(n7740) );
  XOR U8115 ( .A(n7739), .B(n7740), .Z(n7741) );
  AND U8116 ( .A(\stack[1][33] ), .B(o[6]), .Z(n7742) );
  XOR U8117 ( .A(n7741), .B(n7742), .Z(n7735) );
  XOR U8118 ( .A(n7736), .B(n7735), .Z(n7770) );
  XNOR U8119 ( .A(n7771), .B(n7770), .Z(n7772) );
  XNOR U8120 ( .A(n7773), .B(n7772), .Z(n7729) );
  NANDN U8121 ( .A(n2987), .B(o[9]), .Z(n7727) );
  OR U8122 ( .A(n7552), .B(n7551), .Z(n7556) );
  OR U8123 ( .A(n7554), .B(n7553), .Z(n7555) );
  NAND U8124 ( .A(n7556), .B(n7555), .Z(n7728) );
  XOR U8125 ( .A(n7727), .B(n7728), .Z(n7730) );
  XNOR U8126 ( .A(n7729), .B(n7730), .Z(n7721) );
  XNOR U8127 ( .A(n7722), .B(n7721), .Z(n7723) );
  XNOR U8128 ( .A(n7724), .B(n7723), .Z(n7717) );
  NANDN U8129 ( .A(n2985), .B(o[11]), .Z(n7715) );
  OR U8130 ( .A(n7558), .B(n7557), .Z(n7562) );
  OR U8131 ( .A(n7560), .B(n7559), .Z(n7561) );
  NAND U8132 ( .A(n7562), .B(n7561), .Z(n7716) );
  XOR U8133 ( .A(n7715), .B(n7716), .Z(n7718) );
  XNOR U8134 ( .A(n7717), .B(n7718), .Z(n7776) );
  XNOR U8135 ( .A(n7777), .B(n7776), .Z(n7778) );
  XNOR U8136 ( .A(n7779), .B(n7778), .Z(n7711) );
  NANDN U8137 ( .A(n2983), .B(o[13]), .Z(n7709) );
  OR U8138 ( .A(n7564), .B(n7563), .Z(n7568) );
  OR U8139 ( .A(n7566), .B(n7565), .Z(n7567) );
  NAND U8140 ( .A(n7568), .B(n7567), .Z(n7710) );
  XOR U8141 ( .A(n7709), .B(n7710), .Z(n7712) );
  XNOR U8142 ( .A(n7711), .B(n7712), .Z(n7782) );
  XNOR U8143 ( .A(n7783), .B(n7782), .Z(n7784) );
  XNOR U8144 ( .A(n7785), .B(n7784), .Z(n7705) );
  NANDN U8145 ( .A(n2981), .B(o[15]), .Z(n7703) );
  OR U8146 ( .A(n7570), .B(n7569), .Z(n7574) );
  OR U8147 ( .A(n7572), .B(n7571), .Z(n7573) );
  NAND U8148 ( .A(n7574), .B(n7573), .Z(n7704) );
  XOR U8149 ( .A(n7703), .B(n7704), .Z(n7706) );
  XNOR U8150 ( .A(n7705), .B(n7706), .Z(n7789) );
  XNOR U8151 ( .A(n7788), .B(n7789), .Z(n7790) );
  XOR U8152 ( .A(n7699), .B(n7700), .Z(n7794) );
  OR U8153 ( .A(n7576), .B(n7575), .Z(n7580) );
  NANDN U8154 ( .A(n7578), .B(n7577), .Z(n7579) );
  AND U8155 ( .A(n7580), .B(n7579), .Z(n7795) );
  XOR U8156 ( .A(n7794), .B(n7795), .Z(n7797) );
  AND U8157 ( .A(\stack[1][21] ), .B(o[18]), .Z(n7796) );
  XOR U8158 ( .A(n7797), .B(n7796), .Z(n7693) );
  XOR U8159 ( .A(n7694), .B(n7693), .Z(n7801) );
  XOR U8160 ( .A(n7800), .B(n7801), .Z(n7802) );
  XOR U8161 ( .A(n7803), .B(n7802), .Z(n7688) );
  NANDN U8162 ( .A(n3015), .B(\stack[1][18] ), .Z(n7685) );
  NANDN U8163 ( .A(n7582), .B(n7581), .Z(n7586) );
  NANDN U8164 ( .A(n7584), .B(n7583), .Z(n7585) );
  NAND U8165 ( .A(n7586), .B(n7585), .Z(n7686) );
  XOR U8166 ( .A(n7685), .B(n7686), .Z(n7687) );
  XNOR U8167 ( .A(n7688), .B(n7687), .Z(n7806) );
  XOR U8168 ( .A(n7807), .B(n7806), .Z(n7808) );
  XNOR U8169 ( .A(n7809), .B(n7808), .Z(n7682) );
  OR U8170 ( .A(n7588), .B(n7587), .Z(n7592) );
  OR U8171 ( .A(n7590), .B(n7589), .Z(n7591) );
  AND U8172 ( .A(n7592), .B(n7591), .Z(n7674) );
  XNOR U8173 ( .A(n7673), .B(n7674), .Z(n7676) );
  AND U8174 ( .A(o[24]), .B(\stack[1][15] ), .Z(n7675) );
  XOR U8175 ( .A(n7676), .B(n7675), .Z(n7814) );
  XOR U8176 ( .A(n7815), .B(n7814), .Z(n7668) );
  XOR U8177 ( .A(n7667), .B(n7668), .Z(n7669) );
  XOR U8178 ( .A(n7670), .B(n7669), .Z(n7664) );
  AND U8179 ( .A(o[27]), .B(\stack[1][12] ), .Z(n7661) );
  OR U8180 ( .A(n7594), .B(n7593), .Z(n7598) );
  OR U8181 ( .A(n7596), .B(n7595), .Z(n7597) );
  NAND U8182 ( .A(n7598), .B(n7597), .Z(n7662) );
  XNOR U8183 ( .A(n7661), .B(n7662), .Z(n7663) );
  XOR U8184 ( .A(n7664), .B(n7663), .Z(n7818) );
  XNOR U8185 ( .A(n7819), .B(n7818), .Z(n7820) );
  XNOR U8186 ( .A(n7821), .B(n7820), .Z(n7657) );
  NANDN U8187 ( .A(n17101), .B(o[29]), .Z(n7655) );
  OR U8188 ( .A(n7600), .B(n7599), .Z(n7604) );
  OR U8189 ( .A(n7602), .B(n7601), .Z(n7603) );
  NAND U8190 ( .A(n7604), .B(n7603), .Z(n7656) );
  XOR U8191 ( .A(n7655), .B(n7656), .Z(n7658) );
  XNOR U8192 ( .A(n7657), .B(n7658), .Z(n7824) );
  XNOR U8193 ( .A(n7825), .B(n7824), .Z(n7826) );
  XNOR U8194 ( .A(n7827), .B(n7826), .Z(n7651) );
  NANDN U8195 ( .A(n17179), .B(o[31]), .Z(n7649) );
  OR U8196 ( .A(n7606), .B(n7605), .Z(n7610) );
  OR U8197 ( .A(n7608), .B(n7607), .Z(n7609) );
  NAND U8198 ( .A(n7610), .B(n7609), .Z(n7650) );
  XOR U8199 ( .A(n7649), .B(n7650), .Z(n7652) );
  XNOR U8200 ( .A(n7651), .B(n7652), .Z(n7830) );
  XNOR U8201 ( .A(n7831), .B(n7830), .Z(n7832) );
  XNOR U8202 ( .A(n7833), .B(n7832), .Z(n7645) );
  NANDN U8203 ( .A(n17256), .B(o[33]), .Z(n7643) );
  OR U8204 ( .A(n7612), .B(n7611), .Z(n7616) );
  OR U8205 ( .A(n7614), .B(n7613), .Z(n7615) );
  NAND U8206 ( .A(n7616), .B(n7615), .Z(n7644) );
  XOR U8207 ( .A(n7643), .B(n7644), .Z(n7646) );
  XNOR U8208 ( .A(n7645), .B(n7646), .Z(n7836) );
  XNOR U8209 ( .A(n7837), .B(n7836), .Z(n7838) );
  XNOR U8210 ( .A(n7839), .B(n7838), .Z(n7639) );
  AND U8211 ( .A(o[35]), .B(\stack[1][4] ), .Z(n7637) );
  OR U8212 ( .A(n7618), .B(n7617), .Z(n7622) );
  OR U8213 ( .A(n7620), .B(n7619), .Z(n7621) );
  NAND U8214 ( .A(n7622), .B(n7621), .Z(n7638) );
  XNOR U8215 ( .A(n7637), .B(n7638), .Z(n7640) );
  XNOR U8216 ( .A(n7639), .B(n7640), .Z(n7842) );
  XNOR U8217 ( .A(n7843), .B(n7842), .Z(n7844) );
  XOR U8218 ( .A(n7845), .B(n7844), .Z(n7634) );
  AND U8219 ( .A(o[37]), .B(\stack[1][2] ), .Z(n7631) );
  OR U8220 ( .A(n7624), .B(n7623), .Z(n7628) );
  OR U8221 ( .A(n7626), .B(n7625), .Z(n7627) );
  NAND U8222 ( .A(n7628), .B(n7627), .Z(n7632) );
  XOR U8223 ( .A(n7631), .B(n7632), .Z(n7633) );
  XNOR U8224 ( .A(n7634), .B(n7633), .Z(n7848) );
  XNOR U8225 ( .A(n7849), .B(n7848), .Z(n7850) );
  XOR U8226 ( .A(n7851), .B(n7850), .Z(n15977) );
  OR U8227 ( .A(n15976), .B(n15977), .Z(n7629) );
  AND U8228 ( .A(n7630), .B(n7629), .Z(n7855) );
  NANDN U8229 ( .A(n2970), .B(o[38]), .Z(n8089) );
  OR U8230 ( .A(n7632), .B(n7631), .Z(n7636) );
  NANDN U8231 ( .A(n7634), .B(n7633), .Z(n7635) );
  NAND U8232 ( .A(n7636), .B(n7635), .Z(n8087) );
  NANDN U8233 ( .A(n2971), .B(o[36]), .Z(n8083) );
  OR U8234 ( .A(n7638), .B(n7637), .Z(n7642) );
  NANDN U8235 ( .A(n7640), .B(n7639), .Z(n7641) );
  NAND U8236 ( .A(n7642), .B(n7641), .Z(n8081) );
  NANDN U8237 ( .A(n17256), .B(o[34]), .Z(n8077) );
  NANDN U8238 ( .A(n7644), .B(n7643), .Z(n7648) );
  NANDN U8239 ( .A(n7646), .B(n7645), .Z(n7647) );
  NAND U8240 ( .A(n7648), .B(n7647), .Z(n8075) );
  NANDN U8241 ( .A(n17179), .B(o[32]), .Z(n8071) );
  NANDN U8242 ( .A(n7650), .B(n7649), .Z(n7654) );
  NANDN U8243 ( .A(n7652), .B(n7651), .Z(n7653) );
  NAND U8244 ( .A(n7654), .B(n7653), .Z(n8069) );
  NANDN U8245 ( .A(n17101), .B(o[30]), .Z(n8065) );
  NANDN U8246 ( .A(n7656), .B(n7655), .Z(n7660) );
  NANDN U8247 ( .A(n7658), .B(n7657), .Z(n7659) );
  NAND U8248 ( .A(n7660), .B(n7659), .Z(n8063) );
  AND U8249 ( .A(o[28]), .B(\stack[1][12] ), .Z(n8059) );
  OR U8250 ( .A(n7662), .B(n7661), .Z(n7666) );
  OR U8251 ( .A(n7664), .B(n7663), .Z(n7665) );
  AND U8252 ( .A(n7666), .B(n7665), .Z(n8056) );
  OR U8253 ( .A(n7668), .B(n7667), .Z(n7672) );
  NANDN U8254 ( .A(n7670), .B(n7669), .Z(n7671) );
  AND U8255 ( .A(n7672), .B(n7671), .Z(n7896) );
  AND U8256 ( .A(o[27]), .B(\stack[1][13] ), .Z(n7897) );
  XNOR U8257 ( .A(n7896), .B(n7897), .Z(n7899) );
  OR U8258 ( .A(n7674), .B(n7673), .Z(n7678) );
  OR U8259 ( .A(n7676), .B(n7675), .Z(n7677) );
  NAND U8260 ( .A(n7678), .B(n7677), .Z(n7903) );
  ANDN U8261 ( .B(\stack[1][15] ), .A(n3019), .Z(n7902) );
  XNOR U8262 ( .A(n7903), .B(n7902), .Z(n7904) );
  NANDN U8263 ( .A(n2977), .B(o[24]), .Z(n8047) );
  NANDN U8264 ( .A(n7680), .B(n7679), .Z(n7684) );
  OR U8265 ( .A(n7682), .B(n7681), .Z(n7683) );
  AND U8266 ( .A(n7684), .B(n7683), .Z(n8044) );
  NANDN U8267 ( .A(n16786), .B(o[22]), .Z(n8041) );
  NANDN U8268 ( .A(n7686), .B(n7685), .Z(n7690) );
  OR U8269 ( .A(n7688), .B(n7687), .Z(n7689) );
  NAND U8270 ( .A(n7690), .B(n7689), .Z(n8039) );
  NOR U8271 ( .A(n3014), .B(n16712), .Z(n8034) );
  OR U8272 ( .A(n7692), .B(n7691), .Z(n7696) );
  NANDN U8273 ( .A(n7694), .B(n7693), .Z(n7695) );
  NAND U8274 ( .A(n7696), .B(n7695), .Z(n8033) );
  NANDN U8275 ( .A(n3012), .B(\stack[1][22] ), .Z(n8029) );
  NANDN U8276 ( .A(n7698), .B(n7697), .Z(n7702) );
  NANDN U8277 ( .A(n7700), .B(n7699), .Z(n7701) );
  AND U8278 ( .A(n7702), .B(n7701), .Z(n8026) );
  NANDN U8279 ( .A(n3010), .B(\stack[1][24] ), .Z(n8023) );
  NANDN U8280 ( .A(n7704), .B(n7703), .Z(n7708) );
  NANDN U8281 ( .A(n7706), .B(n7705), .Z(n7707) );
  NAND U8282 ( .A(n7708), .B(n7707), .Z(n8021) );
  NANDN U8283 ( .A(n3008), .B(\stack[1][26] ), .Z(n8017) );
  NANDN U8284 ( .A(n7710), .B(n7709), .Z(n7714) );
  NANDN U8285 ( .A(n7712), .B(n7711), .Z(n7713) );
  NAND U8286 ( .A(n7714), .B(n7713), .Z(n8015) );
  AND U8287 ( .A(\stack[1][28] ), .B(o[12]), .Z(n7947) );
  NANDN U8288 ( .A(n7716), .B(n7715), .Z(n7720) );
  NANDN U8289 ( .A(n7718), .B(n7717), .Z(n7719) );
  AND U8290 ( .A(n7720), .B(n7719), .Z(n7944) );
  AND U8291 ( .A(\stack[1][29] ), .B(o[11]), .Z(n8008) );
  OR U8292 ( .A(n7722), .B(n7721), .Z(n7726) );
  OR U8293 ( .A(n7724), .B(n7723), .Z(n7725) );
  NAND U8294 ( .A(n7726), .B(n7725), .Z(n8009) );
  XNOR U8295 ( .A(n8008), .B(n8009), .Z(n8011) );
  NANDN U8296 ( .A(n7728), .B(n7727), .Z(n7732) );
  NANDN U8297 ( .A(n7730), .B(n7729), .Z(n7731) );
  AND U8298 ( .A(n7732), .B(n7731), .Z(n7950) );
  OR U8299 ( .A(n7734), .B(n7733), .Z(n7738) );
  OR U8300 ( .A(n7736), .B(n7735), .Z(n7737) );
  NAND U8301 ( .A(n7738), .B(n7737), .Z(n8003) );
  OR U8302 ( .A(n7740), .B(n7739), .Z(n7744) );
  NANDN U8303 ( .A(n7742), .B(n7741), .Z(n7743) );
  AND U8304 ( .A(n7744), .B(n7743), .Z(n7962) );
  AND U8305 ( .A(\stack[1][33] ), .B(o[7]), .Z(n7963) );
  XNOR U8306 ( .A(n7962), .B(n7963), .Z(n7965) );
  NANDN U8307 ( .A(n2999), .B(\stack[1][35] ), .Z(n7969) );
  NANDN U8308 ( .A(n7746), .B(n7745), .Z(n7750) );
  NANDN U8309 ( .A(n7748), .B(n7747), .Z(n7749) );
  AND U8310 ( .A(n7750), .B(n7749), .Z(n7968) );
  XNOR U8311 ( .A(n7969), .B(n7968), .Z(n7970) );
  OR U8312 ( .A(n7752), .B(n7751), .Z(n7756) );
  OR U8313 ( .A(n7754), .B(n7753), .Z(n7755) );
  NAND U8314 ( .A(n7756), .B(n7755), .Z(n7975) );
  OR U8315 ( .A(n7758), .B(n7757), .Z(n7760) );
  ANDN U8316 ( .B(n7760), .A(n7759), .Z(n7990) );
  AND U8317 ( .A(\stack[1][37] ), .B(o[3]), .Z(n7991) );
  XNOR U8318 ( .A(n7990), .B(n7991), .Z(n7993) );
  NANDN U8319 ( .A(n2996), .B(\stack[1][38] ), .Z(n7986) );
  AND U8320 ( .A(\stack[1][40] ), .B(o[1]), .Z(n7981) );
  AND U8321 ( .A(n7981), .B(n7761), .Z(n8233) );
  XOR U8322 ( .A(n8233), .B(n7983), .Z(n7763) );
  NAND U8323 ( .A(\stack[1][40] ), .B(o[0]), .Z(n7980) );
  NANDN U8324 ( .A(n7762), .B(n7980), .Z(n7985) );
  NAND U8325 ( .A(n7763), .B(n7985), .Z(n7987) );
  XOR U8326 ( .A(n7986), .B(n7987), .Z(n7992) );
  XOR U8327 ( .A(n7993), .B(n7992), .Z(n7974) );
  XNOR U8328 ( .A(n7975), .B(n7974), .Z(n7977) );
  NANDN U8329 ( .A(n2998), .B(\stack[1][36] ), .Z(n7976) );
  XNOR U8330 ( .A(n7977), .B(n7976), .Z(n7971) );
  OR U8331 ( .A(n7765), .B(n7764), .Z(n7769) );
  OR U8332 ( .A(n7767), .B(n7766), .Z(n7768) );
  AND U8333 ( .A(n7769), .B(n7768), .Z(n7997) );
  XNOR U8334 ( .A(n7996), .B(n7997), .Z(n7999) );
  AND U8335 ( .A(\stack[1][34] ), .B(o[6]), .Z(n7998) );
  XNOR U8336 ( .A(n7999), .B(n7998), .Z(n7964) );
  XOR U8337 ( .A(n8003), .B(n8002), .Z(n8005) );
  AND U8338 ( .A(\stack[1][32] ), .B(o[8]), .Z(n8004) );
  XNOR U8339 ( .A(n8005), .B(n8004), .Z(n7958) );
  AND U8340 ( .A(\stack[1][31] ), .B(o[9]), .Z(n7956) );
  OR U8341 ( .A(n7771), .B(n7770), .Z(n7775) );
  OR U8342 ( .A(n7773), .B(n7772), .Z(n7774) );
  NAND U8343 ( .A(n7775), .B(n7774), .Z(n7957) );
  XNOR U8344 ( .A(n7956), .B(n7957), .Z(n7959) );
  XNOR U8345 ( .A(n7958), .B(n7959), .Z(n7951) );
  XNOR U8346 ( .A(n7950), .B(n7951), .Z(n7952) );
  AND U8347 ( .A(\stack[1][30] ), .B(o[10]), .Z(n7953) );
  XNOR U8348 ( .A(n8011), .B(n8010), .Z(n7945) );
  XOR U8349 ( .A(n7944), .B(n7945), .Z(n7946) );
  XOR U8350 ( .A(n7947), .B(n7946), .Z(n7941) );
  AND U8351 ( .A(\stack[1][27] ), .B(o[13]), .Z(n7938) );
  OR U8352 ( .A(n7777), .B(n7776), .Z(n7781) );
  OR U8353 ( .A(n7779), .B(n7778), .Z(n7780) );
  NAND U8354 ( .A(n7781), .B(n7780), .Z(n7939) );
  XNOR U8355 ( .A(n7938), .B(n7939), .Z(n7940) );
  XOR U8356 ( .A(n7941), .B(n7940), .Z(n8014) );
  XNOR U8357 ( .A(n8015), .B(n8014), .Z(n8016) );
  XNOR U8358 ( .A(n8017), .B(n8016), .Z(n7934) );
  NANDN U8359 ( .A(n2982), .B(o[15]), .Z(n7932) );
  OR U8360 ( .A(n7783), .B(n7782), .Z(n7787) );
  OR U8361 ( .A(n7785), .B(n7784), .Z(n7786) );
  NAND U8362 ( .A(n7787), .B(n7786), .Z(n7933) );
  XOR U8363 ( .A(n7932), .B(n7933), .Z(n7935) );
  XNOR U8364 ( .A(n7934), .B(n7935), .Z(n8020) );
  XNOR U8365 ( .A(n8021), .B(n8020), .Z(n8022) );
  XOR U8366 ( .A(n8023), .B(n8022), .Z(n7928) );
  AND U8367 ( .A(\stack[1][23] ), .B(o[17]), .Z(n7926) );
  OR U8368 ( .A(n7789), .B(n7788), .Z(n7793) );
  OR U8369 ( .A(n7791), .B(n7790), .Z(n7792) );
  NAND U8370 ( .A(n7793), .B(n7792), .Z(n7927) );
  XNOR U8371 ( .A(n7926), .B(n7927), .Z(n7929) );
  XNOR U8372 ( .A(n8026), .B(n8027), .Z(n8028) );
  XNOR U8373 ( .A(n8029), .B(n8028), .Z(n7922) );
  NANDN U8374 ( .A(n7795), .B(n7794), .Z(n7799) );
  OR U8375 ( .A(n7797), .B(n7796), .Z(n7798) );
  AND U8376 ( .A(n7799), .B(n7798), .Z(n7921) );
  NANDN U8377 ( .A(n2978), .B(o[19]), .Z(n7920) );
  XOR U8378 ( .A(n7921), .B(n7920), .Z(n7923) );
  XNOR U8379 ( .A(n7922), .B(n7923), .Z(n8032) );
  XNOR U8380 ( .A(n8033), .B(n8032), .Z(n8035) );
  XOR U8381 ( .A(n8034), .B(n8035), .Z(n7916) );
  OR U8382 ( .A(n7801), .B(n7800), .Z(n7805) );
  NANDN U8383 ( .A(n7803), .B(n7802), .Z(n7804) );
  AND U8384 ( .A(n7805), .B(n7804), .Z(n7915) );
  NANDN U8385 ( .A(n3015), .B(\stack[1][19] ), .Z(n7914) );
  XOR U8386 ( .A(n7915), .B(n7914), .Z(n7917) );
  XNOR U8387 ( .A(n7916), .B(n7917), .Z(n8038) );
  XNOR U8388 ( .A(n8039), .B(n8038), .Z(n8040) );
  XNOR U8389 ( .A(n8041), .B(n8040), .Z(n7910) );
  NANDN U8390 ( .A(n3017), .B(\stack[1][17] ), .Z(n7908) );
  NANDN U8391 ( .A(n7807), .B(n7806), .Z(n7811) );
  OR U8392 ( .A(n7809), .B(n7808), .Z(n7810) );
  NAND U8393 ( .A(n7811), .B(n7810), .Z(n7909) );
  XOR U8394 ( .A(n7908), .B(n7909), .Z(n7911) );
  XNOR U8395 ( .A(n7910), .B(n7911), .Z(n8045) );
  XNOR U8396 ( .A(n8044), .B(n8045), .Z(n8046) );
  XOR U8397 ( .A(n7904), .B(n7905), .Z(n8050) );
  OR U8398 ( .A(n7813), .B(n7812), .Z(n7817) );
  NANDN U8399 ( .A(n7815), .B(n7814), .Z(n7816) );
  AND U8400 ( .A(n7817), .B(n7816), .Z(n8051) );
  XOR U8401 ( .A(n8050), .B(n8051), .Z(n8053) );
  AND U8402 ( .A(o[26]), .B(\stack[1][14] ), .Z(n8052) );
  XOR U8403 ( .A(n8053), .B(n8052), .Z(n7898) );
  XOR U8404 ( .A(n7899), .B(n7898), .Z(n8057) );
  XOR U8405 ( .A(n8056), .B(n8057), .Z(n8058) );
  XOR U8406 ( .A(n8059), .B(n8058), .Z(n7893) );
  AND U8407 ( .A(o[29]), .B(\stack[1][11] ), .Z(n7890) );
  OR U8408 ( .A(n7819), .B(n7818), .Z(n7823) );
  OR U8409 ( .A(n7821), .B(n7820), .Z(n7822) );
  NAND U8410 ( .A(n7823), .B(n7822), .Z(n7891) );
  XNOR U8411 ( .A(n7890), .B(n7891), .Z(n7892) );
  XOR U8412 ( .A(n7893), .B(n7892), .Z(n8062) );
  XNOR U8413 ( .A(n8063), .B(n8062), .Z(n8064) );
  XNOR U8414 ( .A(n8065), .B(n8064), .Z(n7886) );
  NANDN U8415 ( .A(n17145), .B(o[31]), .Z(n7884) );
  OR U8416 ( .A(n7825), .B(n7824), .Z(n7829) );
  OR U8417 ( .A(n7827), .B(n7826), .Z(n7828) );
  NAND U8418 ( .A(n7829), .B(n7828), .Z(n7885) );
  XOR U8419 ( .A(n7884), .B(n7885), .Z(n7887) );
  XNOR U8420 ( .A(n7886), .B(n7887), .Z(n8068) );
  XNOR U8421 ( .A(n8069), .B(n8068), .Z(n8070) );
  XNOR U8422 ( .A(n8071), .B(n8070), .Z(n7880) );
  NANDN U8423 ( .A(n17219), .B(o[33]), .Z(n7878) );
  OR U8424 ( .A(n7831), .B(n7830), .Z(n7835) );
  OR U8425 ( .A(n7833), .B(n7832), .Z(n7834) );
  NAND U8426 ( .A(n7835), .B(n7834), .Z(n7879) );
  XOR U8427 ( .A(n7878), .B(n7879), .Z(n7881) );
  XNOR U8428 ( .A(n7880), .B(n7881), .Z(n8074) );
  XNOR U8429 ( .A(n8075), .B(n8074), .Z(n8076) );
  XNOR U8430 ( .A(n8077), .B(n8076), .Z(n7874) );
  NANDN U8431 ( .A(n17296), .B(o[35]), .Z(n7872) );
  OR U8432 ( .A(n7837), .B(n7836), .Z(n7841) );
  OR U8433 ( .A(n7839), .B(n7838), .Z(n7840) );
  NAND U8434 ( .A(n7841), .B(n7840), .Z(n7873) );
  XOR U8435 ( .A(n7872), .B(n7873), .Z(n7875) );
  XNOR U8436 ( .A(n7874), .B(n7875), .Z(n8080) );
  XNOR U8437 ( .A(n8081), .B(n8080), .Z(n8082) );
  XNOR U8438 ( .A(n8083), .B(n8082), .Z(n7868) );
  NANDN U8439 ( .A(n17375), .B(o[37]), .Z(n7866) );
  OR U8440 ( .A(n7843), .B(n7842), .Z(n7847) );
  OR U8441 ( .A(n7845), .B(n7844), .Z(n7846) );
  NAND U8442 ( .A(n7847), .B(n7846), .Z(n7867) );
  XOR U8443 ( .A(n7866), .B(n7867), .Z(n7869) );
  XNOR U8444 ( .A(n7868), .B(n7869), .Z(n8086) );
  XNOR U8445 ( .A(n8087), .B(n8086), .Z(n8088) );
  AND U8446 ( .A(o[39]), .B(\stack[1][1] ), .Z(n7860) );
  OR U8447 ( .A(n7849), .B(n7848), .Z(n7853) );
  OR U8448 ( .A(n7851), .B(n7850), .Z(n7852) );
  NAND U8449 ( .A(n7853), .B(n7852), .Z(n7861) );
  XNOR U8450 ( .A(n7860), .B(n7861), .Z(n7863) );
  XOR U8451 ( .A(n7862), .B(n7863), .Z(n7854) );
  NANDN U8452 ( .A(n7855), .B(n7854), .Z(n7857) );
  XOR U8453 ( .A(n7855), .B(n7854), .Z(n15938) );
  AND U8454 ( .A(o[40]), .B(\stack[1][0] ), .Z(n15939) );
  OR U8455 ( .A(n15938), .B(n15939), .Z(n7856) );
  AND U8456 ( .A(n7857), .B(n7856), .Z(n7859) );
  OR U8457 ( .A(n7858), .B(n7859), .Z(n8093) );
  XNOR U8458 ( .A(n7859), .B(n7858), .Z(n15899) );
  NANDN U8459 ( .A(n2969), .B(o[40]), .Z(n8330) );
  OR U8460 ( .A(n7861), .B(n7860), .Z(n7865) );
  OR U8461 ( .A(n7863), .B(n7862), .Z(n7864) );
  NAND U8462 ( .A(n7865), .B(n7864), .Z(n8328) );
  NANDN U8463 ( .A(n17375), .B(o[38]), .Z(n8324) );
  NANDN U8464 ( .A(n7867), .B(n7866), .Z(n7871) );
  NANDN U8465 ( .A(n7869), .B(n7868), .Z(n7870) );
  NAND U8466 ( .A(n7871), .B(n7870), .Z(n8322) );
  NANDN U8467 ( .A(n17296), .B(o[36]), .Z(n8318) );
  NANDN U8468 ( .A(n7873), .B(n7872), .Z(n7877) );
  NANDN U8469 ( .A(n7875), .B(n7874), .Z(n7876) );
  NAND U8470 ( .A(n7877), .B(n7876), .Z(n8316) );
  NANDN U8471 ( .A(n17219), .B(o[34]), .Z(n8312) );
  NANDN U8472 ( .A(n7879), .B(n7878), .Z(n7883) );
  NANDN U8473 ( .A(n7881), .B(n7880), .Z(n7882) );
  NAND U8474 ( .A(n7883), .B(n7882), .Z(n8310) );
  NANDN U8475 ( .A(n17145), .B(o[32]), .Z(n8306) );
  NANDN U8476 ( .A(n7885), .B(n7884), .Z(n7889) );
  NANDN U8477 ( .A(n7887), .B(n7886), .Z(n7888) );
  NAND U8478 ( .A(n7889), .B(n7888), .Z(n8304) );
  NANDN U8479 ( .A(n2972), .B(o[30]), .Z(n8300) );
  OR U8480 ( .A(n7891), .B(n7890), .Z(n7895) );
  OR U8481 ( .A(n7893), .B(n7892), .Z(n7894) );
  NAND U8482 ( .A(n7895), .B(n7894), .Z(n8298) );
  NANDN U8483 ( .A(n2974), .B(o[28]), .Z(n8294) );
  OR U8484 ( .A(n7897), .B(n7896), .Z(n7901) );
  NANDN U8485 ( .A(n7899), .B(n7898), .Z(n7900) );
  NAND U8486 ( .A(n7901), .B(n7900), .Z(n8292) );
  NANDN U8487 ( .A(n2976), .B(o[26]), .Z(n8288) );
  NANDN U8488 ( .A(n7903), .B(n7902), .Z(n7907) );
  NANDN U8489 ( .A(n7905), .B(n7904), .Z(n7906) );
  AND U8490 ( .A(n7907), .B(n7906), .Z(n8285) );
  NANDN U8491 ( .A(n16826), .B(o[24]), .Z(n8145) );
  NANDN U8492 ( .A(n7909), .B(n7908), .Z(n7913) );
  NANDN U8493 ( .A(n7911), .B(n7910), .Z(n7912) );
  NAND U8494 ( .A(n7913), .B(n7912), .Z(n8143) );
  NANDN U8495 ( .A(n16746), .B(o[22]), .Z(n8282) );
  NANDN U8496 ( .A(n7915), .B(n7914), .Z(n7919) );
  NANDN U8497 ( .A(n7917), .B(n7916), .Z(n7918) );
  NAND U8498 ( .A(n7919), .B(n7918), .Z(n8280) );
  NANDN U8499 ( .A(n3014), .B(\stack[1][21] ), .Z(n8276) );
  NANDN U8500 ( .A(n7921), .B(n7920), .Z(n7925) );
  NANDN U8501 ( .A(n7923), .B(n7922), .Z(n7924) );
  NAND U8502 ( .A(n7925), .B(n7924), .Z(n8274) );
  NANDN U8503 ( .A(n3012), .B(\stack[1][23] ), .Z(n8270) );
  OR U8504 ( .A(n7927), .B(n7926), .Z(n7931) );
  OR U8505 ( .A(n7929), .B(n7928), .Z(n7930) );
  NAND U8506 ( .A(n7931), .B(n7930), .Z(n8268) );
  NANDN U8507 ( .A(n3010), .B(\stack[1][25] ), .Z(n8264) );
  NANDN U8508 ( .A(n7933), .B(n7932), .Z(n7937) );
  NANDN U8509 ( .A(n7935), .B(n7934), .Z(n7936) );
  NAND U8510 ( .A(n7937), .B(n7936), .Z(n8262) );
  AND U8511 ( .A(\stack[1][27] ), .B(o[14]), .Z(n8181) );
  OR U8512 ( .A(n7939), .B(n7938), .Z(n7943) );
  OR U8513 ( .A(n7941), .B(n7940), .Z(n7942) );
  AND U8514 ( .A(n7943), .B(n7942), .Z(n8178) );
  OR U8515 ( .A(n7945), .B(n7944), .Z(n7949) );
  NANDN U8516 ( .A(n7947), .B(n7946), .Z(n7948) );
  AND U8517 ( .A(n7949), .B(n7948), .Z(n8255) );
  AND U8518 ( .A(\stack[1][28] ), .B(o[13]), .Z(n8256) );
  XNOR U8519 ( .A(n8255), .B(n8256), .Z(n8258) );
  OR U8520 ( .A(n7951), .B(n7950), .Z(n7955) );
  OR U8521 ( .A(n7953), .B(n7952), .Z(n7954) );
  NAND U8522 ( .A(n7955), .B(n7954), .Z(n8191) );
  ANDN U8523 ( .B(o[11]), .A(n2987), .Z(n8190) );
  XOR U8524 ( .A(n8191), .B(n8190), .Z(n8192) );
  NANDN U8525 ( .A(n3004), .B(\stack[1][31] ), .Z(n8252) );
  OR U8526 ( .A(n7957), .B(n7956), .Z(n7961) );
  OR U8527 ( .A(n7959), .B(n7958), .Z(n7960) );
  NAND U8528 ( .A(n7961), .B(n7960), .Z(n8250) );
  NANDN U8529 ( .A(n3002), .B(\stack[1][33] ), .Z(n8205) );
  OR U8530 ( .A(n7963), .B(n7962), .Z(n7967) );
  OR U8531 ( .A(n7965), .B(n7964), .Z(n7966) );
  NAND U8532 ( .A(n7967), .B(n7966), .Z(n8203) );
  OR U8533 ( .A(n7969), .B(n7968), .Z(n7973) );
  OR U8534 ( .A(n7971), .B(n7970), .Z(n7972) );
  AND U8535 ( .A(n7973), .B(n7972), .Z(n8208) );
  AND U8536 ( .A(\stack[1][36] ), .B(o[5]), .Z(n8214) );
  OR U8537 ( .A(n7975), .B(n7974), .Z(n7979) );
  OR U8538 ( .A(n7977), .B(n7976), .Z(n7978) );
  NAND U8539 ( .A(n7979), .B(n7978), .Z(n8215) );
  XNOR U8540 ( .A(n8214), .B(n8215), .Z(n8217) );
  AND U8541 ( .A(\stack[1][37] ), .B(o[4]), .Z(n8223) );
  ANDN U8542 ( .B(\stack[1][38] ), .A(n2997), .Z(n8229) );
  AND U8543 ( .A(\stack[1][41] ), .B(o[1]), .Z(n8241) );
  NANDN U8544 ( .A(n7980), .B(n8241), .Z(n8232) );
  IV U8545 ( .A(n8232), .Z(n8470) );
  XNOR U8546 ( .A(n8470), .B(n8233), .Z(n7982) );
  NAND U8547 ( .A(\stack[1][41] ), .B(o[0]), .Z(n8240) );
  NANDN U8548 ( .A(n7981), .B(n8240), .Z(n8235) );
  NAND U8549 ( .A(n7982), .B(n8235), .Z(n8237) );
  AND U8550 ( .A(\stack[1][39] ), .B(o[2]), .Z(n8236) );
  XNOR U8551 ( .A(n8237), .B(n8236), .Z(n8227) );
  NAND U8552 ( .A(n7983), .B(n8233), .Z(n7984) );
  AND U8553 ( .A(n7985), .B(n7984), .Z(n7989) );
  NANDN U8554 ( .A(n7987), .B(n7986), .Z(n7988) );
  AND U8555 ( .A(n7989), .B(n7988), .Z(n8226) );
  XOR U8556 ( .A(n8227), .B(n8226), .Z(n8228) );
  XOR U8557 ( .A(n8229), .B(n8228), .Z(n8221) );
  OR U8558 ( .A(n7991), .B(n7990), .Z(n7995) );
  OR U8559 ( .A(n7993), .B(n7992), .Z(n7994) );
  AND U8560 ( .A(n7995), .B(n7994), .Z(n8220) );
  XOR U8561 ( .A(n8221), .B(n8220), .Z(n8222) );
  XOR U8562 ( .A(n8223), .B(n8222), .Z(n8216) );
  XOR U8563 ( .A(n8217), .B(n8216), .Z(n8209) );
  XNOR U8564 ( .A(n8208), .B(n8209), .Z(n8211) );
  ANDN U8565 ( .B(o[6]), .A(n2992), .Z(n8210) );
  XOR U8566 ( .A(n8211), .B(n8210), .Z(n8245) );
  OR U8567 ( .A(n7997), .B(n7996), .Z(n8001) );
  OR U8568 ( .A(n7999), .B(n7998), .Z(n8000) );
  AND U8569 ( .A(n8001), .B(n8000), .Z(n8244) );
  NANDN U8570 ( .A(n2991), .B(o[7]), .Z(n8243) );
  XOR U8571 ( .A(n8244), .B(n8243), .Z(n8246) );
  XNOR U8572 ( .A(n8245), .B(n8246), .Z(n8202) );
  XNOR U8573 ( .A(n8203), .B(n8202), .Z(n8204) );
  XNOR U8574 ( .A(n8205), .B(n8204), .Z(n8198) );
  AND U8575 ( .A(\stack[1][32] ), .B(o[9]), .Z(n8196) );
  NANDN U8576 ( .A(n8003), .B(n8002), .Z(n8007) );
  NANDN U8577 ( .A(n8005), .B(n8004), .Z(n8006) );
  NAND U8578 ( .A(n8007), .B(n8006), .Z(n8197) );
  XNOR U8579 ( .A(n8196), .B(n8197), .Z(n8199) );
  XNOR U8580 ( .A(n8198), .B(n8199), .Z(n8249) );
  XNOR U8581 ( .A(n8250), .B(n8249), .Z(n8251) );
  XNOR U8582 ( .A(n8252), .B(n8251), .Z(n8193) );
  OR U8583 ( .A(n8009), .B(n8008), .Z(n8013) );
  OR U8584 ( .A(n8011), .B(n8010), .Z(n8012) );
  AND U8585 ( .A(n8013), .B(n8012), .Z(n8185) );
  XNOR U8586 ( .A(n8184), .B(n8185), .Z(n8187) );
  AND U8587 ( .A(\stack[1][29] ), .B(o[12]), .Z(n8186) );
  XOR U8588 ( .A(n8187), .B(n8186), .Z(n8257) );
  XOR U8589 ( .A(n8258), .B(n8257), .Z(n8179) );
  XOR U8590 ( .A(n8178), .B(n8179), .Z(n8180) );
  XOR U8591 ( .A(n8181), .B(n8180), .Z(n8175) );
  AND U8592 ( .A(\stack[1][26] ), .B(o[15]), .Z(n8172) );
  OR U8593 ( .A(n8015), .B(n8014), .Z(n8019) );
  OR U8594 ( .A(n8017), .B(n8016), .Z(n8018) );
  NAND U8595 ( .A(n8019), .B(n8018), .Z(n8173) );
  XNOR U8596 ( .A(n8172), .B(n8173), .Z(n8174) );
  XOR U8597 ( .A(n8175), .B(n8174), .Z(n8261) );
  XNOR U8598 ( .A(n8262), .B(n8261), .Z(n8263) );
  XNOR U8599 ( .A(n8264), .B(n8263), .Z(n8168) );
  NANDN U8600 ( .A(n2981), .B(o[17]), .Z(n8166) );
  OR U8601 ( .A(n8021), .B(n8020), .Z(n8025) );
  OR U8602 ( .A(n8023), .B(n8022), .Z(n8024) );
  NAND U8603 ( .A(n8025), .B(n8024), .Z(n8167) );
  XOR U8604 ( .A(n8166), .B(n8167), .Z(n8169) );
  XNOR U8605 ( .A(n8168), .B(n8169), .Z(n8267) );
  XNOR U8606 ( .A(n8268), .B(n8267), .Z(n8269) );
  XNOR U8607 ( .A(n8270), .B(n8269), .Z(n8162) );
  NANDN U8608 ( .A(n2979), .B(o[19]), .Z(n8160) );
  OR U8609 ( .A(n8027), .B(n8026), .Z(n8031) );
  OR U8610 ( .A(n8029), .B(n8028), .Z(n8030) );
  NAND U8611 ( .A(n8031), .B(n8030), .Z(n8161) );
  XOR U8612 ( .A(n8160), .B(n8161), .Z(n8163) );
  XNOR U8613 ( .A(n8162), .B(n8163), .Z(n8273) );
  XNOR U8614 ( .A(n8274), .B(n8273), .Z(n8275) );
  XNOR U8615 ( .A(n8276), .B(n8275), .Z(n8156) );
  NANDN U8616 ( .A(n3015), .B(\stack[1][20] ), .Z(n8154) );
  OR U8617 ( .A(n8033), .B(n8032), .Z(n8037) );
  IV U8618 ( .A(n8034), .Z(n16706) );
  OR U8619 ( .A(n8035), .B(n16706), .Z(n8036) );
  NAND U8620 ( .A(n8037), .B(n8036), .Z(n8155) );
  XOR U8621 ( .A(n8154), .B(n8155), .Z(n8157) );
  XNOR U8622 ( .A(n8156), .B(n8157), .Z(n8279) );
  XNOR U8623 ( .A(n8280), .B(n8279), .Z(n8281) );
  XNOR U8624 ( .A(n8282), .B(n8281), .Z(n8150) );
  NANDN U8625 ( .A(n3017), .B(\stack[1][18] ), .Z(n8148) );
  OR U8626 ( .A(n8039), .B(n8038), .Z(n8043) );
  OR U8627 ( .A(n8041), .B(n8040), .Z(n8042) );
  NAND U8628 ( .A(n8043), .B(n8042), .Z(n8149) );
  XOR U8629 ( .A(n8148), .B(n8149), .Z(n8151) );
  XNOR U8630 ( .A(n8150), .B(n8151), .Z(n8142) );
  XNOR U8631 ( .A(n8143), .B(n8142), .Z(n8144) );
  XOR U8632 ( .A(n8145), .B(n8144), .Z(n8138) );
  AND U8633 ( .A(o[25]), .B(\stack[1][16] ), .Z(n8136) );
  OR U8634 ( .A(n8045), .B(n8044), .Z(n8049) );
  OR U8635 ( .A(n8047), .B(n8046), .Z(n8048) );
  NAND U8636 ( .A(n8049), .B(n8048), .Z(n8137) );
  XNOR U8637 ( .A(n8136), .B(n8137), .Z(n8139) );
  XNOR U8638 ( .A(n8285), .B(n8286), .Z(n8287) );
  XNOR U8639 ( .A(n8288), .B(n8287), .Z(n8132) );
  NANDN U8640 ( .A(n8051), .B(n8050), .Z(n8055) );
  OR U8641 ( .A(n8053), .B(n8052), .Z(n8054) );
  AND U8642 ( .A(n8055), .B(n8054), .Z(n8131) );
  NANDN U8643 ( .A(n2975), .B(o[27]), .Z(n8130) );
  XOR U8644 ( .A(n8131), .B(n8130), .Z(n8133) );
  XNOR U8645 ( .A(n8132), .B(n8133), .Z(n8291) );
  XNOR U8646 ( .A(n8292), .B(n8291), .Z(n8293) );
  XNOR U8647 ( .A(n8294), .B(n8293), .Z(n8126) );
  OR U8648 ( .A(n8057), .B(n8056), .Z(n8061) );
  NANDN U8649 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U8650 ( .A(n8061), .B(n8060), .Z(n8125) );
  NANDN U8651 ( .A(n2973), .B(o[29]), .Z(n8124) );
  XOR U8652 ( .A(n8125), .B(n8124), .Z(n8127) );
  XNOR U8653 ( .A(n8126), .B(n8127), .Z(n8297) );
  XNOR U8654 ( .A(n8298), .B(n8297), .Z(n8299) );
  XNOR U8655 ( .A(n8300), .B(n8299), .Z(n8120) );
  NANDN U8656 ( .A(n17101), .B(o[31]), .Z(n8118) );
  OR U8657 ( .A(n8063), .B(n8062), .Z(n8067) );
  OR U8658 ( .A(n8065), .B(n8064), .Z(n8066) );
  NAND U8659 ( .A(n8067), .B(n8066), .Z(n8119) );
  XOR U8660 ( .A(n8118), .B(n8119), .Z(n8121) );
  XNOR U8661 ( .A(n8120), .B(n8121), .Z(n8303) );
  XNOR U8662 ( .A(n8304), .B(n8303), .Z(n8305) );
  XNOR U8663 ( .A(n8306), .B(n8305), .Z(n8114) );
  NANDN U8664 ( .A(n17179), .B(o[33]), .Z(n8112) );
  OR U8665 ( .A(n8069), .B(n8068), .Z(n8073) );
  OR U8666 ( .A(n8071), .B(n8070), .Z(n8072) );
  NAND U8667 ( .A(n8073), .B(n8072), .Z(n8113) );
  XOR U8668 ( .A(n8112), .B(n8113), .Z(n8115) );
  XNOR U8669 ( .A(n8114), .B(n8115), .Z(n8309) );
  XNOR U8670 ( .A(n8310), .B(n8309), .Z(n8311) );
  XNOR U8671 ( .A(n8312), .B(n8311), .Z(n8108) );
  NANDN U8672 ( .A(n17256), .B(o[35]), .Z(n8106) );
  OR U8673 ( .A(n8075), .B(n8074), .Z(n8079) );
  OR U8674 ( .A(n8077), .B(n8076), .Z(n8078) );
  NAND U8675 ( .A(n8079), .B(n8078), .Z(n8107) );
  XOR U8676 ( .A(n8106), .B(n8107), .Z(n8109) );
  XNOR U8677 ( .A(n8108), .B(n8109), .Z(n8315) );
  XNOR U8678 ( .A(n8316), .B(n8315), .Z(n8317) );
  XNOR U8679 ( .A(n8318), .B(n8317), .Z(n8102) );
  AND U8680 ( .A(o[37]), .B(\stack[1][4] ), .Z(n8100) );
  OR U8681 ( .A(n8081), .B(n8080), .Z(n8085) );
  OR U8682 ( .A(n8083), .B(n8082), .Z(n8084) );
  NAND U8683 ( .A(n8085), .B(n8084), .Z(n8101) );
  XNOR U8684 ( .A(n8100), .B(n8101), .Z(n8103) );
  XNOR U8685 ( .A(n8102), .B(n8103), .Z(n8321) );
  XNOR U8686 ( .A(n8322), .B(n8321), .Z(n8323) );
  XOR U8687 ( .A(n8324), .B(n8323), .Z(n8097) );
  AND U8688 ( .A(o[39]), .B(\stack[1][2] ), .Z(n8094) );
  OR U8689 ( .A(n8087), .B(n8086), .Z(n8091) );
  OR U8690 ( .A(n8089), .B(n8088), .Z(n8090) );
  NAND U8691 ( .A(n8091), .B(n8090), .Z(n8095) );
  XOR U8692 ( .A(n8094), .B(n8095), .Z(n8096) );
  XNOR U8693 ( .A(n8097), .B(n8096), .Z(n8327) );
  XNOR U8694 ( .A(n8328), .B(n8327), .Z(n8329) );
  XOR U8695 ( .A(n8330), .B(n8329), .Z(n15900) );
  OR U8696 ( .A(n15899), .B(n15900), .Z(n8092) );
  AND U8697 ( .A(n8093), .B(n8092), .Z(n8334) );
  NANDN U8698 ( .A(n2970), .B(o[40]), .Z(n8580) );
  OR U8699 ( .A(n8095), .B(n8094), .Z(n8099) );
  NANDN U8700 ( .A(n8097), .B(n8096), .Z(n8098) );
  NAND U8701 ( .A(n8099), .B(n8098), .Z(n8578) );
  NANDN U8702 ( .A(n2971), .B(o[38]), .Z(n8574) );
  OR U8703 ( .A(n8101), .B(n8100), .Z(n8105) );
  NANDN U8704 ( .A(n8103), .B(n8102), .Z(n8104) );
  NAND U8705 ( .A(n8105), .B(n8104), .Z(n8572) );
  NANDN U8706 ( .A(n17256), .B(o[36]), .Z(n8568) );
  NANDN U8707 ( .A(n8107), .B(n8106), .Z(n8111) );
  NANDN U8708 ( .A(n8109), .B(n8108), .Z(n8110) );
  NAND U8709 ( .A(n8111), .B(n8110), .Z(n8566) );
  NANDN U8710 ( .A(n17179), .B(o[34]), .Z(n8562) );
  NANDN U8711 ( .A(n8113), .B(n8112), .Z(n8117) );
  NANDN U8712 ( .A(n8115), .B(n8114), .Z(n8116) );
  NAND U8713 ( .A(n8117), .B(n8116), .Z(n8560) );
  NANDN U8714 ( .A(n17101), .B(o[32]), .Z(n8556) );
  NANDN U8715 ( .A(n8119), .B(n8118), .Z(n8123) );
  NANDN U8716 ( .A(n8121), .B(n8120), .Z(n8122) );
  NAND U8717 ( .A(n8123), .B(n8122), .Z(n8554) );
  NANDN U8718 ( .A(n2973), .B(o[30]), .Z(n8550) );
  NANDN U8719 ( .A(n8125), .B(n8124), .Z(n8129) );
  NANDN U8720 ( .A(n8127), .B(n8126), .Z(n8128) );
  NAND U8721 ( .A(n8129), .B(n8128), .Z(n8548) );
  NANDN U8722 ( .A(n2975), .B(o[28]), .Z(n8544) );
  NANDN U8723 ( .A(n8131), .B(n8130), .Z(n8135) );
  NANDN U8724 ( .A(n8133), .B(n8132), .Z(n8134) );
  NAND U8725 ( .A(n8135), .B(n8134), .Z(n8542) );
  AND U8726 ( .A(o[26]), .B(\stack[1][16] ), .Z(n8390) );
  OR U8727 ( .A(n8137), .B(n8136), .Z(n8141) );
  OR U8728 ( .A(n8139), .B(n8138), .Z(n8140) );
  AND U8729 ( .A(n8141), .B(n8140), .Z(n8387) );
  AND U8730 ( .A(o[25]), .B(\stack[1][17] ), .Z(n8535) );
  OR U8731 ( .A(n8143), .B(n8142), .Z(n8147) );
  OR U8732 ( .A(n8145), .B(n8144), .Z(n8146) );
  NAND U8733 ( .A(n8147), .B(n8146), .Z(n8536) );
  XNOR U8734 ( .A(n8535), .B(n8536), .Z(n8538) );
  NANDN U8735 ( .A(n8149), .B(n8148), .Z(n8153) );
  NANDN U8736 ( .A(n8151), .B(n8150), .Z(n8152) );
  AND U8737 ( .A(n8153), .B(n8152), .Z(n8393) );
  NANDN U8738 ( .A(n8155), .B(n8154), .Z(n8159) );
  NANDN U8739 ( .A(n8157), .B(n8156), .Z(n8158) );
  NAND U8740 ( .A(n8159), .B(n8158), .Z(n8530) );
  NANDN U8741 ( .A(n3014), .B(\stack[1][22] ), .Z(n8526) );
  NANDN U8742 ( .A(n8161), .B(n8160), .Z(n8165) );
  NANDN U8743 ( .A(n8163), .B(n8162), .Z(n8164) );
  NAND U8744 ( .A(n8165), .B(n8164), .Z(n8524) );
  NANDN U8745 ( .A(n3012), .B(\stack[1][24] ), .Z(n8520) );
  NANDN U8746 ( .A(n8167), .B(n8166), .Z(n8171) );
  NANDN U8747 ( .A(n8169), .B(n8168), .Z(n8170) );
  NAND U8748 ( .A(n8171), .B(n8170), .Z(n8518) );
  AND U8749 ( .A(\stack[1][26] ), .B(o[16]), .Z(n8425) );
  OR U8750 ( .A(n8173), .B(n8172), .Z(n8177) );
  OR U8751 ( .A(n8175), .B(n8174), .Z(n8176) );
  AND U8752 ( .A(n8177), .B(n8176), .Z(n8422) );
  OR U8753 ( .A(n8179), .B(n8178), .Z(n8183) );
  NANDN U8754 ( .A(n8181), .B(n8180), .Z(n8182) );
  AND U8755 ( .A(n8183), .B(n8182), .Z(n8511) );
  AND U8756 ( .A(\stack[1][27] ), .B(o[15]), .Z(n8512) );
  XNOR U8757 ( .A(n8511), .B(n8512), .Z(n8514) );
  OR U8758 ( .A(n8185), .B(n8184), .Z(n8189) );
  OR U8759 ( .A(n8187), .B(n8186), .Z(n8188) );
  NAND U8760 ( .A(n8189), .B(n8188), .Z(n8435) );
  ANDN U8761 ( .B(o[13]), .A(n2986), .Z(n8434) );
  XNOR U8762 ( .A(n8435), .B(n8434), .Z(n8436) );
  NANDN U8763 ( .A(n3006), .B(\stack[1][30] ), .Z(n8508) );
  NANDN U8764 ( .A(n8191), .B(n8190), .Z(n8195) );
  OR U8765 ( .A(n8193), .B(n8192), .Z(n8194) );
  AND U8766 ( .A(n8195), .B(n8194), .Z(n8505) );
  NANDN U8767 ( .A(n3004), .B(\stack[1][32] ), .Z(n8502) );
  OR U8768 ( .A(n8197), .B(n8196), .Z(n8201) );
  NANDN U8769 ( .A(n8199), .B(n8198), .Z(n8200) );
  NAND U8770 ( .A(n8201), .B(n8200), .Z(n8500) );
  AND U8771 ( .A(\stack[1][33] ), .B(o[9]), .Z(n8446) );
  OR U8772 ( .A(n8203), .B(n8202), .Z(n8207) );
  OR U8773 ( .A(n8205), .B(n8204), .Z(n8206) );
  NAND U8774 ( .A(n8207), .B(n8206), .Z(n8447) );
  XNOR U8775 ( .A(n8446), .B(n8447), .Z(n8449) );
  NANDN U8776 ( .A(n3001), .B(\stack[1][35] ), .Z(n8494) );
  OR U8777 ( .A(n8209), .B(n8208), .Z(n8213) );
  NANDN U8778 ( .A(n8211), .B(n8210), .Z(n8212) );
  AND U8779 ( .A(n8213), .B(n8212), .Z(n8493) );
  XNOR U8780 ( .A(n8494), .B(n8493), .Z(n8495) );
  OR U8781 ( .A(n8215), .B(n8214), .Z(n8219) );
  OR U8782 ( .A(n8217), .B(n8216), .Z(n8218) );
  NAND U8783 ( .A(n8219), .B(n8218), .Z(n8488) );
  OR U8784 ( .A(n8221), .B(n8220), .Z(n8225) );
  NANDN U8785 ( .A(n8223), .B(n8222), .Z(n8224) );
  AND U8786 ( .A(n8225), .B(n8224), .Z(n8458) );
  AND U8787 ( .A(\stack[1][37] ), .B(o[5]), .Z(n8459) );
  XNOR U8788 ( .A(n8458), .B(n8459), .Z(n8461) );
  NANDN U8789 ( .A(n2998), .B(\stack[1][38] ), .Z(n8466) );
  OR U8790 ( .A(n8227), .B(n8226), .Z(n8231) );
  NANDN U8791 ( .A(n8229), .B(n8228), .Z(n8230) );
  AND U8792 ( .A(n8231), .B(n8230), .Z(n8465) );
  NANDN U8793 ( .A(n2997), .B(\stack[1][39] ), .Z(n8482) );
  OR U8794 ( .A(n8233), .B(n8232), .Z(n8234) );
  AND U8795 ( .A(n8235), .B(n8234), .Z(n8239) );
  OR U8796 ( .A(n8237), .B(n8236), .Z(n8238) );
  AND U8797 ( .A(n8239), .B(n8238), .Z(n8481) );
  AND U8798 ( .A(\stack[1][42] ), .B(o[1]), .Z(n8478) );
  ANDN U8799 ( .B(n8478), .A(n8240), .Z(n8729) );
  XNOR U8800 ( .A(n8729), .B(n8470), .Z(n8242) );
  NAND U8801 ( .A(\stack[1][42] ), .B(o[0]), .Z(n8477) );
  NANDN U8802 ( .A(n8241), .B(n8477), .Z(n8472) );
  NAND U8803 ( .A(n8242), .B(n8472), .Z(n8474) );
  AND U8804 ( .A(\stack[1][40] ), .B(o[2]), .Z(n8473) );
  XOR U8805 ( .A(n8474), .B(n8473), .Z(n8480) );
  XOR U8806 ( .A(n8481), .B(n8480), .Z(n8483) );
  XNOR U8807 ( .A(n8482), .B(n8483), .Z(n8464) );
  XOR U8808 ( .A(n8465), .B(n8464), .Z(n8467) );
  XOR U8809 ( .A(n8466), .B(n8467), .Z(n8460) );
  XOR U8810 ( .A(n8488), .B(n8487), .Z(n8490) );
  NANDN U8811 ( .A(n3000), .B(\stack[1][36] ), .Z(n8489) );
  XNOR U8812 ( .A(n8490), .B(n8489), .Z(n8496) );
  NANDN U8813 ( .A(n8244), .B(n8243), .Z(n8248) );
  NANDN U8814 ( .A(n8246), .B(n8245), .Z(n8247) );
  AND U8815 ( .A(n8248), .B(n8247), .Z(n8453) );
  XNOR U8816 ( .A(n8452), .B(n8453), .Z(n8455) );
  AND U8817 ( .A(\stack[1][34] ), .B(o[8]), .Z(n8454) );
  XNOR U8818 ( .A(n8455), .B(n8454), .Z(n8448) );
  XOR U8819 ( .A(n8449), .B(n8448), .Z(n8499) );
  XNOR U8820 ( .A(n8500), .B(n8499), .Z(n8501) );
  XNOR U8821 ( .A(n8502), .B(n8501), .Z(n8442) );
  NANDN U8822 ( .A(n2988), .B(o[11]), .Z(n8440) );
  OR U8823 ( .A(n8250), .B(n8249), .Z(n8254) );
  OR U8824 ( .A(n8252), .B(n8251), .Z(n8253) );
  NAND U8825 ( .A(n8254), .B(n8253), .Z(n8441) );
  XOR U8826 ( .A(n8440), .B(n8441), .Z(n8443) );
  XNOR U8827 ( .A(n8442), .B(n8443), .Z(n8506) );
  XNOR U8828 ( .A(n8505), .B(n8506), .Z(n8507) );
  XOR U8829 ( .A(n8436), .B(n8437), .Z(n8428) );
  OR U8830 ( .A(n8256), .B(n8255), .Z(n8260) );
  NANDN U8831 ( .A(n8258), .B(n8257), .Z(n8259) );
  AND U8832 ( .A(n8260), .B(n8259), .Z(n8429) );
  XOR U8833 ( .A(n8428), .B(n8429), .Z(n8431) );
  AND U8834 ( .A(\stack[1][28] ), .B(o[14]), .Z(n8430) );
  XOR U8835 ( .A(n8431), .B(n8430), .Z(n8513) );
  XOR U8836 ( .A(n8514), .B(n8513), .Z(n8423) );
  XOR U8837 ( .A(n8422), .B(n8423), .Z(n8424) );
  XOR U8838 ( .A(n8425), .B(n8424), .Z(n8419) );
  AND U8839 ( .A(\stack[1][25] ), .B(o[17]), .Z(n8416) );
  OR U8840 ( .A(n8262), .B(n8261), .Z(n8266) );
  OR U8841 ( .A(n8264), .B(n8263), .Z(n8265) );
  NAND U8842 ( .A(n8266), .B(n8265), .Z(n8417) );
  XNOR U8843 ( .A(n8416), .B(n8417), .Z(n8418) );
  XOR U8844 ( .A(n8419), .B(n8418), .Z(n8517) );
  XNOR U8845 ( .A(n8518), .B(n8517), .Z(n8519) );
  XNOR U8846 ( .A(n8520), .B(n8519), .Z(n8412) );
  NANDN U8847 ( .A(n2980), .B(o[19]), .Z(n8410) );
  OR U8848 ( .A(n8268), .B(n8267), .Z(n8272) );
  OR U8849 ( .A(n8270), .B(n8269), .Z(n8271) );
  NAND U8850 ( .A(n8272), .B(n8271), .Z(n8411) );
  XOR U8851 ( .A(n8410), .B(n8411), .Z(n8413) );
  XNOR U8852 ( .A(n8412), .B(n8413), .Z(n8523) );
  XNOR U8853 ( .A(n8524), .B(n8523), .Z(n8525) );
  XNOR U8854 ( .A(n8526), .B(n8525), .Z(n8406) );
  AND U8855 ( .A(\stack[1][21] ), .B(o[21]), .Z(n16672) );
  OR U8856 ( .A(n8274), .B(n8273), .Z(n8278) );
  OR U8857 ( .A(n8276), .B(n8275), .Z(n8277) );
  NAND U8858 ( .A(n8278), .B(n8277), .Z(n8405) );
  XNOR U8859 ( .A(n16672), .B(n8405), .Z(n8407) );
  XNOR U8860 ( .A(n8406), .B(n8407), .Z(n8529) );
  XNOR U8861 ( .A(n8530), .B(n8529), .Z(n8532) );
  AND U8862 ( .A(o[22]), .B(\stack[1][20] ), .Z(n8531) );
  XNOR U8863 ( .A(n8532), .B(n8531), .Z(n8401) );
  AND U8864 ( .A(o[23]), .B(\stack[1][19] ), .Z(n8399) );
  OR U8865 ( .A(n8280), .B(n8279), .Z(n8284) );
  OR U8866 ( .A(n8282), .B(n8281), .Z(n8283) );
  NAND U8867 ( .A(n8284), .B(n8283), .Z(n8400) );
  XNOR U8868 ( .A(n8399), .B(n8400), .Z(n8402) );
  XNOR U8869 ( .A(n8401), .B(n8402), .Z(n8394) );
  XNOR U8870 ( .A(n8393), .B(n8394), .Z(n8395) );
  AND U8871 ( .A(o[24]), .B(\stack[1][18] ), .Z(n8396) );
  XNOR U8872 ( .A(n8538), .B(n8537), .Z(n8388) );
  XOR U8873 ( .A(n8387), .B(n8388), .Z(n8389) );
  XOR U8874 ( .A(n8390), .B(n8389), .Z(n8384) );
  AND U8875 ( .A(o[27]), .B(\stack[1][15] ), .Z(n8381) );
  OR U8876 ( .A(n8286), .B(n8285), .Z(n8290) );
  OR U8877 ( .A(n8288), .B(n8287), .Z(n8289) );
  NAND U8878 ( .A(n8290), .B(n8289), .Z(n8382) );
  XNOR U8879 ( .A(n8381), .B(n8382), .Z(n8383) );
  XOR U8880 ( .A(n8384), .B(n8383), .Z(n8541) );
  XNOR U8881 ( .A(n8542), .B(n8541), .Z(n8543) );
  XNOR U8882 ( .A(n8544), .B(n8543), .Z(n8377) );
  NANDN U8883 ( .A(n2974), .B(o[29]), .Z(n8375) );
  OR U8884 ( .A(n8292), .B(n8291), .Z(n8296) );
  OR U8885 ( .A(n8294), .B(n8293), .Z(n8295) );
  NAND U8886 ( .A(n8296), .B(n8295), .Z(n8376) );
  XOR U8887 ( .A(n8375), .B(n8376), .Z(n8378) );
  XNOR U8888 ( .A(n8377), .B(n8378), .Z(n8547) );
  XNOR U8889 ( .A(n8548), .B(n8547), .Z(n8549) );
  XNOR U8890 ( .A(n8550), .B(n8549), .Z(n8371) );
  NANDN U8891 ( .A(n2972), .B(o[31]), .Z(n8369) );
  OR U8892 ( .A(n8298), .B(n8297), .Z(n8302) );
  OR U8893 ( .A(n8300), .B(n8299), .Z(n8301) );
  NAND U8894 ( .A(n8302), .B(n8301), .Z(n8370) );
  XOR U8895 ( .A(n8369), .B(n8370), .Z(n8372) );
  XNOR U8896 ( .A(n8371), .B(n8372), .Z(n8553) );
  XNOR U8897 ( .A(n8554), .B(n8553), .Z(n8555) );
  XNOR U8898 ( .A(n8556), .B(n8555), .Z(n8365) );
  NANDN U8899 ( .A(n17145), .B(o[33]), .Z(n8363) );
  OR U8900 ( .A(n8304), .B(n8303), .Z(n8308) );
  OR U8901 ( .A(n8306), .B(n8305), .Z(n8307) );
  NAND U8902 ( .A(n8308), .B(n8307), .Z(n8364) );
  XOR U8903 ( .A(n8363), .B(n8364), .Z(n8366) );
  XNOR U8904 ( .A(n8365), .B(n8366), .Z(n8559) );
  XNOR U8905 ( .A(n8560), .B(n8559), .Z(n8561) );
  XNOR U8906 ( .A(n8562), .B(n8561), .Z(n8359) );
  NANDN U8907 ( .A(n17219), .B(o[35]), .Z(n8357) );
  OR U8908 ( .A(n8310), .B(n8309), .Z(n8314) );
  OR U8909 ( .A(n8312), .B(n8311), .Z(n8313) );
  NAND U8910 ( .A(n8314), .B(n8313), .Z(n8358) );
  XOR U8911 ( .A(n8357), .B(n8358), .Z(n8360) );
  XNOR U8912 ( .A(n8359), .B(n8360), .Z(n8565) );
  XNOR U8913 ( .A(n8566), .B(n8565), .Z(n8567) );
  XNOR U8914 ( .A(n8568), .B(n8567), .Z(n8353) );
  NANDN U8915 ( .A(n17296), .B(o[37]), .Z(n8351) );
  OR U8916 ( .A(n8316), .B(n8315), .Z(n8320) );
  OR U8917 ( .A(n8318), .B(n8317), .Z(n8319) );
  NAND U8918 ( .A(n8320), .B(n8319), .Z(n8352) );
  XOR U8919 ( .A(n8351), .B(n8352), .Z(n8354) );
  XNOR U8920 ( .A(n8353), .B(n8354), .Z(n8571) );
  XNOR U8921 ( .A(n8572), .B(n8571), .Z(n8573) );
  XNOR U8922 ( .A(n8574), .B(n8573), .Z(n8347) );
  NANDN U8923 ( .A(n17375), .B(o[39]), .Z(n8345) );
  OR U8924 ( .A(n8322), .B(n8321), .Z(n8326) );
  OR U8925 ( .A(n8324), .B(n8323), .Z(n8325) );
  NAND U8926 ( .A(n8326), .B(n8325), .Z(n8346) );
  XOR U8927 ( .A(n8345), .B(n8346), .Z(n8348) );
  XNOR U8928 ( .A(n8347), .B(n8348), .Z(n8577) );
  XNOR U8929 ( .A(n8578), .B(n8577), .Z(n8579) );
  AND U8930 ( .A(o[41]), .B(\stack[1][1] ), .Z(n8339) );
  OR U8931 ( .A(n8328), .B(n8327), .Z(n8332) );
  OR U8932 ( .A(n8330), .B(n8329), .Z(n8331) );
  NAND U8933 ( .A(n8332), .B(n8331), .Z(n8340) );
  XNOR U8934 ( .A(n8339), .B(n8340), .Z(n8342) );
  XOR U8935 ( .A(n8341), .B(n8342), .Z(n8333) );
  NANDN U8936 ( .A(n8334), .B(n8333), .Z(n8336) );
  XOR U8937 ( .A(n8334), .B(n8333), .Z(n15860) );
  AND U8938 ( .A(o[42]), .B(\stack[1][0] ), .Z(n15861) );
  OR U8939 ( .A(n15860), .B(n15861), .Z(n8335) );
  AND U8940 ( .A(n8336), .B(n8335), .Z(n8338) );
  OR U8941 ( .A(n8337), .B(n8338), .Z(n8584) );
  XNOR U8942 ( .A(n8338), .B(n8337), .Z(n15821) );
  NANDN U8943 ( .A(n2969), .B(o[42]), .Z(n8832) );
  OR U8944 ( .A(n8340), .B(n8339), .Z(n8344) );
  OR U8945 ( .A(n8342), .B(n8341), .Z(n8343) );
  NAND U8946 ( .A(n8344), .B(n8343), .Z(n8830) );
  NANDN U8947 ( .A(n17375), .B(o[40]), .Z(n8826) );
  NANDN U8948 ( .A(n8346), .B(n8345), .Z(n8350) );
  NANDN U8949 ( .A(n8348), .B(n8347), .Z(n8349) );
  NAND U8950 ( .A(n8350), .B(n8349), .Z(n8824) );
  NANDN U8951 ( .A(n17296), .B(o[38]), .Z(n8820) );
  NANDN U8952 ( .A(n8352), .B(n8351), .Z(n8356) );
  NANDN U8953 ( .A(n8354), .B(n8353), .Z(n8355) );
  NAND U8954 ( .A(n8356), .B(n8355), .Z(n8818) );
  NANDN U8955 ( .A(n17219), .B(o[36]), .Z(n8814) );
  NANDN U8956 ( .A(n8358), .B(n8357), .Z(n8362) );
  NANDN U8957 ( .A(n8360), .B(n8359), .Z(n8361) );
  NAND U8958 ( .A(n8362), .B(n8361), .Z(n8812) );
  NANDN U8959 ( .A(n17145), .B(o[34]), .Z(n8808) );
  NANDN U8960 ( .A(n8364), .B(n8363), .Z(n8368) );
  NANDN U8961 ( .A(n8366), .B(n8365), .Z(n8367) );
  NAND U8962 ( .A(n8368), .B(n8367), .Z(n8806) );
  NANDN U8963 ( .A(n2972), .B(o[32]), .Z(n8802) );
  NANDN U8964 ( .A(n8370), .B(n8369), .Z(n8374) );
  NANDN U8965 ( .A(n8372), .B(n8371), .Z(n8373) );
  NAND U8966 ( .A(n8374), .B(n8373), .Z(n8800) );
  NANDN U8967 ( .A(n2974), .B(o[30]), .Z(n8796) );
  NANDN U8968 ( .A(n8376), .B(n8375), .Z(n8380) );
  NANDN U8969 ( .A(n8378), .B(n8377), .Z(n8379) );
  NAND U8970 ( .A(n8380), .B(n8379), .Z(n8794) );
  AND U8971 ( .A(o[28]), .B(\stack[1][15] ), .Z(n8630) );
  OR U8972 ( .A(n8382), .B(n8381), .Z(n8386) );
  OR U8973 ( .A(n8384), .B(n8383), .Z(n8385) );
  AND U8974 ( .A(n8386), .B(n8385), .Z(n8627) );
  OR U8975 ( .A(n8388), .B(n8387), .Z(n8392) );
  NANDN U8976 ( .A(n8390), .B(n8389), .Z(n8391) );
  AND U8977 ( .A(n8392), .B(n8391), .Z(n8787) );
  AND U8978 ( .A(o[27]), .B(\stack[1][16] ), .Z(n8788) );
  XNOR U8979 ( .A(n8787), .B(n8788), .Z(n8790) );
  OR U8980 ( .A(n8394), .B(n8393), .Z(n8398) );
  OR U8981 ( .A(n8396), .B(n8395), .Z(n8397) );
  NAND U8982 ( .A(n8398), .B(n8397), .Z(n8640) );
  ANDN U8983 ( .B(\stack[1][18] ), .A(n3019), .Z(n8639) );
  XOR U8984 ( .A(n8640), .B(n8639), .Z(n8641) );
  NANDN U8985 ( .A(n16746), .B(o[24]), .Z(n8784) );
  OR U8986 ( .A(n8400), .B(n8399), .Z(n8404) );
  OR U8987 ( .A(n8402), .B(n8401), .Z(n8403) );
  NAND U8988 ( .A(n8404), .B(n8403), .Z(n8782) );
  NANDN U8989 ( .A(n2978), .B(o[22]), .Z(n8778) );
  OR U8990 ( .A(n8405), .B(n16672), .Z(n8409) );
  NANDN U8991 ( .A(n8407), .B(n8406), .Z(n8408) );
  NAND U8992 ( .A(n8409), .B(n8408), .Z(n8776) );
  NANDN U8993 ( .A(n3014), .B(\stack[1][23] ), .Z(n8772) );
  NANDN U8994 ( .A(n8411), .B(n8410), .Z(n8415) );
  NANDN U8995 ( .A(n8413), .B(n8412), .Z(n8414) );
  NAND U8996 ( .A(n8415), .B(n8414), .Z(n8770) );
  AND U8997 ( .A(\stack[1][25] ), .B(o[18]), .Z(n8666) );
  OR U8998 ( .A(n8417), .B(n8416), .Z(n8421) );
  OR U8999 ( .A(n8419), .B(n8418), .Z(n8420) );
  AND U9000 ( .A(n8421), .B(n8420), .Z(n8663) );
  OR U9001 ( .A(n8423), .B(n8422), .Z(n8427) );
  NANDN U9002 ( .A(n8425), .B(n8424), .Z(n8426) );
  AND U9003 ( .A(n8427), .B(n8426), .Z(n8763) );
  AND U9004 ( .A(\stack[1][26] ), .B(o[17]), .Z(n8764) );
  XNOR U9005 ( .A(n8763), .B(n8764), .Z(n8766) );
  NANDN U9006 ( .A(n8429), .B(n8428), .Z(n8433) );
  OR U9007 ( .A(n8431), .B(n8430), .Z(n8432) );
  NAND U9008 ( .A(n8433), .B(n8432), .Z(n8676) );
  ANDN U9009 ( .B(o[15]), .A(n2985), .Z(n8675) );
  XNOR U9010 ( .A(n8676), .B(n8675), .Z(n8677) );
  NANDN U9011 ( .A(n3008), .B(\stack[1][29] ), .Z(n8760) );
  NANDN U9012 ( .A(n8435), .B(n8434), .Z(n8439) );
  NANDN U9013 ( .A(n8437), .B(n8436), .Z(n8438) );
  AND U9014 ( .A(n8439), .B(n8438), .Z(n8757) );
  NANDN U9015 ( .A(n3006), .B(\stack[1][31] ), .Z(n8690) );
  NANDN U9016 ( .A(n8441), .B(n8440), .Z(n8445) );
  NANDN U9017 ( .A(n8443), .B(n8442), .Z(n8444) );
  NAND U9018 ( .A(n8445), .B(n8444), .Z(n8688) );
  NANDN U9019 ( .A(n3004), .B(\stack[1][33] ), .Z(n8696) );
  OR U9020 ( .A(n8447), .B(n8446), .Z(n8451) );
  OR U9021 ( .A(n8449), .B(n8448), .Z(n8450) );
  NAND U9022 ( .A(n8451), .B(n8450), .Z(n8694) );
  OR U9023 ( .A(n8453), .B(n8452), .Z(n8457) );
  OR U9024 ( .A(n8455), .B(n8454), .Z(n8456) );
  AND U9025 ( .A(n8457), .B(n8456), .Z(n8699) );
  AND U9026 ( .A(\stack[1][34] ), .B(o[9]), .Z(n8700) );
  XNOR U9027 ( .A(n8699), .B(n8700), .Z(n8702) );
  OR U9028 ( .A(n8459), .B(n8458), .Z(n8463) );
  OR U9029 ( .A(n8461), .B(n8460), .Z(n8462) );
  NAND U9030 ( .A(n8463), .B(n8462), .Z(n8712) );
  ANDN U9031 ( .B(\stack[1][38] ), .A(n2999), .Z(n8720) );
  NANDN U9032 ( .A(n8465), .B(n8464), .Z(n8469) );
  NANDN U9033 ( .A(n8467), .B(n8466), .Z(n8468) );
  AND U9034 ( .A(n8469), .B(n8468), .Z(n8717) );
  AND U9035 ( .A(\stack[1][39] ), .B(o[4]), .Z(n8726) );
  AND U9036 ( .A(\stack[1][40] ), .B(o[3]), .Z(n8742) );
  NANDN U9037 ( .A(n8470), .B(n8729), .Z(n8471) );
  AND U9038 ( .A(n8472), .B(n8471), .Z(n8476) );
  OR U9039 ( .A(n8474), .B(n8473), .Z(n8475) );
  AND U9040 ( .A(n8476), .B(n8475), .Z(n8739) );
  AND U9041 ( .A(\stack[1][43] ), .B(o[1]), .Z(n8737) );
  ANDN U9042 ( .B(n8737), .A(n8477), .Z(n8979) );
  XNOR U9043 ( .A(n8979), .B(n8729), .Z(n8479) );
  NAND U9044 ( .A(\stack[1][43] ), .B(o[0]), .Z(n8736) );
  NANDN U9045 ( .A(n8478), .B(n8736), .Z(n8731) );
  NAND U9046 ( .A(n8479), .B(n8731), .Z(n8733) );
  AND U9047 ( .A(\stack[1][41] ), .B(o[2]), .Z(n8732) );
  XNOR U9048 ( .A(n8733), .B(n8732), .Z(n8740) );
  XOR U9049 ( .A(n8739), .B(n8740), .Z(n8741) );
  XOR U9050 ( .A(n8742), .B(n8741), .Z(n8724) );
  NANDN U9051 ( .A(n8481), .B(n8480), .Z(n8485) );
  NANDN U9052 ( .A(n8483), .B(n8482), .Z(n8484) );
  AND U9053 ( .A(n8485), .B(n8484), .Z(n8723) );
  XOR U9054 ( .A(n8724), .B(n8723), .Z(n8725) );
  XOR U9055 ( .A(n8726), .B(n8725), .Z(n8718) );
  XNOR U9056 ( .A(n8717), .B(n8718), .Z(n8719) );
  IV U9057 ( .A(n8719), .Z(n8486) );
  XOR U9058 ( .A(n8720), .B(n8486), .Z(n8711) );
  XOR U9059 ( .A(n8712), .B(n8711), .Z(n8714) );
  AND U9060 ( .A(\stack[1][37] ), .B(o[6]), .Z(n8713) );
  XNOR U9061 ( .A(n8714), .B(n8713), .Z(n8707) );
  AND U9062 ( .A(\stack[1][36] ), .B(o[7]), .Z(n8705) );
  NANDN U9063 ( .A(n8488), .B(n8487), .Z(n8492) );
  OR U9064 ( .A(n8490), .B(n8489), .Z(n8491) );
  NAND U9065 ( .A(n8492), .B(n8491), .Z(n8706) );
  XNOR U9066 ( .A(n8705), .B(n8706), .Z(n8708) );
  XNOR U9067 ( .A(n8707), .B(n8708), .Z(n8746) );
  OR U9068 ( .A(n8494), .B(n8493), .Z(n8498) );
  OR U9069 ( .A(n8496), .B(n8495), .Z(n8497) );
  NAND U9070 ( .A(n8498), .B(n8497), .Z(n8745) );
  XOR U9071 ( .A(n8746), .B(n8745), .Z(n8747) );
  AND U9072 ( .A(\stack[1][35] ), .B(o[8]), .Z(n8748) );
  XOR U9073 ( .A(n8747), .B(n8748), .Z(n8701) );
  XOR U9074 ( .A(n8702), .B(n8701), .Z(n8693) );
  XNOR U9075 ( .A(n8694), .B(n8693), .Z(n8695) );
  XNOR U9076 ( .A(n8696), .B(n8695), .Z(n8753) );
  NANDN U9077 ( .A(n2989), .B(o[11]), .Z(n8751) );
  OR U9078 ( .A(n8500), .B(n8499), .Z(n8504) );
  OR U9079 ( .A(n8502), .B(n8501), .Z(n8503) );
  NAND U9080 ( .A(n8504), .B(n8503), .Z(n8752) );
  XOR U9081 ( .A(n8751), .B(n8752), .Z(n8754) );
  XNOR U9082 ( .A(n8753), .B(n8754), .Z(n8687) );
  XNOR U9083 ( .A(n8688), .B(n8687), .Z(n8689) );
  XNOR U9084 ( .A(n8690), .B(n8689), .Z(n8683) );
  NANDN U9085 ( .A(n2987), .B(o[13]), .Z(n8681) );
  OR U9086 ( .A(n8506), .B(n8505), .Z(n8510) );
  OR U9087 ( .A(n8508), .B(n8507), .Z(n8509) );
  NAND U9088 ( .A(n8510), .B(n8509), .Z(n8682) );
  XOR U9089 ( .A(n8681), .B(n8682), .Z(n8684) );
  XNOR U9090 ( .A(n8683), .B(n8684), .Z(n8758) );
  XNOR U9091 ( .A(n8757), .B(n8758), .Z(n8759) );
  XOR U9092 ( .A(n8677), .B(n8678), .Z(n8669) );
  OR U9093 ( .A(n8512), .B(n8511), .Z(n8516) );
  NANDN U9094 ( .A(n8514), .B(n8513), .Z(n8515) );
  AND U9095 ( .A(n8516), .B(n8515), .Z(n8670) );
  XOR U9096 ( .A(n8669), .B(n8670), .Z(n8672) );
  AND U9097 ( .A(\stack[1][27] ), .B(o[16]), .Z(n8671) );
  XOR U9098 ( .A(n8672), .B(n8671), .Z(n8765) );
  XOR U9099 ( .A(n8766), .B(n8765), .Z(n8664) );
  XOR U9100 ( .A(n8663), .B(n8664), .Z(n8665) );
  XOR U9101 ( .A(n8666), .B(n8665), .Z(n8660) );
  AND U9102 ( .A(\stack[1][24] ), .B(o[19]), .Z(n8657) );
  OR U9103 ( .A(n8518), .B(n8517), .Z(n8522) );
  OR U9104 ( .A(n8520), .B(n8519), .Z(n8521) );
  NAND U9105 ( .A(n8522), .B(n8521), .Z(n8658) );
  XNOR U9106 ( .A(n8657), .B(n8658), .Z(n8659) );
  XOR U9107 ( .A(n8660), .B(n8659), .Z(n8769) );
  XNOR U9108 ( .A(n8770), .B(n8769), .Z(n8771) );
  XNOR U9109 ( .A(n8772), .B(n8771), .Z(n8653) );
  NANDN U9110 ( .A(n2979), .B(o[21]), .Z(n8651) );
  OR U9111 ( .A(n8524), .B(n8523), .Z(n8528) );
  OR U9112 ( .A(n8526), .B(n8525), .Z(n8527) );
  NAND U9113 ( .A(n8528), .B(n8527), .Z(n8652) );
  XOR U9114 ( .A(n8651), .B(n8652), .Z(n8654) );
  XNOR U9115 ( .A(n8653), .B(n8654), .Z(n8775) );
  XNOR U9116 ( .A(n8776), .B(n8775), .Z(n8777) );
  XNOR U9117 ( .A(n8778), .B(n8777), .Z(n8647) );
  AND U9118 ( .A(o[23]), .B(\stack[1][20] ), .Z(n8645) );
  OR U9119 ( .A(n8530), .B(n8529), .Z(n8534) );
  NANDN U9120 ( .A(n8532), .B(n8531), .Z(n8533) );
  NAND U9121 ( .A(n8534), .B(n8533), .Z(n8646) );
  XNOR U9122 ( .A(n8645), .B(n8646), .Z(n8648) );
  XNOR U9123 ( .A(n8647), .B(n8648), .Z(n8781) );
  XNOR U9124 ( .A(n8782), .B(n8781), .Z(n8783) );
  XNOR U9125 ( .A(n8784), .B(n8783), .Z(n8642) );
  OR U9126 ( .A(n8536), .B(n8535), .Z(n8540) );
  OR U9127 ( .A(n8538), .B(n8537), .Z(n8539) );
  AND U9128 ( .A(n8540), .B(n8539), .Z(n8634) );
  XNOR U9129 ( .A(n8633), .B(n8634), .Z(n8636) );
  AND U9130 ( .A(o[26]), .B(\stack[1][17] ), .Z(n8635) );
  XOR U9131 ( .A(n8636), .B(n8635), .Z(n8789) );
  XOR U9132 ( .A(n8790), .B(n8789), .Z(n8628) );
  XOR U9133 ( .A(n8627), .B(n8628), .Z(n8629) );
  XOR U9134 ( .A(n8630), .B(n8629), .Z(n8624) );
  AND U9135 ( .A(o[29]), .B(\stack[1][14] ), .Z(n8621) );
  OR U9136 ( .A(n8542), .B(n8541), .Z(n8546) );
  OR U9137 ( .A(n8544), .B(n8543), .Z(n8545) );
  NAND U9138 ( .A(n8546), .B(n8545), .Z(n8622) );
  XNOR U9139 ( .A(n8621), .B(n8622), .Z(n8623) );
  XOR U9140 ( .A(n8624), .B(n8623), .Z(n8793) );
  XNOR U9141 ( .A(n8794), .B(n8793), .Z(n8795) );
  XNOR U9142 ( .A(n8796), .B(n8795), .Z(n8617) );
  NANDN U9143 ( .A(n2973), .B(o[31]), .Z(n8615) );
  OR U9144 ( .A(n8548), .B(n8547), .Z(n8552) );
  OR U9145 ( .A(n8550), .B(n8549), .Z(n8551) );
  NAND U9146 ( .A(n8552), .B(n8551), .Z(n8616) );
  XOR U9147 ( .A(n8615), .B(n8616), .Z(n8618) );
  XNOR U9148 ( .A(n8617), .B(n8618), .Z(n8799) );
  XNOR U9149 ( .A(n8800), .B(n8799), .Z(n8801) );
  XNOR U9150 ( .A(n8802), .B(n8801), .Z(n8611) );
  NANDN U9151 ( .A(n17101), .B(o[33]), .Z(n8609) );
  OR U9152 ( .A(n8554), .B(n8553), .Z(n8558) );
  OR U9153 ( .A(n8556), .B(n8555), .Z(n8557) );
  NAND U9154 ( .A(n8558), .B(n8557), .Z(n8610) );
  XOR U9155 ( .A(n8609), .B(n8610), .Z(n8612) );
  XNOR U9156 ( .A(n8611), .B(n8612), .Z(n8805) );
  XNOR U9157 ( .A(n8806), .B(n8805), .Z(n8807) );
  XNOR U9158 ( .A(n8808), .B(n8807), .Z(n8605) );
  NANDN U9159 ( .A(n17179), .B(o[35]), .Z(n8603) );
  OR U9160 ( .A(n8560), .B(n8559), .Z(n8564) );
  OR U9161 ( .A(n8562), .B(n8561), .Z(n8563) );
  NAND U9162 ( .A(n8564), .B(n8563), .Z(n8604) );
  XOR U9163 ( .A(n8603), .B(n8604), .Z(n8606) );
  XNOR U9164 ( .A(n8605), .B(n8606), .Z(n8811) );
  XNOR U9165 ( .A(n8812), .B(n8811), .Z(n8813) );
  XNOR U9166 ( .A(n8814), .B(n8813), .Z(n8599) );
  NANDN U9167 ( .A(n17256), .B(o[37]), .Z(n8597) );
  OR U9168 ( .A(n8566), .B(n8565), .Z(n8570) );
  OR U9169 ( .A(n8568), .B(n8567), .Z(n8569) );
  NAND U9170 ( .A(n8570), .B(n8569), .Z(n8598) );
  XOR U9171 ( .A(n8597), .B(n8598), .Z(n8600) );
  XNOR U9172 ( .A(n8599), .B(n8600), .Z(n8817) );
  XNOR U9173 ( .A(n8818), .B(n8817), .Z(n8819) );
  XNOR U9174 ( .A(n8820), .B(n8819), .Z(n8593) );
  AND U9175 ( .A(o[39]), .B(\stack[1][4] ), .Z(n8591) );
  OR U9176 ( .A(n8572), .B(n8571), .Z(n8576) );
  OR U9177 ( .A(n8574), .B(n8573), .Z(n8575) );
  NAND U9178 ( .A(n8576), .B(n8575), .Z(n8592) );
  XNOR U9179 ( .A(n8591), .B(n8592), .Z(n8594) );
  XNOR U9180 ( .A(n8593), .B(n8594), .Z(n8823) );
  XNOR U9181 ( .A(n8824), .B(n8823), .Z(n8825) );
  XOR U9182 ( .A(n8826), .B(n8825), .Z(n8588) );
  AND U9183 ( .A(o[41]), .B(\stack[1][2] ), .Z(n8585) );
  OR U9184 ( .A(n8578), .B(n8577), .Z(n8582) );
  OR U9185 ( .A(n8580), .B(n8579), .Z(n8581) );
  NAND U9186 ( .A(n8582), .B(n8581), .Z(n8586) );
  XOR U9187 ( .A(n8585), .B(n8586), .Z(n8587) );
  XNOR U9188 ( .A(n8588), .B(n8587), .Z(n8829) );
  XNOR U9189 ( .A(n8830), .B(n8829), .Z(n8831) );
  XOR U9190 ( .A(n8832), .B(n8831), .Z(n15822) );
  OR U9191 ( .A(n15821), .B(n15822), .Z(n8583) );
  AND U9192 ( .A(n8584), .B(n8583), .Z(n8836) );
  NANDN U9193 ( .A(n2970), .B(o[42]), .Z(n9094) );
  OR U9194 ( .A(n8586), .B(n8585), .Z(n8590) );
  NANDN U9195 ( .A(n8588), .B(n8587), .Z(n8589) );
  NAND U9196 ( .A(n8590), .B(n8589), .Z(n9092) );
  NANDN U9197 ( .A(n2971), .B(o[40]), .Z(n9088) );
  OR U9198 ( .A(n8592), .B(n8591), .Z(n8596) );
  NANDN U9199 ( .A(n8594), .B(n8593), .Z(n8595) );
  NAND U9200 ( .A(n8596), .B(n8595), .Z(n9086) );
  NANDN U9201 ( .A(n17256), .B(o[38]), .Z(n9082) );
  NANDN U9202 ( .A(n8598), .B(n8597), .Z(n8602) );
  NANDN U9203 ( .A(n8600), .B(n8599), .Z(n8601) );
  NAND U9204 ( .A(n8602), .B(n8601), .Z(n9080) );
  NANDN U9205 ( .A(n17179), .B(o[36]), .Z(n9076) );
  NANDN U9206 ( .A(n8604), .B(n8603), .Z(n8608) );
  NANDN U9207 ( .A(n8606), .B(n8605), .Z(n8607) );
  NAND U9208 ( .A(n8608), .B(n8607), .Z(n9074) );
  NANDN U9209 ( .A(n17101), .B(o[34]), .Z(n9070) );
  NANDN U9210 ( .A(n8610), .B(n8609), .Z(n8614) );
  NANDN U9211 ( .A(n8612), .B(n8611), .Z(n8613) );
  NAND U9212 ( .A(n8614), .B(n8613), .Z(n9068) );
  NANDN U9213 ( .A(n2973), .B(o[32]), .Z(n9064) );
  NANDN U9214 ( .A(n8616), .B(n8615), .Z(n8620) );
  NANDN U9215 ( .A(n8618), .B(n8617), .Z(n8619) );
  NAND U9216 ( .A(n8620), .B(n8619), .Z(n9062) );
  AND U9217 ( .A(o[30]), .B(\stack[1][14] ), .Z(n8886) );
  OR U9218 ( .A(n8622), .B(n8621), .Z(n8626) );
  OR U9219 ( .A(n8624), .B(n8623), .Z(n8625) );
  AND U9220 ( .A(n8626), .B(n8625), .Z(n8883) );
  OR U9221 ( .A(n8628), .B(n8627), .Z(n8632) );
  NANDN U9222 ( .A(n8630), .B(n8629), .Z(n8631) );
  AND U9223 ( .A(n8632), .B(n8631), .Z(n9055) );
  AND U9224 ( .A(o[29]), .B(\stack[1][15] ), .Z(n9056) );
  XNOR U9225 ( .A(n9055), .B(n9056), .Z(n9058) );
  OR U9226 ( .A(n8634), .B(n8633), .Z(n8638) );
  OR U9227 ( .A(n8636), .B(n8635), .Z(n8637) );
  NAND U9228 ( .A(n8638), .B(n8637), .Z(n8896) );
  ANDN U9229 ( .B(o[27]), .A(n16826), .Z(n8895) );
  XNOR U9230 ( .A(n8896), .B(n8895), .Z(n8897) );
  NANDN U9231 ( .A(n16786), .B(o[26]), .Z(n9052) );
  NANDN U9232 ( .A(n8640), .B(n8639), .Z(n8644) );
  OR U9233 ( .A(n8642), .B(n8641), .Z(n8643) );
  AND U9234 ( .A(n8644), .B(n8643), .Z(n9049) );
  NANDN U9235 ( .A(n16712), .B(o[24]), .Z(n9046) );
  OR U9236 ( .A(n8646), .B(n8645), .Z(n8650) );
  NANDN U9237 ( .A(n8648), .B(n8647), .Z(n8649) );
  NAND U9238 ( .A(n8650), .B(n8649), .Z(n9044) );
  NOR U9239 ( .A(n3016), .B(n2979), .Z(n9039) );
  NANDN U9240 ( .A(n8652), .B(n8651), .Z(n8656) );
  NANDN U9241 ( .A(n8654), .B(n8653), .Z(n8655) );
  NAND U9242 ( .A(n8656), .B(n8655), .Z(n9038) );
  AND U9243 ( .A(\stack[1][24] ), .B(o[20]), .Z(n8922) );
  OR U9244 ( .A(n8658), .B(n8657), .Z(n8662) );
  OR U9245 ( .A(n8660), .B(n8659), .Z(n8661) );
  AND U9246 ( .A(n8662), .B(n8661), .Z(n8919) );
  OR U9247 ( .A(n8664), .B(n8663), .Z(n8668) );
  NANDN U9248 ( .A(n8666), .B(n8665), .Z(n8667) );
  AND U9249 ( .A(n8668), .B(n8667), .Z(n9031) );
  AND U9250 ( .A(\stack[1][25] ), .B(o[19]), .Z(n9032) );
  XNOR U9251 ( .A(n9031), .B(n9032), .Z(n9034) );
  NANDN U9252 ( .A(n8670), .B(n8669), .Z(n8674) );
  OR U9253 ( .A(n8672), .B(n8671), .Z(n8673) );
  NAND U9254 ( .A(n8674), .B(n8673), .Z(n8932) );
  ANDN U9255 ( .B(o[17]), .A(n2984), .Z(n8931) );
  XNOR U9256 ( .A(n8932), .B(n8931), .Z(n8933) );
  NANDN U9257 ( .A(n3010), .B(\stack[1][28] ), .Z(n8940) );
  NANDN U9258 ( .A(n8676), .B(n8675), .Z(n8680) );
  NANDN U9259 ( .A(n8678), .B(n8677), .Z(n8679) );
  AND U9260 ( .A(n8680), .B(n8679), .Z(n8937) );
  NANDN U9261 ( .A(n3008), .B(\stack[1][30] ), .Z(n8946) );
  NANDN U9262 ( .A(n8682), .B(n8681), .Z(n8686) );
  NANDN U9263 ( .A(n8684), .B(n8683), .Z(n8685) );
  NAND U9264 ( .A(n8686), .B(n8685), .Z(n8944) );
  AND U9265 ( .A(\stack[1][31] ), .B(o[13]), .Z(n8949) );
  OR U9266 ( .A(n8688), .B(n8687), .Z(n8692) );
  OR U9267 ( .A(n8690), .B(n8689), .Z(n8691) );
  NAND U9268 ( .A(n8692), .B(n8691), .Z(n8950) );
  XNOR U9269 ( .A(n8949), .B(n8950), .Z(n8952) );
  NANDN U9270 ( .A(n3005), .B(\stack[1][33] ), .Z(n9020) );
  OR U9271 ( .A(n8694), .B(n8693), .Z(n8698) );
  OR U9272 ( .A(n8696), .B(n8695), .Z(n8697) );
  AND U9273 ( .A(n8698), .B(n8697), .Z(n9019) );
  XNOR U9274 ( .A(n9020), .B(n9019), .Z(n9021) );
  OR U9275 ( .A(n8700), .B(n8699), .Z(n8704) );
  OR U9276 ( .A(n8702), .B(n8701), .Z(n8703) );
  NAND U9277 ( .A(n8704), .B(n8703), .Z(n9014) );
  AND U9278 ( .A(\stack[1][36] ), .B(o[8]), .Z(n9010) );
  OR U9279 ( .A(n8706), .B(n8705), .Z(n8710) );
  OR U9280 ( .A(n8708), .B(n8707), .Z(n8709) );
  AND U9281 ( .A(n8710), .B(n8709), .Z(n9007) );
  AND U9282 ( .A(\stack[1][37] ), .B(o[7]), .Z(n9001) );
  NANDN U9283 ( .A(n8712), .B(n8711), .Z(n8716) );
  NANDN U9284 ( .A(n8714), .B(n8713), .Z(n8715) );
  NAND U9285 ( .A(n8716), .B(n8715), .Z(n9002) );
  XNOR U9286 ( .A(n9001), .B(n9002), .Z(n9004) );
  NANDN U9287 ( .A(n3000), .B(\stack[1][38] ), .Z(n8969) );
  OR U9288 ( .A(n8718), .B(n8717), .Z(n8722) );
  OR U9289 ( .A(n8720), .B(n8719), .Z(n8721) );
  AND U9290 ( .A(n8722), .B(n8721), .Z(n8968) );
  NANDN U9291 ( .A(n2999), .B(\stack[1][39] ), .Z(n8997) );
  OR U9292 ( .A(n8724), .B(n8723), .Z(n8728) );
  NANDN U9293 ( .A(n8726), .B(n8725), .Z(n8727) );
  AND U9294 ( .A(n8728), .B(n8727), .Z(n8996) );
  IV U9295 ( .A(\stack[1][40] ), .Z(n15935) );
  NANDN U9296 ( .A(n15935), .B(o[4]), .Z(n8975) );
  AND U9297 ( .A(\stack[1][41] ), .B(o[3]), .Z(n8992) );
  NANDN U9298 ( .A(n8729), .B(n8979), .Z(n8730) );
  AND U9299 ( .A(n8731), .B(n8730), .Z(n8735) );
  OR U9300 ( .A(n8733), .B(n8732), .Z(n8734) );
  AND U9301 ( .A(n8735), .B(n8734), .Z(n8989) );
  AND U9302 ( .A(\stack[1][44] ), .B(o[1]), .Z(n8987) );
  ANDN U9303 ( .B(n8987), .A(n8736), .Z(n9243) );
  XNOR U9304 ( .A(n9243), .B(n8979), .Z(n8738) );
  NAND U9305 ( .A(\stack[1][44] ), .B(o[0]), .Z(n8986) );
  NANDN U9306 ( .A(n8737), .B(n8986), .Z(n8981) );
  NAND U9307 ( .A(n8738), .B(n8981), .Z(n8983) );
  AND U9308 ( .A(\stack[1][42] ), .B(o[2]), .Z(n8982) );
  XNOR U9309 ( .A(n8983), .B(n8982), .Z(n8990) );
  XOR U9310 ( .A(n8989), .B(n8990), .Z(n8991) );
  XOR U9311 ( .A(n8992), .B(n8991), .Z(n8974) );
  OR U9312 ( .A(n8740), .B(n8739), .Z(n8744) );
  NANDN U9313 ( .A(n8742), .B(n8741), .Z(n8743) );
  AND U9314 ( .A(n8744), .B(n8743), .Z(n8973) );
  XNOR U9315 ( .A(n8974), .B(n8973), .Z(n8976) );
  XNOR U9316 ( .A(n8975), .B(n8976), .Z(n8995) );
  XOR U9317 ( .A(n8996), .B(n8995), .Z(n8998) );
  XNOR U9318 ( .A(n8997), .B(n8998), .Z(n8967) );
  XOR U9319 ( .A(n8968), .B(n8967), .Z(n8970) );
  XNOR U9320 ( .A(n8969), .B(n8970), .Z(n9003) );
  XOR U9321 ( .A(n9004), .B(n9003), .Z(n9008) );
  XOR U9322 ( .A(n9007), .B(n9008), .Z(n9009) );
  XOR U9323 ( .A(n9010), .B(n9009), .Z(n8964) );
  OR U9324 ( .A(n8746), .B(n8745), .Z(n8750) );
  NANDN U9325 ( .A(n8748), .B(n8747), .Z(n8749) );
  AND U9326 ( .A(n8750), .B(n8749), .Z(n8962) );
  NANDN U9327 ( .A(n2992), .B(o[9]), .Z(n8961) );
  XOR U9328 ( .A(n8962), .B(n8961), .Z(n8963) );
  XNOR U9329 ( .A(n8964), .B(n8963), .Z(n9013) );
  XOR U9330 ( .A(n9014), .B(n9013), .Z(n9016) );
  NANDN U9331 ( .A(n3004), .B(\stack[1][34] ), .Z(n9015) );
  XNOR U9332 ( .A(n9016), .B(n9015), .Z(n9022) );
  NANDN U9333 ( .A(n8752), .B(n8751), .Z(n8756) );
  NANDN U9334 ( .A(n8754), .B(n8753), .Z(n8755) );
  AND U9335 ( .A(n8756), .B(n8755), .Z(n8956) );
  XNOR U9336 ( .A(n8955), .B(n8956), .Z(n8958) );
  AND U9337 ( .A(\stack[1][32] ), .B(o[12]), .Z(n8957) );
  XNOR U9338 ( .A(n8958), .B(n8957), .Z(n8951) );
  XOR U9339 ( .A(n8952), .B(n8951), .Z(n8943) );
  XNOR U9340 ( .A(n8944), .B(n8943), .Z(n8945) );
  XNOR U9341 ( .A(n8946), .B(n8945), .Z(n9027) );
  NANDN U9342 ( .A(n2986), .B(o[15]), .Z(n9025) );
  OR U9343 ( .A(n8758), .B(n8757), .Z(n8762) );
  OR U9344 ( .A(n8760), .B(n8759), .Z(n8761) );
  NAND U9345 ( .A(n8762), .B(n8761), .Z(n9026) );
  XOR U9346 ( .A(n9025), .B(n9026), .Z(n9028) );
  XNOR U9347 ( .A(n9027), .B(n9028), .Z(n8938) );
  XNOR U9348 ( .A(n8937), .B(n8938), .Z(n8939) );
  XOR U9349 ( .A(n8933), .B(n8934), .Z(n8925) );
  OR U9350 ( .A(n8764), .B(n8763), .Z(n8768) );
  NANDN U9351 ( .A(n8766), .B(n8765), .Z(n8767) );
  AND U9352 ( .A(n8768), .B(n8767), .Z(n8926) );
  XOR U9353 ( .A(n8925), .B(n8926), .Z(n8928) );
  AND U9354 ( .A(\stack[1][26] ), .B(o[18]), .Z(n8927) );
  XOR U9355 ( .A(n8928), .B(n8927), .Z(n9033) );
  XOR U9356 ( .A(n9034), .B(n9033), .Z(n8920) );
  XOR U9357 ( .A(n8919), .B(n8920), .Z(n8921) );
  XOR U9358 ( .A(n8922), .B(n8921), .Z(n8916) );
  AND U9359 ( .A(\stack[1][23] ), .B(o[21]), .Z(n8913) );
  OR U9360 ( .A(n8770), .B(n8769), .Z(n8774) );
  OR U9361 ( .A(n8772), .B(n8771), .Z(n8773) );
  NAND U9362 ( .A(n8774), .B(n8773), .Z(n8914) );
  XNOR U9363 ( .A(n8913), .B(n8914), .Z(n8915) );
  XOR U9364 ( .A(n8916), .B(n8915), .Z(n9037) );
  XNOR U9365 ( .A(n9038), .B(n9037), .Z(n9040) );
  XOR U9366 ( .A(n9039), .B(n9040), .Z(n8909) );
  NANDN U9367 ( .A(n3017), .B(\stack[1][21] ), .Z(n8907) );
  OR U9368 ( .A(n8776), .B(n8775), .Z(n8780) );
  OR U9369 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U9370 ( .A(n8780), .B(n8779), .Z(n8908) );
  XOR U9371 ( .A(n8907), .B(n8908), .Z(n8910) );
  XNOR U9372 ( .A(n8909), .B(n8910), .Z(n9043) );
  XNOR U9373 ( .A(n9044), .B(n9043), .Z(n9045) );
  XNOR U9374 ( .A(n9046), .B(n9045), .Z(n8903) );
  NANDN U9375 ( .A(n3019), .B(\stack[1][19] ), .Z(n8901) );
  OR U9376 ( .A(n8782), .B(n8781), .Z(n8786) );
  OR U9377 ( .A(n8784), .B(n8783), .Z(n8785) );
  NAND U9378 ( .A(n8786), .B(n8785), .Z(n8902) );
  XOR U9379 ( .A(n8901), .B(n8902), .Z(n8904) );
  XNOR U9380 ( .A(n8903), .B(n8904), .Z(n9050) );
  XNOR U9381 ( .A(n9049), .B(n9050), .Z(n9051) );
  XOR U9382 ( .A(n8897), .B(n8898), .Z(n8889) );
  OR U9383 ( .A(n8788), .B(n8787), .Z(n8792) );
  NANDN U9384 ( .A(n8790), .B(n8789), .Z(n8791) );
  AND U9385 ( .A(n8792), .B(n8791), .Z(n8890) );
  XOR U9386 ( .A(n8889), .B(n8890), .Z(n8892) );
  AND U9387 ( .A(o[28]), .B(\stack[1][16] ), .Z(n8891) );
  XOR U9388 ( .A(n8892), .B(n8891), .Z(n9057) );
  XOR U9389 ( .A(n9058), .B(n9057), .Z(n8884) );
  XOR U9390 ( .A(n8883), .B(n8884), .Z(n8885) );
  XOR U9391 ( .A(n8886), .B(n8885), .Z(n8880) );
  AND U9392 ( .A(o[31]), .B(\stack[1][13] ), .Z(n8877) );
  OR U9393 ( .A(n8794), .B(n8793), .Z(n8798) );
  OR U9394 ( .A(n8796), .B(n8795), .Z(n8797) );
  NAND U9395 ( .A(n8798), .B(n8797), .Z(n8878) );
  XNOR U9396 ( .A(n8877), .B(n8878), .Z(n8879) );
  XOR U9397 ( .A(n8880), .B(n8879), .Z(n9061) );
  XNOR U9398 ( .A(n9062), .B(n9061), .Z(n9063) );
  XNOR U9399 ( .A(n9064), .B(n9063), .Z(n8873) );
  NANDN U9400 ( .A(n2972), .B(o[33]), .Z(n8871) );
  OR U9401 ( .A(n8800), .B(n8799), .Z(n8804) );
  OR U9402 ( .A(n8802), .B(n8801), .Z(n8803) );
  NAND U9403 ( .A(n8804), .B(n8803), .Z(n8872) );
  XOR U9404 ( .A(n8871), .B(n8872), .Z(n8874) );
  XNOR U9405 ( .A(n8873), .B(n8874), .Z(n9067) );
  XNOR U9406 ( .A(n9068), .B(n9067), .Z(n9069) );
  XNOR U9407 ( .A(n9070), .B(n9069), .Z(n8867) );
  NANDN U9408 ( .A(n17145), .B(o[35]), .Z(n8865) );
  OR U9409 ( .A(n8806), .B(n8805), .Z(n8810) );
  OR U9410 ( .A(n8808), .B(n8807), .Z(n8809) );
  NAND U9411 ( .A(n8810), .B(n8809), .Z(n8866) );
  XOR U9412 ( .A(n8865), .B(n8866), .Z(n8868) );
  XNOR U9413 ( .A(n8867), .B(n8868), .Z(n9073) );
  XNOR U9414 ( .A(n9074), .B(n9073), .Z(n9075) );
  XNOR U9415 ( .A(n9076), .B(n9075), .Z(n8861) );
  NANDN U9416 ( .A(n17219), .B(o[37]), .Z(n8859) );
  OR U9417 ( .A(n8812), .B(n8811), .Z(n8816) );
  OR U9418 ( .A(n8814), .B(n8813), .Z(n8815) );
  NAND U9419 ( .A(n8816), .B(n8815), .Z(n8860) );
  XOR U9420 ( .A(n8859), .B(n8860), .Z(n8862) );
  XNOR U9421 ( .A(n8861), .B(n8862), .Z(n9079) );
  XNOR U9422 ( .A(n9080), .B(n9079), .Z(n9081) );
  XNOR U9423 ( .A(n9082), .B(n9081), .Z(n8855) );
  NANDN U9424 ( .A(n17296), .B(o[39]), .Z(n8853) );
  OR U9425 ( .A(n8818), .B(n8817), .Z(n8822) );
  OR U9426 ( .A(n8820), .B(n8819), .Z(n8821) );
  NAND U9427 ( .A(n8822), .B(n8821), .Z(n8854) );
  XOR U9428 ( .A(n8853), .B(n8854), .Z(n8856) );
  XNOR U9429 ( .A(n8855), .B(n8856), .Z(n9085) );
  XNOR U9430 ( .A(n9086), .B(n9085), .Z(n9087) );
  XNOR U9431 ( .A(n9088), .B(n9087), .Z(n8849) );
  NANDN U9432 ( .A(n17375), .B(o[41]), .Z(n8847) );
  OR U9433 ( .A(n8824), .B(n8823), .Z(n8828) );
  OR U9434 ( .A(n8826), .B(n8825), .Z(n8827) );
  NAND U9435 ( .A(n8828), .B(n8827), .Z(n8848) );
  XOR U9436 ( .A(n8847), .B(n8848), .Z(n8850) );
  XNOR U9437 ( .A(n8849), .B(n8850), .Z(n9091) );
  XNOR U9438 ( .A(n9092), .B(n9091), .Z(n9093) );
  AND U9439 ( .A(o[43]), .B(\stack[1][1] ), .Z(n8841) );
  OR U9440 ( .A(n8830), .B(n8829), .Z(n8834) );
  OR U9441 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U9442 ( .A(n8834), .B(n8833), .Z(n8842) );
  XNOR U9443 ( .A(n8841), .B(n8842), .Z(n8844) );
  XOR U9444 ( .A(n8843), .B(n8844), .Z(n8835) );
  NANDN U9445 ( .A(n8836), .B(n8835), .Z(n8838) );
  XOR U9446 ( .A(n8836), .B(n8835), .Z(n15782) );
  AND U9447 ( .A(o[44]), .B(\stack[1][0] ), .Z(n15783) );
  OR U9448 ( .A(n15782), .B(n15783), .Z(n8837) );
  AND U9449 ( .A(n8838), .B(n8837), .Z(n8840) );
  OR U9450 ( .A(n8839), .B(n8840), .Z(n9098) );
  XNOR U9451 ( .A(n8840), .B(n8839), .Z(n15743) );
  NANDN U9452 ( .A(n2969), .B(o[44]), .Z(n9358) );
  OR U9453 ( .A(n8842), .B(n8841), .Z(n8846) );
  OR U9454 ( .A(n8844), .B(n8843), .Z(n8845) );
  NAND U9455 ( .A(n8846), .B(n8845), .Z(n9356) );
  NANDN U9456 ( .A(n17375), .B(o[42]), .Z(n9352) );
  NANDN U9457 ( .A(n8848), .B(n8847), .Z(n8852) );
  NANDN U9458 ( .A(n8850), .B(n8849), .Z(n8851) );
  NAND U9459 ( .A(n8852), .B(n8851), .Z(n9350) );
  NANDN U9460 ( .A(n17296), .B(o[40]), .Z(n9346) );
  NANDN U9461 ( .A(n8854), .B(n8853), .Z(n8858) );
  NANDN U9462 ( .A(n8856), .B(n8855), .Z(n8857) );
  NAND U9463 ( .A(n8858), .B(n8857), .Z(n9344) );
  NANDN U9464 ( .A(n17219), .B(o[38]), .Z(n9340) );
  NANDN U9465 ( .A(n8860), .B(n8859), .Z(n8864) );
  NANDN U9466 ( .A(n8862), .B(n8861), .Z(n8863) );
  NAND U9467 ( .A(n8864), .B(n8863), .Z(n9338) );
  NANDN U9468 ( .A(n17145), .B(o[36]), .Z(n9334) );
  NANDN U9469 ( .A(n8866), .B(n8865), .Z(n8870) );
  NANDN U9470 ( .A(n8868), .B(n8867), .Z(n8869) );
  NAND U9471 ( .A(n8870), .B(n8869), .Z(n9332) );
  NANDN U9472 ( .A(n2972), .B(o[34]), .Z(n9328) );
  NANDN U9473 ( .A(n8872), .B(n8871), .Z(n8876) );
  NANDN U9474 ( .A(n8874), .B(n8873), .Z(n8875) );
  NAND U9475 ( .A(n8876), .B(n8875), .Z(n9326) );
  AND U9476 ( .A(o[32]), .B(\stack[1][13] ), .Z(n9138) );
  OR U9477 ( .A(n8878), .B(n8877), .Z(n8882) );
  OR U9478 ( .A(n8880), .B(n8879), .Z(n8881) );
  AND U9479 ( .A(n8882), .B(n8881), .Z(n9135) );
  OR U9480 ( .A(n8884), .B(n8883), .Z(n8888) );
  NANDN U9481 ( .A(n8886), .B(n8885), .Z(n8887) );
  AND U9482 ( .A(n8888), .B(n8887), .Z(n9319) );
  AND U9483 ( .A(o[31]), .B(\stack[1][14] ), .Z(n9320) );
  XNOR U9484 ( .A(n9319), .B(n9320), .Z(n9322) );
  NANDN U9485 ( .A(n8890), .B(n8889), .Z(n8894) );
  OR U9486 ( .A(n8892), .B(n8891), .Z(n8893) );
  NAND U9487 ( .A(n8894), .B(n8893), .Z(n9148) );
  ANDN U9488 ( .B(o[29]), .A(n2977), .Z(n9147) );
  XNOR U9489 ( .A(n9148), .B(n9147), .Z(n9149) );
  NANDN U9490 ( .A(n16826), .B(o[28]), .Z(n9316) );
  NANDN U9491 ( .A(n8896), .B(n8895), .Z(n8900) );
  NANDN U9492 ( .A(n8898), .B(n8897), .Z(n8899) );
  AND U9493 ( .A(n8900), .B(n8899), .Z(n9313) );
  NANDN U9494 ( .A(n16746), .B(o[26]), .Z(n9310) );
  NANDN U9495 ( .A(n8902), .B(n8901), .Z(n8906) );
  NANDN U9496 ( .A(n8904), .B(n8903), .Z(n8905) );
  NAND U9497 ( .A(n8906), .B(n8905), .Z(n9308) );
  NANDN U9498 ( .A(n2978), .B(o[24]), .Z(n9304) );
  NANDN U9499 ( .A(n8908), .B(n8907), .Z(n8912) );
  NANDN U9500 ( .A(n8910), .B(n8909), .Z(n8911) );
  NAND U9501 ( .A(n8912), .B(n8911), .Z(n9302) );
  AND U9502 ( .A(\stack[1][23] ), .B(o[22]), .Z(n9174) );
  OR U9503 ( .A(n8914), .B(n8913), .Z(n8918) );
  OR U9504 ( .A(n8916), .B(n8915), .Z(n8917) );
  AND U9505 ( .A(n8918), .B(n8917), .Z(n9171) );
  OR U9506 ( .A(n8920), .B(n8919), .Z(n8924) );
  NANDN U9507 ( .A(n8922), .B(n8921), .Z(n8923) );
  AND U9508 ( .A(n8924), .B(n8923), .Z(n9295) );
  AND U9509 ( .A(\stack[1][24] ), .B(o[21]), .Z(n9296) );
  XNOR U9510 ( .A(n9295), .B(n9296), .Z(n9298) );
  NANDN U9511 ( .A(n8926), .B(n8925), .Z(n8930) );
  OR U9512 ( .A(n8928), .B(n8927), .Z(n8929) );
  NAND U9513 ( .A(n8930), .B(n8929), .Z(n9184) );
  ANDN U9514 ( .B(o[19]), .A(n2983), .Z(n9183) );
  XNOR U9515 ( .A(n9184), .B(n9183), .Z(n9185) );
  NANDN U9516 ( .A(n3012), .B(\stack[1][27] ), .Z(n9192) );
  NANDN U9517 ( .A(n8932), .B(n8931), .Z(n8936) );
  NANDN U9518 ( .A(n8934), .B(n8933), .Z(n8935) );
  AND U9519 ( .A(n8936), .B(n8935), .Z(n9189) );
  AND U9520 ( .A(\stack[1][28] ), .B(o[17]), .Z(n9289) );
  OR U9521 ( .A(n8938), .B(n8937), .Z(n8942) );
  OR U9522 ( .A(n8940), .B(n8939), .Z(n8941) );
  NAND U9523 ( .A(n8942), .B(n8941), .Z(n9290) );
  XNOR U9524 ( .A(n9289), .B(n9290), .Z(n9292) );
  NANDN U9525 ( .A(n3009), .B(\stack[1][30] ), .Z(n9202) );
  OR U9526 ( .A(n8944), .B(n8943), .Z(n8948) );
  OR U9527 ( .A(n8946), .B(n8945), .Z(n8947) );
  AND U9528 ( .A(n8948), .B(n8947), .Z(n9201) );
  XNOR U9529 ( .A(n9202), .B(n9201), .Z(n9203) );
  OR U9530 ( .A(n8950), .B(n8949), .Z(n8954) );
  OR U9531 ( .A(n8952), .B(n8951), .Z(n8953) );
  NAND U9532 ( .A(n8954), .B(n8953), .Z(n9208) );
  OR U9533 ( .A(n8956), .B(n8955), .Z(n8960) );
  OR U9534 ( .A(n8958), .B(n8957), .Z(n8959) );
  AND U9535 ( .A(n8960), .B(n8959), .Z(n9213) );
  AND U9536 ( .A(\stack[1][32] ), .B(o[13]), .Z(n9214) );
  XNOR U9537 ( .A(n9213), .B(n9214), .Z(n9216) );
  NANDN U9538 ( .A(n8962), .B(n8961), .Z(n8966) );
  OR U9539 ( .A(n8964), .B(n8963), .Z(n8965) );
  NAND U9540 ( .A(n8966), .B(n8965), .Z(n9278) );
  ANDN U9541 ( .B(\stack[1][38] ), .A(n3001), .Z(n9234) );
  NANDN U9542 ( .A(n8968), .B(n8967), .Z(n8972) );
  NANDN U9543 ( .A(n8970), .B(n8969), .Z(n8971) );
  AND U9544 ( .A(n8972), .B(n8971), .Z(n9231) );
  AND U9545 ( .A(\stack[1][40] ), .B(o[5]), .Z(n9262) );
  OR U9546 ( .A(n8974), .B(n8973), .Z(n8978) );
  NANDN U9547 ( .A(n8976), .B(n8975), .Z(n8977) );
  AND U9548 ( .A(n8978), .B(n8977), .Z(n9259) );
  AND U9549 ( .A(\stack[1][41] ), .B(o[4]), .Z(n9240) );
  AND U9550 ( .A(\stack[1][42] ), .B(o[3]), .Z(n9256) );
  NANDN U9551 ( .A(n8979), .B(n9243), .Z(n8980) );
  AND U9552 ( .A(n8981), .B(n8980), .Z(n8985) );
  OR U9553 ( .A(n8983), .B(n8982), .Z(n8984) );
  AND U9554 ( .A(n8985), .B(n8984), .Z(n9253) );
  AND U9555 ( .A(\stack[1][45] ), .B(o[1]), .Z(n9251) );
  ANDN U9556 ( .B(n9251), .A(n8986), .Z(n9522) );
  XNOR U9557 ( .A(n9522), .B(n9243), .Z(n8988) );
  NAND U9558 ( .A(\stack[1][45] ), .B(o[0]), .Z(n9250) );
  NANDN U9559 ( .A(n8987), .B(n9250), .Z(n9245) );
  NAND U9560 ( .A(n8988), .B(n9245), .Z(n9247) );
  AND U9561 ( .A(\stack[1][43] ), .B(o[2]), .Z(n9246) );
  XNOR U9562 ( .A(n9247), .B(n9246), .Z(n9254) );
  XOR U9563 ( .A(n9253), .B(n9254), .Z(n9255) );
  XOR U9564 ( .A(n9256), .B(n9255), .Z(n9238) );
  OR U9565 ( .A(n8990), .B(n8989), .Z(n8994) );
  NANDN U9566 ( .A(n8992), .B(n8991), .Z(n8993) );
  AND U9567 ( .A(n8994), .B(n8993), .Z(n9237) );
  XOR U9568 ( .A(n9238), .B(n9237), .Z(n9239) );
  XOR U9569 ( .A(n9240), .B(n9239), .Z(n9260) );
  XOR U9570 ( .A(n9259), .B(n9260), .Z(n9261) );
  XOR U9571 ( .A(n9262), .B(n9261), .Z(n9267) );
  NANDN U9572 ( .A(n8996), .B(n8995), .Z(n9000) );
  NANDN U9573 ( .A(n8998), .B(n8997), .Z(n8999) );
  NAND U9574 ( .A(n9000), .B(n8999), .Z(n9266) );
  NANDN U9575 ( .A(n3000), .B(\stack[1][39] ), .Z(n9265) );
  XNOR U9576 ( .A(n9266), .B(n9265), .Z(n9268) );
  XNOR U9577 ( .A(n9267), .B(n9268), .Z(n9232) );
  XNOR U9578 ( .A(n9231), .B(n9232), .Z(n9233) );
  OR U9579 ( .A(n9002), .B(n9001), .Z(n9006) );
  NANDN U9580 ( .A(n9004), .B(n9003), .Z(n9005) );
  NAND U9581 ( .A(n9006), .B(n9005), .Z(n9272) );
  ANDN U9582 ( .B(\stack[1][37] ), .A(n3002), .Z(n9271) );
  XOR U9583 ( .A(n9272), .B(n9271), .Z(n9274) );
  OR U9584 ( .A(n9008), .B(n9007), .Z(n9012) );
  NANDN U9585 ( .A(n9010), .B(n9009), .Z(n9011) );
  AND U9586 ( .A(n9012), .B(n9011), .Z(n9225) );
  AND U9587 ( .A(\stack[1][36] ), .B(o[9]), .Z(n9226) );
  XNOR U9588 ( .A(n9225), .B(n9226), .Z(n9228) );
  XOR U9589 ( .A(n9227), .B(n9228), .Z(n9277) );
  XOR U9590 ( .A(n9278), .B(n9277), .Z(n9280) );
  AND U9591 ( .A(\stack[1][35] ), .B(o[10]), .Z(n9279) );
  XNOR U9592 ( .A(n9280), .B(n9279), .Z(n9221) );
  AND U9593 ( .A(\stack[1][34] ), .B(o[11]), .Z(n9219) );
  NANDN U9594 ( .A(n9014), .B(n9013), .Z(n9018) );
  OR U9595 ( .A(n9016), .B(n9015), .Z(n9017) );
  NAND U9596 ( .A(n9018), .B(n9017), .Z(n9220) );
  XNOR U9597 ( .A(n9219), .B(n9220), .Z(n9222) );
  XNOR U9598 ( .A(n9221), .B(n9222), .Z(n9284) );
  OR U9599 ( .A(n9020), .B(n9019), .Z(n9024) );
  OR U9600 ( .A(n9022), .B(n9021), .Z(n9023) );
  NAND U9601 ( .A(n9024), .B(n9023), .Z(n9283) );
  XNOR U9602 ( .A(n9284), .B(n9283), .Z(n9285) );
  AND U9603 ( .A(\stack[1][33] ), .B(o[12]), .Z(n9286) );
  XNOR U9604 ( .A(n9216), .B(n9215), .Z(n9207) );
  XOR U9605 ( .A(n9208), .B(n9207), .Z(n9210) );
  NANDN U9606 ( .A(n3008), .B(\stack[1][31] ), .Z(n9209) );
  XNOR U9607 ( .A(n9210), .B(n9209), .Z(n9204) );
  NANDN U9608 ( .A(n9026), .B(n9025), .Z(n9030) );
  NANDN U9609 ( .A(n9028), .B(n9027), .Z(n9029) );
  AND U9610 ( .A(n9030), .B(n9029), .Z(n9196) );
  XNOR U9611 ( .A(n9195), .B(n9196), .Z(n9198) );
  AND U9612 ( .A(\stack[1][29] ), .B(o[16]), .Z(n9197) );
  XNOR U9613 ( .A(n9198), .B(n9197), .Z(n9291) );
  XOR U9614 ( .A(n9292), .B(n9291), .Z(n9190) );
  XNOR U9615 ( .A(n9189), .B(n9190), .Z(n9191) );
  XOR U9616 ( .A(n9185), .B(n9186), .Z(n9177) );
  OR U9617 ( .A(n9032), .B(n9031), .Z(n9036) );
  NANDN U9618 ( .A(n9034), .B(n9033), .Z(n9035) );
  AND U9619 ( .A(n9036), .B(n9035), .Z(n9178) );
  XOR U9620 ( .A(n9177), .B(n9178), .Z(n9180) );
  AND U9621 ( .A(\stack[1][25] ), .B(o[20]), .Z(n9179) );
  XOR U9622 ( .A(n9180), .B(n9179), .Z(n9297) );
  XOR U9623 ( .A(n9298), .B(n9297), .Z(n9172) );
  XOR U9624 ( .A(n9171), .B(n9172), .Z(n9173) );
  XOR U9625 ( .A(n9174), .B(n9173), .Z(n9168) );
  AND U9626 ( .A(o[23]), .B(\stack[1][22] ), .Z(n9165) );
  OR U9627 ( .A(n9038), .B(n9037), .Z(n9042) );
  IV U9628 ( .A(n9039), .Z(n16633) );
  OR U9629 ( .A(n9040), .B(n16633), .Z(n9041) );
  NAND U9630 ( .A(n9042), .B(n9041), .Z(n9166) );
  XNOR U9631 ( .A(n9165), .B(n9166), .Z(n9167) );
  XOR U9632 ( .A(n9168), .B(n9167), .Z(n9301) );
  XNOR U9633 ( .A(n9302), .B(n9301), .Z(n9303) );
  XNOR U9634 ( .A(n9304), .B(n9303), .Z(n9161) );
  NANDN U9635 ( .A(n3019), .B(\stack[1][20] ), .Z(n9159) );
  OR U9636 ( .A(n9044), .B(n9043), .Z(n9048) );
  OR U9637 ( .A(n9046), .B(n9045), .Z(n9047) );
  NAND U9638 ( .A(n9048), .B(n9047), .Z(n9160) );
  XOR U9639 ( .A(n9159), .B(n9160), .Z(n9162) );
  XNOR U9640 ( .A(n9161), .B(n9162), .Z(n9307) );
  XNOR U9641 ( .A(n9308), .B(n9307), .Z(n9309) );
  XNOR U9642 ( .A(n9310), .B(n9309), .Z(n9155) );
  NANDN U9643 ( .A(n16786), .B(o[27]), .Z(n9153) );
  OR U9644 ( .A(n9050), .B(n9049), .Z(n9054) );
  OR U9645 ( .A(n9052), .B(n9051), .Z(n9053) );
  NAND U9646 ( .A(n9054), .B(n9053), .Z(n9154) );
  XOR U9647 ( .A(n9153), .B(n9154), .Z(n9156) );
  XNOR U9648 ( .A(n9155), .B(n9156), .Z(n9314) );
  XNOR U9649 ( .A(n9313), .B(n9314), .Z(n9315) );
  XOR U9650 ( .A(n9149), .B(n9150), .Z(n9141) );
  OR U9651 ( .A(n9056), .B(n9055), .Z(n9060) );
  NANDN U9652 ( .A(n9058), .B(n9057), .Z(n9059) );
  AND U9653 ( .A(n9060), .B(n9059), .Z(n9142) );
  XOR U9654 ( .A(n9141), .B(n9142), .Z(n9144) );
  AND U9655 ( .A(o[30]), .B(\stack[1][15] ), .Z(n9143) );
  XOR U9656 ( .A(n9144), .B(n9143), .Z(n9321) );
  XOR U9657 ( .A(n9322), .B(n9321), .Z(n9136) );
  XOR U9658 ( .A(n9135), .B(n9136), .Z(n9137) );
  XOR U9659 ( .A(n9138), .B(n9137), .Z(n9132) );
  AND U9660 ( .A(o[33]), .B(\stack[1][12] ), .Z(n9129) );
  OR U9661 ( .A(n9062), .B(n9061), .Z(n9066) );
  OR U9662 ( .A(n9064), .B(n9063), .Z(n9065) );
  NAND U9663 ( .A(n9066), .B(n9065), .Z(n9130) );
  XNOR U9664 ( .A(n9129), .B(n9130), .Z(n9131) );
  XOR U9665 ( .A(n9132), .B(n9131), .Z(n9325) );
  XNOR U9666 ( .A(n9326), .B(n9325), .Z(n9327) );
  XNOR U9667 ( .A(n9328), .B(n9327), .Z(n9125) );
  NANDN U9668 ( .A(n17101), .B(o[35]), .Z(n9123) );
  OR U9669 ( .A(n9068), .B(n9067), .Z(n9072) );
  OR U9670 ( .A(n9070), .B(n9069), .Z(n9071) );
  NAND U9671 ( .A(n9072), .B(n9071), .Z(n9124) );
  XOR U9672 ( .A(n9123), .B(n9124), .Z(n9126) );
  XNOR U9673 ( .A(n9125), .B(n9126), .Z(n9331) );
  XNOR U9674 ( .A(n9332), .B(n9331), .Z(n9333) );
  XNOR U9675 ( .A(n9334), .B(n9333), .Z(n9119) );
  NANDN U9676 ( .A(n17179), .B(o[37]), .Z(n9117) );
  OR U9677 ( .A(n9074), .B(n9073), .Z(n9078) );
  OR U9678 ( .A(n9076), .B(n9075), .Z(n9077) );
  NAND U9679 ( .A(n9078), .B(n9077), .Z(n9118) );
  XOR U9680 ( .A(n9117), .B(n9118), .Z(n9120) );
  XNOR U9681 ( .A(n9119), .B(n9120), .Z(n9337) );
  XNOR U9682 ( .A(n9338), .B(n9337), .Z(n9339) );
  XNOR U9683 ( .A(n9340), .B(n9339), .Z(n9113) );
  NANDN U9684 ( .A(n17256), .B(o[39]), .Z(n9111) );
  OR U9685 ( .A(n9080), .B(n9079), .Z(n9084) );
  OR U9686 ( .A(n9082), .B(n9081), .Z(n9083) );
  NAND U9687 ( .A(n9084), .B(n9083), .Z(n9112) );
  XOR U9688 ( .A(n9111), .B(n9112), .Z(n9114) );
  XNOR U9689 ( .A(n9113), .B(n9114), .Z(n9343) );
  XNOR U9690 ( .A(n9344), .B(n9343), .Z(n9345) );
  XNOR U9691 ( .A(n9346), .B(n9345), .Z(n9107) );
  AND U9692 ( .A(o[41]), .B(\stack[1][4] ), .Z(n9105) );
  OR U9693 ( .A(n9086), .B(n9085), .Z(n9090) );
  OR U9694 ( .A(n9088), .B(n9087), .Z(n9089) );
  NAND U9695 ( .A(n9090), .B(n9089), .Z(n9106) );
  XNOR U9696 ( .A(n9105), .B(n9106), .Z(n9108) );
  XNOR U9697 ( .A(n9107), .B(n9108), .Z(n9349) );
  XNOR U9698 ( .A(n9350), .B(n9349), .Z(n9351) );
  XOR U9699 ( .A(n9352), .B(n9351), .Z(n9102) );
  AND U9700 ( .A(o[43]), .B(\stack[1][2] ), .Z(n9099) );
  OR U9701 ( .A(n9092), .B(n9091), .Z(n9096) );
  OR U9702 ( .A(n9094), .B(n9093), .Z(n9095) );
  NAND U9703 ( .A(n9096), .B(n9095), .Z(n9100) );
  XOR U9704 ( .A(n9099), .B(n9100), .Z(n9101) );
  XNOR U9705 ( .A(n9102), .B(n9101), .Z(n9355) );
  XNOR U9706 ( .A(n9356), .B(n9355), .Z(n9357) );
  XOR U9707 ( .A(n9358), .B(n9357), .Z(n15744) );
  OR U9708 ( .A(n15743), .B(n15744), .Z(n9097) );
  AND U9709 ( .A(n9098), .B(n9097), .Z(n9362) );
  NANDN U9710 ( .A(n2970), .B(o[44]), .Z(n9631) );
  OR U9711 ( .A(n9100), .B(n9099), .Z(n9104) );
  NANDN U9712 ( .A(n9102), .B(n9101), .Z(n9103) );
  NAND U9713 ( .A(n9104), .B(n9103), .Z(n9629) );
  NANDN U9714 ( .A(n2971), .B(o[42]), .Z(n9625) );
  OR U9715 ( .A(n9106), .B(n9105), .Z(n9110) );
  NANDN U9716 ( .A(n9108), .B(n9107), .Z(n9109) );
  NAND U9717 ( .A(n9110), .B(n9109), .Z(n9623) );
  NANDN U9718 ( .A(n17256), .B(o[40]), .Z(n9619) );
  NANDN U9719 ( .A(n9112), .B(n9111), .Z(n9116) );
  NANDN U9720 ( .A(n9114), .B(n9113), .Z(n9115) );
  NAND U9721 ( .A(n9116), .B(n9115), .Z(n9617) );
  NANDN U9722 ( .A(n17179), .B(o[38]), .Z(n9613) );
  NANDN U9723 ( .A(n9118), .B(n9117), .Z(n9122) );
  NANDN U9724 ( .A(n9120), .B(n9119), .Z(n9121) );
  NAND U9725 ( .A(n9122), .B(n9121), .Z(n9611) );
  NANDN U9726 ( .A(n17101), .B(o[36]), .Z(n9607) );
  NANDN U9727 ( .A(n9124), .B(n9123), .Z(n9128) );
  NANDN U9728 ( .A(n9126), .B(n9125), .Z(n9127) );
  NAND U9729 ( .A(n9128), .B(n9127), .Z(n9605) );
  AND U9730 ( .A(o[34]), .B(\stack[1][12] ), .Z(n9406) );
  OR U9731 ( .A(n9130), .B(n9129), .Z(n9134) );
  OR U9732 ( .A(n9132), .B(n9131), .Z(n9133) );
  AND U9733 ( .A(n9134), .B(n9133), .Z(n9403) );
  OR U9734 ( .A(n9136), .B(n9135), .Z(n9140) );
  NANDN U9735 ( .A(n9138), .B(n9137), .Z(n9139) );
  AND U9736 ( .A(n9140), .B(n9139), .Z(n9598) );
  AND U9737 ( .A(o[33]), .B(\stack[1][13] ), .Z(n9599) );
  XNOR U9738 ( .A(n9598), .B(n9599), .Z(n9601) );
  NANDN U9739 ( .A(n9142), .B(n9141), .Z(n9146) );
  OR U9740 ( .A(n9144), .B(n9143), .Z(n9145) );
  NAND U9741 ( .A(n9146), .B(n9145), .Z(n9416) );
  ANDN U9742 ( .B(o[31]), .A(n2976), .Z(n9415) );
  XNOR U9743 ( .A(n9416), .B(n9415), .Z(n9417) );
  NANDN U9744 ( .A(n2977), .B(o[30]), .Z(n9595) );
  NANDN U9745 ( .A(n9148), .B(n9147), .Z(n9152) );
  NANDN U9746 ( .A(n9150), .B(n9149), .Z(n9151) );
  AND U9747 ( .A(n9152), .B(n9151), .Z(n9592) );
  NANDN U9748 ( .A(n16786), .B(o[28]), .Z(n9589) );
  NANDN U9749 ( .A(n9154), .B(n9153), .Z(n9158) );
  NANDN U9750 ( .A(n9156), .B(n9155), .Z(n9157) );
  NAND U9751 ( .A(n9158), .B(n9157), .Z(n9587) );
  NANDN U9752 ( .A(n16712), .B(o[26]), .Z(n9583) );
  NANDN U9753 ( .A(n9160), .B(n9159), .Z(n9164) );
  NANDN U9754 ( .A(n9162), .B(n9161), .Z(n9163) );
  NAND U9755 ( .A(n9164), .B(n9163), .Z(n9581) );
  AND U9756 ( .A(o[24]), .B(\stack[1][22] ), .Z(n9577) );
  OR U9757 ( .A(n9166), .B(n9165), .Z(n9170) );
  OR U9758 ( .A(n9168), .B(n9167), .Z(n9169) );
  AND U9759 ( .A(n9170), .B(n9169), .Z(n9574) );
  AND U9760 ( .A(\stack[1][23] ), .B(o[23]), .Z(n16589) );
  OR U9761 ( .A(n9172), .B(n9171), .Z(n9176) );
  NANDN U9762 ( .A(n9174), .B(n9173), .Z(n9175) );
  AND U9763 ( .A(n9176), .B(n9175), .Z(n9439) );
  XNOR U9764 ( .A(n16589), .B(n9439), .Z(n9441) );
  NANDN U9765 ( .A(n9178), .B(n9177), .Z(n9182) );
  OR U9766 ( .A(n9180), .B(n9179), .Z(n9181) );
  NAND U9767 ( .A(n9182), .B(n9181), .Z(n9445) );
  ANDN U9768 ( .B(o[21]), .A(n2982), .Z(n9444) );
  XNOR U9769 ( .A(n9445), .B(n9444), .Z(n9446) );
  NANDN U9770 ( .A(n3014), .B(\stack[1][26] ), .Z(n9453) );
  NANDN U9771 ( .A(n9184), .B(n9183), .Z(n9188) );
  NANDN U9772 ( .A(n9186), .B(n9185), .Z(n9187) );
  AND U9773 ( .A(n9188), .B(n9187), .Z(n9450) );
  AND U9774 ( .A(\stack[1][27] ), .B(o[19]), .Z(n9562) );
  OR U9775 ( .A(n9190), .B(n9189), .Z(n9194) );
  OR U9776 ( .A(n9192), .B(n9191), .Z(n9193) );
  NAND U9777 ( .A(n9194), .B(n9193), .Z(n9563) );
  XNOR U9778 ( .A(n9562), .B(n9563), .Z(n9565) );
  OR U9779 ( .A(n9196), .B(n9195), .Z(n9200) );
  OR U9780 ( .A(n9198), .B(n9197), .Z(n9199) );
  NAND U9781 ( .A(n9200), .B(n9199), .Z(n9463) );
  ANDN U9782 ( .B(o[17]), .A(n2986), .Z(n9462) );
  XNOR U9783 ( .A(n9463), .B(n9462), .Z(n9464) );
  NANDN U9784 ( .A(n3010), .B(\stack[1][30] ), .Z(n9471) );
  OR U9785 ( .A(n9202), .B(n9201), .Z(n9206) );
  OR U9786 ( .A(n9204), .B(n9203), .Z(n9205) );
  AND U9787 ( .A(n9206), .B(n9205), .Z(n9468) );
  AND U9788 ( .A(\stack[1][31] ), .B(o[15]), .Z(n9556) );
  NANDN U9789 ( .A(n9208), .B(n9207), .Z(n9212) );
  OR U9790 ( .A(n9210), .B(n9209), .Z(n9211) );
  NAND U9791 ( .A(n9212), .B(n9211), .Z(n9557) );
  XNOR U9792 ( .A(n9556), .B(n9557), .Z(n9559) );
  OR U9793 ( .A(n9214), .B(n9213), .Z(n9218) );
  OR U9794 ( .A(n9216), .B(n9215), .Z(n9217) );
  AND U9795 ( .A(n9218), .B(n9217), .Z(n9474) );
  NANDN U9796 ( .A(n3006), .B(\stack[1][34] ), .Z(n9489) );
  OR U9797 ( .A(n9220), .B(n9219), .Z(n9224) );
  OR U9798 ( .A(n9222), .B(n9221), .Z(n9223) );
  NAND U9799 ( .A(n9224), .B(n9223), .Z(n9487) );
  NANDN U9800 ( .A(n3004), .B(\stack[1][36] ), .Z(n9553) );
  OR U9801 ( .A(n9226), .B(n9225), .Z(n9230) );
  NANDN U9802 ( .A(n9228), .B(n9227), .Z(n9229) );
  NAND U9803 ( .A(n9230), .B(n9229), .Z(n9551) );
  ANDN U9804 ( .B(\stack[1][38] ), .A(n3002), .Z(n9507) );
  OR U9805 ( .A(n9232), .B(n9231), .Z(n9236) );
  OR U9806 ( .A(n9234), .B(n9233), .Z(n9235) );
  AND U9807 ( .A(n9236), .B(n9235), .Z(n9504) );
  AND U9808 ( .A(\stack[1][41] ), .B(o[5]), .Z(n9541) );
  OR U9809 ( .A(n9238), .B(n9237), .Z(n9242) );
  NANDN U9810 ( .A(n9240), .B(n9239), .Z(n9241) );
  AND U9811 ( .A(n9242), .B(n9241), .Z(n9538) );
  AND U9812 ( .A(\stack[1][42] ), .B(o[4]), .Z(n9519) );
  AND U9813 ( .A(\stack[1][43] ), .B(o[3]), .Z(n9535) );
  NANDN U9814 ( .A(n9243), .B(n9522), .Z(n9244) );
  AND U9815 ( .A(n9245), .B(n9244), .Z(n9249) );
  OR U9816 ( .A(n9247), .B(n9246), .Z(n9248) );
  AND U9817 ( .A(n9249), .B(n9248), .Z(n9532) );
  AND U9818 ( .A(\stack[1][46] ), .B(o[1]), .Z(n9530) );
  ANDN U9819 ( .B(n9530), .A(n9250), .Z(n9780) );
  XNOR U9820 ( .A(n9780), .B(n9522), .Z(n9252) );
  NAND U9821 ( .A(\stack[1][46] ), .B(o[0]), .Z(n9529) );
  NANDN U9822 ( .A(n9251), .B(n9529), .Z(n9524) );
  NAND U9823 ( .A(n9252), .B(n9524), .Z(n9526) );
  AND U9824 ( .A(\stack[1][44] ), .B(o[2]), .Z(n9525) );
  XNOR U9825 ( .A(n9526), .B(n9525), .Z(n9533) );
  XOR U9826 ( .A(n9532), .B(n9533), .Z(n9534) );
  XOR U9827 ( .A(n9535), .B(n9534), .Z(n9517) );
  OR U9828 ( .A(n9254), .B(n9253), .Z(n9258) );
  NANDN U9829 ( .A(n9256), .B(n9255), .Z(n9257) );
  AND U9830 ( .A(n9258), .B(n9257), .Z(n9516) );
  XOR U9831 ( .A(n9517), .B(n9516), .Z(n9518) );
  XOR U9832 ( .A(n9519), .B(n9518), .Z(n9539) );
  XNOR U9833 ( .A(n9538), .B(n9539), .Z(n9540) );
  OR U9834 ( .A(n9260), .B(n9259), .Z(n9264) );
  NANDN U9835 ( .A(n9262), .B(n9261), .Z(n9263) );
  NAND U9836 ( .A(n9264), .B(n9263), .Z(n9511) );
  ANDN U9837 ( .B(o[6]), .A(n15935), .Z(n9510) );
  XNOR U9838 ( .A(n9511), .B(n9510), .Z(n9513) );
  XNOR U9839 ( .A(n9512), .B(n9513), .Z(n9545) );
  ANDN U9840 ( .B(\stack[1][39] ), .A(n3001), .Z(n9544) );
  XNOR U9841 ( .A(n9545), .B(n9544), .Z(n9546) );
  OR U9842 ( .A(n9266), .B(n9265), .Z(n9270) );
  NANDN U9843 ( .A(n9268), .B(n9267), .Z(n9269) );
  AND U9844 ( .A(n9270), .B(n9269), .Z(n9547) );
  XNOR U9845 ( .A(n9546), .B(n9547), .Z(n9505) );
  XOR U9846 ( .A(n9504), .B(n9505), .Z(n9506) );
  XOR U9847 ( .A(n9507), .B(n9506), .Z(n9501) );
  AND U9848 ( .A(\stack[1][37] ), .B(o[9]), .Z(n9498) );
  NANDN U9849 ( .A(n9272), .B(n9271), .Z(n9276) );
  NANDN U9850 ( .A(n9274), .B(n9273), .Z(n9275) );
  NAND U9851 ( .A(n9276), .B(n9275), .Z(n9499) );
  XNOR U9852 ( .A(n9498), .B(n9499), .Z(n9500) );
  XOR U9853 ( .A(n9501), .B(n9500), .Z(n9550) );
  XNOR U9854 ( .A(n9551), .B(n9550), .Z(n9552) );
  XNOR U9855 ( .A(n9553), .B(n9552), .Z(n9494) );
  NANDN U9856 ( .A(n2992), .B(o[11]), .Z(n9492) );
  NANDN U9857 ( .A(n9278), .B(n9277), .Z(n9282) );
  NANDN U9858 ( .A(n9280), .B(n9279), .Z(n9281) );
  NAND U9859 ( .A(n9282), .B(n9281), .Z(n9493) );
  XOR U9860 ( .A(n9492), .B(n9493), .Z(n9495) );
  XNOR U9861 ( .A(n9494), .B(n9495), .Z(n9486) );
  XNOR U9862 ( .A(n9487), .B(n9486), .Z(n9488) );
  XNOR U9863 ( .A(n9489), .B(n9488), .Z(n9482) );
  OR U9864 ( .A(n9284), .B(n9283), .Z(n9288) );
  OR U9865 ( .A(n9286), .B(n9285), .Z(n9287) );
  AND U9866 ( .A(n9288), .B(n9287), .Z(n9480) );
  AND U9867 ( .A(\stack[1][33] ), .B(o[13]), .Z(n9481) );
  XNOR U9868 ( .A(n9480), .B(n9481), .Z(n9483) );
  XOR U9869 ( .A(n9482), .B(n9483), .Z(n9475) );
  XOR U9870 ( .A(n9474), .B(n9475), .Z(n9476) );
  AND U9871 ( .A(\stack[1][32] ), .B(o[14]), .Z(n9477) );
  XOR U9872 ( .A(n9476), .B(n9477), .Z(n9558) );
  XOR U9873 ( .A(n9559), .B(n9558), .Z(n9469) );
  XNOR U9874 ( .A(n9468), .B(n9469), .Z(n9470) );
  XOR U9875 ( .A(n9464), .B(n9465), .Z(n9456) );
  OR U9876 ( .A(n9290), .B(n9289), .Z(n9294) );
  OR U9877 ( .A(n9292), .B(n9291), .Z(n9293) );
  AND U9878 ( .A(n9294), .B(n9293), .Z(n9457) );
  XOR U9879 ( .A(n9456), .B(n9457), .Z(n9459) );
  AND U9880 ( .A(\stack[1][28] ), .B(o[18]), .Z(n9458) );
  XNOR U9881 ( .A(n9459), .B(n9458), .Z(n9564) );
  XOR U9882 ( .A(n9565), .B(n9564), .Z(n9451) );
  XNOR U9883 ( .A(n9450), .B(n9451), .Z(n9452) );
  XOR U9884 ( .A(n9446), .B(n9447), .Z(n9568) );
  OR U9885 ( .A(n9296), .B(n9295), .Z(n9300) );
  NANDN U9886 ( .A(n9298), .B(n9297), .Z(n9299) );
  AND U9887 ( .A(n9300), .B(n9299), .Z(n9569) );
  XOR U9888 ( .A(n9568), .B(n9569), .Z(n9571) );
  AND U9889 ( .A(\stack[1][24] ), .B(o[22]), .Z(n9570) );
  XOR U9890 ( .A(n9571), .B(n9570), .Z(n9440) );
  XOR U9891 ( .A(n9441), .B(n9440), .Z(n9575) );
  XOR U9892 ( .A(n9574), .B(n9575), .Z(n9576) );
  XOR U9893 ( .A(n9577), .B(n9576), .Z(n9436) );
  AND U9894 ( .A(o[25]), .B(\stack[1][21] ), .Z(n9433) );
  OR U9895 ( .A(n9302), .B(n9301), .Z(n9306) );
  OR U9896 ( .A(n9304), .B(n9303), .Z(n9305) );
  NAND U9897 ( .A(n9306), .B(n9305), .Z(n9434) );
  XNOR U9898 ( .A(n9433), .B(n9434), .Z(n9435) );
  XOR U9899 ( .A(n9436), .B(n9435), .Z(n9580) );
  XNOR U9900 ( .A(n9581), .B(n9580), .Z(n9582) );
  XNOR U9901 ( .A(n9583), .B(n9582), .Z(n9429) );
  NANDN U9902 ( .A(n16746), .B(o[27]), .Z(n9427) );
  OR U9903 ( .A(n9308), .B(n9307), .Z(n9312) );
  OR U9904 ( .A(n9310), .B(n9309), .Z(n9311) );
  NAND U9905 ( .A(n9312), .B(n9311), .Z(n9428) );
  XOR U9906 ( .A(n9427), .B(n9428), .Z(n9430) );
  XNOR U9907 ( .A(n9429), .B(n9430), .Z(n9586) );
  XNOR U9908 ( .A(n9587), .B(n9586), .Z(n9588) );
  XNOR U9909 ( .A(n9589), .B(n9588), .Z(n9423) );
  NANDN U9910 ( .A(n16826), .B(o[29]), .Z(n9421) );
  OR U9911 ( .A(n9314), .B(n9313), .Z(n9318) );
  OR U9912 ( .A(n9316), .B(n9315), .Z(n9317) );
  NAND U9913 ( .A(n9318), .B(n9317), .Z(n9422) );
  XOR U9914 ( .A(n9421), .B(n9422), .Z(n9424) );
  XNOR U9915 ( .A(n9423), .B(n9424), .Z(n9593) );
  XNOR U9916 ( .A(n9592), .B(n9593), .Z(n9594) );
  XOR U9917 ( .A(n9417), .B(n9418), .Z(n9409) );
  OR U9918 ( .A(n9320), .B(n9319), .Z(n9324) );
  NANDN U9919 ( .A(n9322), .B(n9321), .Z(n9323) );
  AND U9920 ( .A(n9324), .B(n9323), .Z(n9410) );
  XOR U9921 ( .A(n9409), .B(n9410), .Z(n9412) );
  AND U9922 ( .A(o[32]), .B(\stack[1][14] ), .Z(n9411) );
  XOR U9923 ( .A(n9412), .B(n9411), .Z(n9600) );
  XOR U9924 ( .A(n9601), .B(n9600), .Z(n9404) );
  XOR U9925 ( .A(n9403), .B(n9404), .Z(n9405) );
  XOR U9926 ( .A(n9406), .B(n9405), .Z(n9400) );
  AND U9927 ( .A(o[35]), .B(\stack[1][11] ), .Z(n9397) );
  OR U9928 ( .A(n9326), .B(n9325), .Z(n9330) );
  OR U9929 ( .A(n9328), .B(n9327), .Z(n9329) );
  NAND U9930 ( .A(n9330), .B(n9329), .Z(n9398) );
  XNOR U9931 ( .A(n9397), .B(n9398), .Z(n9399) );
  XOR U9932 ( .A(n9400), .B(n9399), .Z(n9604) );
  XNOR U9933 ( .A(n9605), .B(n9604), .Z(n9606) );
  XNOR U9934 ( .A(n9607), .B(n9606), .Z(n9393) );
  NANDN U9935 ( .A(n17145), .B(o[37]), .Z(n9391) );
  OR U9936 ( .A(n9332), .B(n9331), .Z(n9336) );
  OR U9937 ( .A(n9334), .B(n9333), .Z(n9335) );
  NAND U9938 ( .A(n9336), .B(n9335), .Z(n9392) );
  XOR U9939 ( .A(n9391), .B(n9392), .Z(n9394) );
  XNOR U9940 ( .A(n9393), .B(n9394), .Z(n9610) );
  XNOR U9941 ( .A(n9611), .B(n9610), .Z(n9612) );
  XNOR U9942 ( .A(n9613), .B(n9612), .Z(n9387) );
  NANDN U9943 ( .A(n17219), .B(o[39]), .Z(n9385) );
  OR U9944 ( .A(n9338), .B(n9337), .Z(n9342) );
  OR U9945 ( .A(n9340), .B(n9339), .Z(n9341) );
  NAND U9946 ( .A(n9342), .B(n9341), .Z(n9386) );
  XOR U9947 ( .A(n9385), .B(n9386), .Z(n9388) );
  XNOR U9948 ( .A(n9387), .B(n9388), .Z(n9616) );
  XNOR U9949 ( .A(n9617), .B(n9616), .Z(n9618) );
  XNOR U9950 ( .A(n9619), .B(n9618), .Z(n9381) );
  NANDN U9951 ( .A(n17296), .B(o[41]), .Z(n9379) );
  OR U9952 ( .A(n9344), .B(n9343), .Z(n9348) );
  OR U9953 ( .A(n9346), .B(n9345), .Z(n9347) );
  NAND U9954 ( .A(n9348), .B(n9347), .Z(n9380) );
  XOR U9955 ( .A(n9379), .B(n9380), .Z(n9382) );
  XNOR U9956 ( .A(n9381), .B(n9382), .Z(n9622) );
  XNOR U9957 ( .A(n9623), .B(n9622), .Z(n9624) );
  XNOR U9958 ( .A(n9625), .B(n9624), .Z(n9375) );
  NANDN U9959 ( .A(n17375), .B(o[43]), .Z(n9373) );
  OR U9960 ( .A(n9350), .B(n9349), .Z(n9354) );
  OR U9961 ( .A(n9352), .B(n9351), .Z(n9353) );
  NAND U9962 ( .A(n9354), .B(n9353), .Z(n9374) );
  XOR U9963 ( .A(n9373), .B(n9374), .Z(n9376) );
  XNOR U9964 ( .A(n9375), .B(n9376), .Z(n9628) );
  XNOR U9965 ( .A(n9629), .B(n9628), .Z(n9630) );
  AND U9966 ( .A(o[45]), .B(\stack[1][1] ), .Z(n9367) );
  OR U9967 ( .A(n9356), .B(n9355), .Z(n9360) );
  OR U9968 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U9969 ( .A(n9360), .B(n9359), .Z(n9368) );
  XNOR U9970 ( .A(n9367), .B(n9368), .Z(n9370) );
  XOR U9971 ( .A(n9369), .B(n9370), .Z(n9361) );
  NANDN U9972 ( .A(n9362), .B(n9361), .Z(n9364) );
  XOR U9973 ( .A(n9362), .B(n9361), .Z(n15704) );
  AND U9974 ( .A(o[46]), .B(\stack[1][0] ), .Z(n15705) );
  OR U9975 ( .A(n15704), .B(n15705), .Z(n9363) );
  AND U9976 ( .A(n9364), .B(n9363), .Z(n9366) );
  OR U9977 ( .A(n9365), .B(n9366), .Z(n9635) );
  XNOR U9978 ( .A(n9366), .B(n9365), .Z(n15665) );
  NANDN U9979 ( .A(n2969), .B(o[46]), .Z(n9907) );
  OR U9980 ( .A(n9368), .B(n9367), .Z(n9372) );
  OR U9981 ( .A(n9370), .B(n9369), .Z(n9371) );
  NAND U9982 ( .A(n9372), .B(n9371), .Z(n9905) );
  NANDN U9983 ( .A(n17375), .B(o[44]), .Z(n9901) );
  NANDN U9984 ( .A(n9374), .B(n9373), .Z(n9378) );
  NANDN U9985 ( .A(n9376), .B(n9375), .Z(n9377) );
  NAND U9986 ( .A(n9378), .B(n9377), .Z(n9899) );
  NANDN U9987 ( .A(n17296), .B(o[42]), .Z(n9895) );
  NANDN U9988 ( .A(n9380), .B(n9379), .Z(n9384) );
  NANDN U9989 ( .A(n9382), .B(n9381), .Z(n9383) );
  NAND U9990 ( .A(n9384), .B(n9383), .Z(n9893) );
  NANDN U9991 ( .A(n17219), .B(o[40]), .Z(n9889) );
  NANDN U9992 ( .A(n9386), .B(n9385), .Z(n9390) );
  NANDN U9993 ( .A(n9388), .B(n9387), .Z(n9389) );
  NAND U9994 ( .A(n9390), .B(n9389), .Z(n9887) );
  NANDN U9995 ( .A(n17145), .B(o[38]), .Z(n9883) );
  NANDN U9996 ( .A(n9392), .B(n9391), .Z(n9396) );
  NANDN U9997 ( .A(n9394), .B(n9393), .Z(n9395) );
  NAND U9998 ( .A(n9396), .B(n9395), .Z(n9881) );
  AND U9999 ( .A(o[36]), .B(\stack[1][11] ), .Z(n9669) );
  OR U10000 ( .A(n9398), .B(n9397), .Z(n9402) );
  OR U10001 ( .A(n9400), .B(n9399), .Z(n9401) );
  AND U10002 ( .A(n9402), .B(n9401), .Z(n9666) );
  OR U10003 ( .A(n9404), .B(n9403), .Z(n9408) );
  NANDN U10004 ( .A(n9406), .B(n9405), .Z(n9407) );
  AND U10005 ( .A(n9408), .B(n9407), .Z(n9874) );
  AND U10006 ( .A(o[35]), .B(\stack[1][12] ), .Z(n9875) );
  XNOR U10007 ( .A(n9874), .B(n9875), .Z(n9877) );
  NANDN U10008 ( .A(n9410), .B(n9409), .Z(n9414) );
  OR U10009 ( .A(n9412), .B(n9411), .Z(n9413) );
  NAND U10010 ( .A(n9414), .B(n9413), .Z(n9679) );
  ANDN U10011 ( .B(o[33]), .A(n2975), .Z(n9678) );
  XNOR U10012 ( .A(n9679), .B(n9678), .Z(n9680) );
  NANDN U10013 ( .A(n2976), .B(o[32]), .Z(n9871) );
  NANDN U10014 ( .A(n9416), .B(n9415), .Z(n9420) );
  NANDN U10015 ( .A(n9418), .B(n9417), .Z(n9419) );
  AND U10016 ( .A(n9420), .B(n9419), .Z(n9868) );
  NANDN U10017 ( .A(n16826), .B(o[30]), .Z(n9865) );
  NANDN U10018 ( .A(n9422), .B(n9421), .Z(n9426) );
  NANDN U10019 ( .A(n9424), .B(n9423), .Z(n9425) );
  NAND U10020 ( .A(n9426), .B(n9425), .Z(n9863) );
  NANDN U10021 ( .A(n16746), .B(o[28]), .Z(n9859) );
  NANDN U10022 ( .A(n9428), .B(n9427), .Z(n9432) );
  NANDN U10023 ( .A(n9430), .B(n9429), .Z(n9431) );
  NAND U10024 ( .A(n9432), .B(n9431), .Z(n9857) );
  NANDN U10025 ( .A(n2978), .B(o[26]), .Z(n9853) );
  OR U10026 ( .A(n9434), .B(n9433), .Z(n9438) );
  OR U10027 ( .A(n9436), .B(n9435), .Z(n9437) );
  NAND U10028 ( .A(n9438), .B(n9437), .Z(n9851) );
  NANDN U10029 ( .A(n2980), .B(o[24]), .Z(n9711) );
  OR U10030 ( .A(n9439), .B(n16589), .Z(n9443) );
  NANDN U10031 ( .A(n9441), .B(n9440), .Z(n9442) );
  NAND U10032 ( .A(n9443), .B(n9442), .Z(n9709) );
  NANDN U10033 ( .A(n3016), .B(\stack[1][25] ), .Z(n9717) );
  NANDN U10034 ( .A(n9445), .B(n9444), .Z(n9449) );
  NANDN U10035 ( .A(n9447), .B(n9446), .Z(n9448) );
  AND U10036 ( .A(n9449), .B(n9448), .Z(n9714) );
  AND U10037 ( .A(\stack[1][26] ), .B(o[21]), .Z(n9720) );
  OR U10038 ( .A(n9451), .B(n9450), .Z(n9455) );
  OR U10039 ( .A(n9453), .B(n9452), .Z(n9454) );
  NAND U10040 ( .A(n9455), .B(n9454), .Z(n9721) );
  XNOR U10041 ( .A(n9720), .B(n9721), .Z(n9723) );
  NANDN U10042 ( .A(n9457), .B(n9456), .Z(n9461) );
  OR U10043 ( .A(n9459), .B(n9458), .Z(n9460) );
  NAND U10044 ( .A(n9461), .B(n9460), .Z(n9727) );
  ANDN U10045 ( .B(o[19]), .A(n2985), .Z(n9726) );
  XNOR U10046 ( .A(n9727), .B(n9726), .Z(n9728) );
  NANDN U10047 ( .A(n3012), .B(\stack[1][29] ), .Z(n9835) );
  NANDN U10048 ( .A(n9463), .B(n9462), .Z(n9467) );
  NANDN U10049 ( .A(n9465), .B(n9464), .Z(n9466) );
  AND U10050 ( .A(n9467), .B(n9466), .Z(n9832) );
  AND U10051 ( .A(\stack[1][30] ), .B(o[17]), .Z(n9732) );
  OR U10052 ( .A(n9469), .B(n9468), .Z(n9473) );
  OR U10053 ( .A(n9471), .B(n9470), .Z(n9472) );
  NAND U10054 ( .A(n9473), .B(n9472), .Z(n9733) );
  XNOR U10055 ( .A(n9732), .B(n9733), .Z(n9735) );
  OR U10056 ( .A(n9475), .B(n9474), .Z(n9479) );
  NANDN U10057 ( .A(n9477), .B(n9476), .Z(n9478) );
  NAND U10058 ( .A(n9479), .B(n9478), .Z(n9827) );
  ANDN U10059 ( .B(o[15]), .A(n2989), .Z(n9826) );
  XOR U10060 ( .A(n9827), .B(n9826), .Z(n9828) );
  NANDN U10061 ( .A(n3008), .B(\stack[1][33] ), .Z(n9823) );
  OR U10062 ( .A(n9481), .B(n9480), .Z(n9485) );
  NANDN U10063 ( .A(n9483), .B(n9482), .Z(n9484) );
  NAND U10064 ( .A(n9485), .B(n9484), .Z(n9821) );
  AND U10065 ( .A(\stack[1][34] ), .B(o[13]), .Z(n9744) );
  OR U10066 ( .A(n9487), .B(n9486), .Z(n9491) );
  OR U10067 ( .A(n9489), .B(n9488), .Z(n9490) );
  NAND U10068 ( .A(n9491), .B(n9490), .Z(n9745) );
  XNOR U10069 ( .A(n9744), .B(n9745), .Z(n9747) );
  NANDN U10070 ( .A(n9493), .B(n9492), .Z(n9497) );
  NANDN U10071 ( .A(n9495), .B(n9494), .Z(n9496) );
  AND U10072 ( .A(n9497), .B(n9496), .Z(n9814) );
  OR U10073 ( .A(n9499), .B(n9498), .Z(n9503) );
  OR U10074 ( .A(n9501), .B(n9500), .Z(n9502) );
  NAND U10075 ( .A(n9503), .B(n9502), .Z(n9757) );
  ANDN U10076 ( .B(\stack[1][38] ), .A(n3003), .Z(n9765) );
  OR U10077 ( .A(n9505), .B(n9504), .Z(n9509) );
  NANDN U10078 ( .A(n9507), .B(n9506), .Z(n9508) );
  AND U10079 ( .A(n9509), .B(n9508), .Z(n9762) );
  NANDN U10080 ( .A(n9511), .B(n9510), .Z(n9515) );
  NAND U10081 ( .A(n9513), .B(n9512), .Z(n9514) );
  AND U10082 ( .A(n9515), .B(n9514), .Z(n9805) );
  AND U10083 ( .A(\stack[1][42] ), .B(o[5]), .Z(n9799) );
  OR U10084 ( .A(n9517), .B(n9516), .Z(n9521) );
  NANDN U10085 ( .A(n9519), .B(n9518), .Z(n9520) );
  AND U10086 ( .A(n9521), .B(n9520), .Z(n9796) );
  AND U10087 ( .A(\stack[1][43] ), .B(o[4]), .Z(n9777) );
  AND U10088 ( .A(\stack[1][44] ), .B(o[3]), .Z(n9793) );
  NANDN U10089 ( .A(n9522), .B(n9780), .Z(n9523) );
  AND U10090 ( .A(n9524), .B(n9523), .Z(n9528) );
  OR U10091 ( .A(n9526), .B(n9525), .Z(n9527) );
  AND U10092 ( .A(n9528), .B(n9527), .Z(n9790) );
  AND U10093 ( .A(\stack[1][47] ), .B(o[1]), .Z(n9788) );
  ANDN U10094 ( .B(n9788), .A(n9529), .Z(n10054) );
  XNOR U10095 ( .A(n10054), .B(n9780), .Z(n9531) );
  NAND U10096 ( .A(\stack[1][47] ), .B(o[0]), .Z(n9787) );
  NANDN U10097 ( .A(n9530), .B(n9787), .Z(n9782) );
  NAND U10098 ( .A(n9531), .B(n9782), .Z(n9784) );
  AND U10099 ( .A(\stack[1][45] ), .B(o[2]), .Z(n9783) );
  XNOR U10100 ( .A(n9784), .B(n9783), .Z(n9791) );
  XOR U10101 ( .A(n9790), .B(n9791), .Z(n9792) );
  XOR U10102 ( .A(n9793), .B(n9792), .Z(n9775) );
  OR U10103 ( .A(n9533), .B(n9532), .Z(n9537) );
  NANDN U10104 ( .A(n9535), .B(n9534), .Z(n9536) );
  AND U10105 ( .A(n9537), .B(n9536), .Z(n9774) );
  XOR U10106 ( .A(n9775), .B(n9774), .Z(n9776) );
  XOR U10107 ( .A(n9777), .B(n9776), .Z(n9797) );
  XNOR U10108 ( .A(n9796), .B(n9797), .Z(n9798) );
  OR U10109 ( .A(n9539), .B(n9538), .Z(n9543) );
  OR U10110 ( .A(n9541), .B(n9540), .Z(n9542) );
  NAND U10111 ( .A(n9543), .B(n9542), .Z(n9769) );
  IV U10112 ( .A(\stack[1][41] ), .Z(n15896) );
  ANDN U10113 ( .B(o[6]), .A(n15896), .Z(n9768) );
  XNOR U10114 ( .A(n9769), .B(n9768), .Z(n9771) );
  XNOR U10115 ( .A(n9770), .B(n9771), .Z(n9803) );
  ANDN U10116 ( .B(o[7]), .A(n15935), .Z(n9802) );
  XOR U10117 ( .A(n9803), .B(n9802), .Z(n9804) );
  NANDN U10118 ( .A(n9545), .B(n9544), .Z(n9549) );
  NANDN U10119 ( .A(n9547), .B(n9546), .Z(n9548) );
  AND U10120 ( .A(n9549), .B(n9548), .Z(n9808) );
  XNOR U10121 ( .A(n9809), .B(n9808), .Z(n9811) );
  NANDN U10122 ( .A(n3002), .B(\stack[1][39] ), .Z(n9810) );
  XOR U10123 ( .A(n9811), .B(n9810), .Z(n9763) );
  XNOR U10124 ( .A(n9762), .B(n9763), .Z(n9764) );
  XOR U10125 ( .A(n9757), .B(n9756), .Z(n9759) );
  AND U10126 ( .A(\stack[1][37] ), .B(o[10]), .Z(n9758) );
  XNOR U10127 ( .A(n9759), .B(n9758), .Z(n9752) );
  AND U10128 ( .A(\stack[1][36] ), .B(o[11]), .Z(n9750) );
  OR U10129 ( .A(n9551), .B(n9550), .Z(n9555) );
  OR U10130 ( .A(n9553), .B(n9552), .Z(n9554) );
  NAND U10131 ( .A(n9555), .B(n9554), .Z(n9751) );
  XNOR U10132 ( .A(n9750), .B(n9751), .Z(n9753) );
  XNOR U10133 ( .A(n9752), .B(n9753), .Z(n9815) );
  XNOR U10134 ( .A(n9814), .B(n9815), .Z(n9816) );
  AND U10135 ( .A(\stack[1][35] ), .B(o[12]), .Z(n9817) );
  XOR U10136 ( .A(n9747), .B(n9746), .Z(n9820) );
  XNOR U10137 ( .A(n9821), .B(n9820), .Z(n9822) );
  XNOR U10138 ( .A(n9823), .B(n9822), .Z(n9829) );
  OR U10139 ( .A(n9557), .B(n9556), .Z(n9561) );
  OR U10140 ( .A(n9559), .B(n9558), .Z(n9560) );
  AND U10141 ( .A(n9561), .B(n9560), .Z(n9739) );
  XNOR U10142 ( .A(n9738), .B(n9739), .Z(n9741) );
  AND U10143 ( .A(\stack[1][31] ), .B(o[16]), .Z(n9740) );
  XNOR U10144 ( .A(n9741), .B(n9740), .Z(n9734) );
  XOR U10145 ( .A(n9735), .B(n9734), .Z(n9833) );
  XNOR U10146 ( .A(n9832), .B(n9833), .Z(n9834) );
  XOR U10147 ( .A(n9728), .B(n9729), .Z(n9838) );
  OR U10148 ( .A(n9563), .B(n9562), .Z(n9567) );
  OR U10149 ( .A(n9565), .B(n9564), .Z(n9566) );
  AND U10150 ( .A(n9567), .B(n9566), .Z(n9839) );
  XOR U10151 ( .A(n9838), .B(n9839), .Z(n9841) );
  AND U10152 ( .A(\stack[1][27] ), .B(o[20]), .Z(n9840) );
  XNOR U10153 ( .A(n9841), .B(n9840), .Z(n9722) );
  XNOR U10154 ( .A(n9714), .B(n9715), .Z(n9716) );
  XNOR U10155 ( .A(n9717), .B(n9716), .Z(n9846) );
  NANDN U10156 ( .A(n9569), .B(n9568), .Z(n9573) );
  OR U10157 ( .A(n9571), .B(n9570), .Z(n9572) );
  AND U10158 ( .A(n9573), .B(n9572), .Z(n9845) );
  NANDN U10159 ( .A(n2981), .B(o[23]), .Z(n9844) );
  XOR U10160 ( .A(n9845), .B(n9844), .Z(n9847) );
  XNOR U10161 ( .A(n9846), .B(n9847), .Z(n9708) );
  XNOR U10162 ( .A(n9709), .B(n9708), .Z(n9710) );
  XNOR U10163 ( .A(n9711), .B(n9710), .Z(n9704) );
  OR U10164 ( .A(n9575), .B(n9574), .Z(n9579) );
  NANDN U10165 ( .A(n9577), .B(n9576), .Z(n9578) );
  AND U10166 ( .A(n9579), .B(n9578), .Z(n9703) );
  NANDN U10167 ( .A(n3019), .B(\stack[1][22] ), .Z(n9702) );
  XOR U10168 ( .A(n9703), .B(n9702), .Z(n9705) );
  XNOR U10169 ( .A(n9704), .B(n9705), .Z(n9850) );
  XNOR U10170 ( .A(n9851), .B(n9850), .Z(n9852) );
  XNOR U10171 ( .A(n9853), .B(n9852), .Z(n9698) );
  NANDN U10172 ( .A(n16712), .B(o[27]), .Z(n9696) );
  OR U10173 ( .A(n9581), .B(n9580), .Z(n9585) );
  OR U10174 ( .A(n9583), .B(n9582), .Z(n9584) );
  NAND U10175 ( .A(n9585), .B(n9584), .Z(n9697) );
  XOR U10176 ( .A(n9696), .B(n9697), .Z(n9699) );
  XNOR U10177 ( .A(n9698), .B(n9699), .Z(n9856) );
  XNOR U10178 ( .A(n9857), .B(n9856), .Z(n9858) );
  XNOR U10179 ( .A(n9859), .B(n9858), .Z(n9692) );
  NANDN U10180 ( .A(n16786), .B(o[29]), .Z(n9690) );
  OR U10181 ( .A(n9587), .B(n9586), .Z(n9591) );
  OR U10182 ( .A(n9589), .B(n9588), .Z(n9590) );
  NAND U10183 ( .A(n9591), .B(n9590), .Z(n9691) );
  XOR U10184 ( .A(n9690), .B(n9691), .Z(n9693) );
  XNOR U10185 ( .A(n9692), .B(n9693), .Z(n9862) );
  XNOR U10186 ( .A(n9863), .B(n9862), .Z(n9864) );
  XNOR U10187 ( .A(n9865), .B(n9864), .Z(n9686) );
  NANDN U10188 ( .A(n2977), .B(o[31]), .Z(n9684) );
  OR U10189 ( .A(n9593), .B(n9592), .Z(n9597) );
  OR U10190 ( .A(n9595), .B(n9594), .Z(n9596) );
  NAND U10191 ( .A(n9597), .B(n9596), .Z(n9685) );
  XOR U10192 ( .A(n9684), .B(n9685), .Z(n9687) );
  XNOR U10193 ( .A(n9686), .B(n9687), .Z(n9869) );
  XNOR U10194 ( .A(n9868), .B(n9869), .Z(n9870) );
  XOR U10195 ( .A(n9680), .B(n9681), .Z(n9672) );
  OR U10196 ( .A(n9599), .B(n9598), .Z(n9603) );
  NANDN U10197 ( .A(n9601), .B(n9600), .Z(n9602) );
  AND U10198 ( .A(n9603), .B(n9602), .Z(n9673) );
  XOR U10199 ( .A(n9672), .B(n9673), .Z(n9675) );
  AND U10200 ( .A(o[34]), .B(\stack[1][13] ), .Z(n9674) );
  XOR U10201 ( .A(n9675), .B(n9674), .Z(n9876) );
  XOR U10202 ( .A(n9877), .B(n9876), .Z(n9667) );
  XOR U10203 ( .A(n9666), .B(n9667), .Z(n9668) );
  XOR U10204 ( .A(n9669), .B(n9668), .Z(n9663) );
  AND U10205 ( .A(o[37]), .B(\stack[1][10] ), .Z(n9660) );
  OR U10206 ( .A(n9605), .B(n9604), .Z(n9609) );
  OR U10207 ( .A(n9607), .B(n9606), .Z(n9608) );
  NAND U10208 ( .A(n9609), .B(n9608), .Z(n9661) );
  XNOR U10209 ( .A(n9660), .B(n9661), .Z(n9662) );
  XOR U10210 ( .A(n9663), .B(n9662), .Z(n9880) );
  XNOR U10211 ( .A(n9881), .B(n9880), .Z(n9882) );
  XNOR U10212 ( .A(n9883), .B(n9882), .Z(n9656) );
  NANDN U10213 ( .A(n17179), .B(o[39]), .Z(n9654) );
  OR U10214 ( .A(n9611), .B(n9610), .Z(n9615) );
  OR U10215 ( .A(n9613), .B(n9612), .Z(n9614) );
  NAND U10216 ( .A(n9615), .B(n9614), .Z(n9655) );
  XOR U10217 ( .A(n9654), .B(n9655), .Z(n9657) );
  XNOR U10218 ( .A(n9656), .B(n9657), .Z(n9886) );
  XNOR U10219 ( .A(n9887), .B(n9886), .Z(n9888) );
  XNOR U10220 ( .A(n9889), .B(n9888), .Z(n9650) );
  NANDN U10221 ( .A(n17256), .B(o[41]), .Z(n9648) );
  OR U10222 ( .A(n9617), .B(n9616), .Z(n9621) );
  OR U10223 ( .A(n9619), .B(n9618), .Z(n9620) );
  NAND U10224 ( .A(n9621), .B(n9620), .Z(n9649) );
  XOR U10225 ( .A(n9648), .B(n9649), .Z(n9651) );
  XNOR U10226 ( .A(n9650), .B(n9651), .Z(n9892) );
  XNOR U10227 ( .A(n9893), .B(n9892), .Z(n9894) );
  XNOR U10228 ( .A(n9895), .B(n9894), .Z(n9644) );
  AND U10229 ( .A(o[43]), .B(\stack[1][4] ), .Z(n9642) );
  OR U10230 ( .A(n9623), .B(n9622), .Z(n9627) );
  OR U10231 ( .A(n9625), .B(n9624), .Z(n9626) );
  NAND U10232 ( .A(n9627), .B(n9626), .Z(n9643) );
  XNOR U10233 ( .A(n9642), .B(n9643), .Z(n9645) );
  XNOR U10234 ( .A(n9644), .B(n9645), .Z(n9898) );
  XNOR U10235 ( .A(n9899), .B(n9898), .Z(n9900) );
  XOR U10236 ( .A(n9901), .B(n9900), .Z(n9639) );
  AND U10237 ( .A(o[45]), .B(\stack[1][2] ), .Z(n9636) );
  OR U10238 ( .A(n9629), .B(n9628), .Z(n9633) );
  OR U10239 ( .A(n9631), .B(n9630), .Z(n9632) );
  NAND U10240 ( .A(n9633), .B(n9632), .Z(n9637) );
  XOR U10241 ( .A(n9636), .B(n9637), .Z(n9638) );
  XNOR U10242 ( .A(n9639), .B(n9638), .Z(n9904) );
  XNOR U10243 ( .A(n9905), .B(n9904), .Z(n9906) );
  XOR U10244 ( .A(n9907), .B(n9906), .Z(n15666) );
  OR U10245 ( .A(n15665), .B(n15666), .Z(n9634) );
  AND U10246 ( .A(n9635), .B(n9634), .Z(n9911) );
  NANDN U10247 ( .A(n2970), .B(o[46]), .Z(n10192) );
  OR U10248 ( .A(n9637), .B(n9636), .Z(n9641) );
  NANDN U10249 ( .A(n9639), .B(n9638), .Z(n9640) );
  NAND U10250 ( .A(n9641), .B(n9640), .Z(n10190) );
  NANDN U10251 ( .A(n2971), .B(o[44]), .Z(n10186) );
  OR U10252 ( .A(n9643), .B(n9642), .Z(n9647) );
  NANDN U10253 ( .A(n9645), .B(n9644), .Z(n9646) );
  NAND U10254 ( .A(n9647), .B(n9646), .Z(n10184) );
  NANDN U10255 ( .A(n17256), .B(o[42]), .Z(n10180) );
  NANDN U10256 ( .A(n9649), .B(n9648), .Z(n9653) );
  NANDN U10257 ( .A(n9651), .B(n9650), .Z(n9652) );
  NAND U10258 ( .A(n9653), .B(n9652), .Z(n10178) );
  NANDN U10259 ( .A(n17179), .B(o[40]), .Z(n10174) );
  NANDN U10260 ( .A(n9655), .B(n9654), .Z(n9659) );
  NANDN U10261 ( .A(n9657), .B(n9656), .Z(n9658) );
  NAND U10262 ( .A(n9659), .B(n9658), .Z(n10172) );
  AND U10263 ( .A(o[38]), .B(\stack[1][10] ), .Z(n9949) );
  OR U10264 ( .A(n9661), .B(n9660), .Z(n9665) );
  OR U10265 ( .A(n9663), .B(n9662), .Z(n9664) );
  AND U10266 ( .A(n9665), .B(n9664), .Z(n9946) );
  OR U10267 ( .A(n9667), .B(n9666), .Z(n9671) );
  NANDN U10268 ( .A(n9669), .B(n9668), .Z(n9670) );
  AND U10269 ( .A(n9671), .B(n9670), .Z(n10165) );
  AND U10270 ( .A(o[37]), .B(\stack[1][11] ), .Z(n10166) );
  XNOR U10271 ( .A(n10165), .B(n10166), .Z(n10168) );
  NANDN U10272 ( .A(n9673), .B(n9672), .Z(n9677) );
  OR U10273 ( .A(n9675), .B(n9674), .Z(n9676) );
  NAND U10274 ( .A(n9677), .B(n9676), .Z(n9959) );
  ANDN U10275 ( .B(o[35]), .A(n2974), .Z(n9958) );
  XNOR U10276 ( .A(n9959), .B(n9958), .Z(n9960) );
  NANDN U10277 ( .A(n2975), .B(o[34]), .Z(n10162) );
  NANDN U10278 ( .A(n9679), .B(n9678), .Z(n9683) );
  NANDN U10279 ( .A(n9681), .B(n9680), .Z(n9682) );
  AND U10280 ( .A(n9683), .B(n9682), .Z(n10159) );
  NANDN U10281 ( .A(n2977), .B(o[32]), .Z(n10156) );
  NANDN U10282 ( .A(n9685), .B(n9684), .Z(n9689) );
  NANDN U10283 ( .A(n9687), .B(n9686), .Z(n9688) );
  NAND U10284 ( .A(n9689), .B(n9688), .Z(n10154) );
  NANDN U10285 ( .A(n16786), .B(o[30]), .Z(n10150) );
  NANDN U10286 ( .A(n9691), .B(n9690), .Z(n9695) );
  NANDN U10287 ( .A(n9693), .B(n9692), .Z(n9694) );
  NAND U10288 ( .A(n9695), .B(n9694), .Z(n10148) );
  NANDN U10289 ( .A(n16712), .B(o[28]), .Z(n10144) );
  NANDN U10290 ( .A(n9697), .B(n9696), .Z(n9701) );
  NANDN U10291 ( .A(n9699), .B(n9698), .Z(n9700) );
  NAND U10292 ( .A(n9701), .B(n9700), .Z(n10142) );
  NANDN U10293 ( .A(n2979), .B(o[26]), .Z(n10138) );
  NANDN U10294 ( .A(n9703), .B(n9702), .Z(n9707) );
  NANDN U10295 ( .A(n9705), .B(n9704), .Z(n9706) );
  NAND U10296 ( .A(n9707), .B(n9706), .Z(n10136) );
  AND U10297 ( .A(o[25]), .B(\stack[1][23] ), .Z(n9988) );
  OR U10298 ( .A(n9709), .B(n9708), .Z(n9713) );
  OR U10299 ( .A(n9711), .B(n9710), .Z(n9712) );
  NAND U10300 ( .A(n9713), .B(n9712), .Z(n9989) );
  XNOR U10301 ( .A(n9988), .B(n9989), .Z(n9991) );
  AND U10302 ( .A(o[24]), .B(\stack[1][24] ), .Z(n16555) );
  NANDN U10303 ( .A(n3017), .B(\stack[1][25] ), .Z(n9995) );
  OR U10304 ( .A(n9715), .B(n9714), .Z(n9719) );
  OR U10305 ( .A(n9717), .B(n9716), .Z(n9718) );
  AND U10306 ( .A(n9719), .B(n9718), .Z(n9994) );
  XNOR U10307 ( .A(n9995), .B(n9994), .Z(n9996) );
  OR U10308 ( .A(n9721), .B(n9720), .Z(n9725) );
  OR U10309 ( .A(n9723), .B(n9722), .Z(n9724) );
  NAND U10310 ( .A(n9725), .B(n9724), .Z(n10125) );
  NANDN U10311 ( .A(n3014), .B(\stack[1][28] ), .Z(n10121) );
  NANDN U10312 ( .A(n9727), .B(n9726), .Z(n9731) );
  NANDN U10313 ( .A(n9729), .B(n9728), .Z(n9730) );
  AND U10314 ( .A(n9731), .B(n9730), .Z(n10118) );
  NANDN U10315 ( .A(n3012), .B(\stack[1][30] ), .Z(n10115) );
  OR U10316 ( .A(n9733), .B(n9732), .Z(n9737) );
  OR U10317 ( .A(n9735), .B(n9734), .Z(n9736) );
  NAND U10318 ( .A(n9737), .B(n9736), .Z(n10113) );
  OR U10319 ( .A(n9739), .B(n9738), .Z(n9743) );
  OR U10320 ( .A(n9741), .B(n9740), .Z(n9742) );
  AND U10321 ( .A(n9743), .B(n9742), .Z(n10012) );
  AND U10322 ( .A(\stack[1][31] ), .B(o[17]), .Z(n10013) );
  XNOR U10323 ( .A(n10012), .B(n10013), .Z(n10015) );
  OR U10324 ( .A(n9745), .B(n9744), .Z(n9749) );
  OR U10325 ( .A(n9747), .B(n9746), .Z(n9748) );
  NAND U10326 ( .A(n9749), .B(n9748), .Z(n10107) );
  AND U10327 ( .A(\stack[1][36] ), .B(o[12]), .Z(n10103) );
  OR U10328 ( .A(n9751), .B(n9750), .Z(n9755) );
  OR U10329 ( .A(n9753), .B(n9752), .Z(n9754) );
  AND U10330 ( .A(n9755), .B(n9754), .Z(n10100) );
  AND U10331 ( .A(\stack[1][37] ), .B(o[11]), .Z(n10094) );
  NANDN U10332 ( .A(n9757), .B(n9756), .Z(n9761) );
  NANDN U10333 ( .A(n9759), .B(n9758), .Z(n9760) );
  NAND U10334 ( .A(n9761), .B(n9760), .Z(n10095) );
  XNOR U10335 ( .A(n10094), .B(n10095), .Z(n10097) );
  NANDN U10336 ( .A(n3004), .B(\stack[1][38] ), .Z(n10038) );
  OR U10337 ( .A(n9763), .B(n9762), .Z(n9767) );
  OR U10338 ( .A(n9765), .B(n9764), .Z(n9766) );
  AND U10339 ( .A(n9767), .B(n9766), .Z(n10037) );
  NANDN U10340 ( .A(n3003), .B(\stack[1][39] ), .Z(n10090) );
  NANDN U10341 ( .A(n9769), .B(n9768), .Z(n9773) );
  NAND U10342 ( .A(n9771), .B(n9770), .Z(n9772) );
  AND U10343 ( .A(n9773), .B(n9772), .Z(n10079) );
  AND U10344 ( .A(\stack[1][43] ), .B(o[5]), .Z(n10073) );
  OR U10345 ( .A(n9775), .B(n9774), .Z(n9779) );
  NANDN U10346 ( .A(n9777), .B(n9776), .Z(n9778) );
  AND U10347 ( .A(n9779), .B(n9778), .Z(n10070) );
  AND U10348 ( .A(\stack[1][44] ), .B(o[4]), .Z(n10051) );
  AND U10349 ( .A(\stack[1][45] ), .B(o[3]), .Z(n10067) );
  NANDN U10350 ( .A(n9780), .B(n10054), .Z(n9781) );
  AND U10351 ( .A(n9782), .B(n9781), .Z(n9786) );
  OR U10352 ( .A(n9784), .B(n9783), .Z(n9785) );
  AND U10353 ( .A(n9786), .B(n9785), .Z(n10064) );
  AND U10354 ( .A(\stack[1][48] ), .B(o[1]), .Z(n10062) );
  ANDN U10355 ( .B(n10062), .A(n9787), .Z(n10335) );
  XNOR U10356 ( .A(n10335), .B(n10054), .Z(n9789) );
  NAND U10357 ( .A(\stack[1][48] ), .B(o[0]), .Z(n10061) );
  NANDN U10358 ( .A(n9788), .B(n10061), .Z(n10056) );
  NAND U10359 ( .A(n9789), .B(n10056), .Z(n10058) );
  AND U10360 ( .A(\stack[1][46] ), .B(o[2]), .Z(n10057) );
  XNOR U10361 ( .A(n10058), .B(n10057), .Z(n10065) );
  XOR U10362 ( .A(n10064), .B(n10065), .Z(n10066) );
  XOR U10363 ( .A(n10067), .B(n10066), .Z(n10049) );
  OR U10364 ( .A(n9791), .B(n9790), .Z(n9795) );
  NANDN U10365 ( .A(n9793), .B(n9792), .Z(n9794) );
  AND U10366 ( .A(n9795), .B(n9794), .Z(n10048) );
  XOR U10367 ( .A(n10049), .B(n10048), .Z(n10050) );
  XOR U10368 ( .A(n10051), .B(n10050), .Z(n10071) );
  XNOR U10369 ( .A(n10070), .B(n10071), .Z(n10072) );
  OR U10370 ( .A(n9797), .B(n9796), .Z(n9801) );
  OR U10371 ( .A(n9799), .B(n9798), .Z(n9800) );
  NAND U10372 ( .A(n9801), .B(n9800), .Z(n10043) );
  IV U10373 ( .A(\stack[1][42] ), .Z(n15857) );
  ANDN U10374 ( .B(o[6]), .A(n15857), .Z(n10042) );
  XNOR U10375 ( .A(n10043), .B(n10042), .Z(n10045) );
  XNOR U10376 ( .A(n10044), .B(n10045), .Z(n10077) );
  ANDN U10377 ( .B(o[7]), .A(n15896), .Z(n10076) );
  XOR U10378 ( .A(n10077), .B(n10076), .Z(n10078) );
  NANDN U10379 ( .A(n9803), .B(n9802), .Z(n9807) );
  OR U10380 ( .A(n9805), .B(n9804), .Z(n9806) );
  AND U10381 ( .A(n9807), .B(n9806), .Z(n10082) );
  XNOR U10382 ( .A(n10083), .B(n10082), .Z(n10085) );
  ANDN U10383 ( .B(o[8]), .A(n15935), .Z(n10084) );
  XOR U10384 ( .A(n10085), .B(n10084), .Z(n10088) );
  OR U10385 ( .A(n9809), .B(n9808), .Z(n9813) );
  OR U10386 ( .A(n9811), .B(n9810), .Z(n9812) );
  NAND U10387 ( .A(n9813), .B(n9812), .Z(n10089) );
  XOR U10388 ( .A(n10088), .B(n10089), .Z(n10091) );
  XNOR U10389 ( .A(n10090), .B(n10091), .Z(n10036) );
  XOR U10390 ( .A(n10037), .B(n10036), .Z(n10039) );
  XNOR U10391 ( .A(n10038), .B(n10039), .Z(n10096) );
  XOR U10392 ( .A(n10097), .B(n10096), .Z(n10101) );
  XOR U10393 ( .A(n10100), .B(n10101), .Z(n10102) );
  XOR U10394 ( .A(n10103), .B(n10102), .Z(n10033) );
  OR U10395 ( .A(n9815), .B(n9814), .Z(n9819) );
  OR U10396 ( .A(n9817), .B(n9816), .Z(n9818) );
  AND U10397 ( .A(n9819), .B(n9818), .Z(n10031) );
  NANDN U10398 ( .A(n2992), .B(o[13]), .Z(n10030) );
  XOR U10399 ( .A(n10031), .B(n10030), .Z(n10032) );
  XNOR U10400 ( .A(n10033), .B(n10032), .Z(n10106) );
  XOR U10401 ( .A(n10107), .B(n10106), .Z(n10109) );
  AND U10402 ( .A(\stack[1][34] ), .B(o[14]), .Z(n10108) );
  XNOR U10403 ( .A(n10109), .B(n10108), .Z(n10026) );
  AND U10404 ( .A(\stack[1][33] ), .B(o[15]), .Z(n10024) );
  OR U10405 ( .A(n9821), .B(n9820), .Z(n9825) );
  OR U10406 ( .A(n9823), .B(n9822), .Z(n9824) );
  NAND U10407 ( .A(n9825), .B(n9824), .Z(n10025) );
  XNOR U10408 ( .A(n10024), .B(n10025), .Z(n10027) );
  XNOR U10409 ( .A(n10026), .B(n10027), .Z(n10019) );
  NANDN U10410 ( .A(n9827), .B(n9826), .Z(n9831) );
  OR U10411 ( .A(n9829), .B(n9828), .Z(n9830) );
  NAND U10412 ( .A(n9831), .B(n9830), .Z(n10018) );
  XOR U10413 ( .A(n10019), .B(n10018), .Z(n10020) );
  AND U10414 ( .A(\stack[1][32] ), .B(o[16]), .Z(n10021) );
  XOR U10415 ( .A(n10020), .B(n10021), .Z(n10014) );
  XOR U10416 ( .A(n10015), .B(n10014), .Z(n10112) );
  XNOR U10417 ( .A(n10113), .B(n10112), .Z(n10114) );
  XOR U10418 ( .A(n10115), .B(n10114), .Z(n10008) );
  AND U10419 ( .A(\stack[1][29] ), .B(o[19]), .Z(n10006) );
  OR U10420 ( .A(n9833), .B(n9832), .Z(n9837) );
  OR U10421 ( .A(n9835), .B(n9834), .Z(n9836) );
  NAND U10422 ( .A(n9837), .B(n9836), .Z(n10007) );
  XNOR U10423 ( .A(n10006), .B(n10007), .Z(n10009) );
  XNOR U10424 ( .A(n10118), .B(n10119), .Z(n10120) );
  XOR U10425 ( .A(n10121), .B(n10120), .Z(n10002) );
  NANDN U10426 ( .A(n9839), .B(n9838), .Z(n9843) );
  OR U10427 ( .A(n9841), .B(n9840), .Z(n9842) );
  AND U10428 ( .A(n9843), .B(n9842), .Z(n10000) );
  AND U10429 ( .A(\stack[1][27] ), .B(o[21]), .Z(n10001) );
  XNOR U10430 ( .A(n10000), .B(n10001), .Z(n10003) );
  XOR U10431 ( .A(n10125), .B(n10124), .Z(n10127) );
  NANDN U10432 ( .A(n3016), .B(\stack[1][26] ), .Z(n10126) );
  XNOR U10433 ( .A(n10127), .B(n10126), .Z(n9997) );
  NANDN U10434 ( .A(n9845), .B(n9844), .Z(n9849) );
  NANDN U10435 ( .A(n9847), .B(n9846), .Z(n9848) );
  AND U10436 ( .A(n9849), .B(n9848), .Z(n10131) );
  XNOR U10437 ( .A(n10130), .B(n10131), .Z(n10132) );
  XNOR U10438 ( .A(n16555), .B(n10132), .Z(n9990) );
  XOR U10439 ( .A(n9991), .B(n9990), .Z(n10135) );
  XNOR U10440 ( .A(n10136), .B(n10135), .Z(n10137) );
  XNOR U10441 ( .A(n10138), .B(n10137), .Z(n9984) );
  NANDN U10442 ( .A(n2978), .B(o[27]), .Z(n9982) );
  OR U10443 ( .A(n9851), .B(n9850), .Z(n9855) );
  OR U10444 ( .A(n9853), .B(n9852), .Z(n9854) );
  NAND U10445 ( .A(n9855), .B(n9854), .Z(n9983) );
  XOR U10446 ( .A(n9982), .B(n9983), .Z(n9985) );
  XNOR U10447 ( .A(n9984), .B(n9985), .Z(n10141) );
  XNOR U10448 ( .A(n10142), .B(n10141), .Z(n10143) );
  XNOR U10449 ( .A(n10144), .B(n10143), .Z(n9978) );
  NANDN U10450 ( .A(n16746), .B(o[29]), .Z(n9976) );
  OR U10451 ( .A(n9857), .B(n9856), .Z(n9861) );
  OR U10452 ( .A(n9859), .B(n9858), .Z(n9860) );
  NAND U10453 ( .A(n9861), .B(n9860), .Z(n9977) );
  XOR U10454 ( .A(n9976), .B(n9977), .Z(n9979) );
  XNOR U10455 ( .A(n9978), .B(n9979), .Z(n10147) );
  XNOR U10456 ( .A(n10148), .B(n10147), .Z(n10149) );
  XNOR U10457 ( .A(n10150), .B(n10149), .Z(n9972) );
  NANDN U10458 ( .A(n16826), .B(o[31]), .Z(n9970) );
  OR U10459 ( .A(n9863), .B(n9862), .Z(n9867) );
  OR U10460 ( .A(n9865), .B(n9864), .Z(n9866) );
  NAND U10461 ( .A(n9867), .B(n9866), .Z(n9971) );
  XOR U10462 ( .A(n9970), .B(n9971), .Z(n9973) );
  XNOR U10463 ( .A(n9972), .B(n9973), .Z(n10153) );
  XNOR U10464 ( .A(n10154), .B(n10153), .Z(n10155) );
  XNOR U10465 ( .A(n10156), .B(n10155), .Z(n9966) );
  NANDN U10466 ( .A(n2976), .B(o[33]), .Z(n9964) );
  OR U10467 ( .A(n9869), .B(n9868), .Z(n9873) );
  OR U10468 ( .A(n9871), .B(n9870), .Z(n9872) );
  NAND U10469 ( .A(n9873), .B(n9872), .Z(n9965) );
  XOR U10470 ( .A(n9964), .B(n9965), .Z(n9967) );
  XNOR U10471 ( .A(n9966), .B(n9967), .Z(n10160) );
  XNOR U10472 ( .A(n10159), .B(n10160), .Z(n10161) );
  XOR U10473 ( .A(n9960), .B(n9961), .Z(n9952) );
  OR U10474 ( .A(n9875), .B(n9874), .Z(n9879) );
  NANDN U10475 ( .A(n9877), .B(n9876), .Z(n9878) );
  AND U10476 ( .A(n9879), .B(n9878), .Z(n9953) );
  XOR U10477 ( .A(n9952), .B(n9953), .Z(n9955) );
  AND U10478 ( .A(o[36]), .B(\stack[1][12] ), .Z(n9954) );
  XOR U10479 ( .A(n9955), .B(n9954), .Z(n10167) );
  XOR U10480 ( .A(n10168), .B(n10167), .Z(n9947) );
  XOR U10481 ( .A(n9946), .B(n9947), .Z(n9948) );
  XOR U10482 ( .A(n9949), .B(n9948), .Z(n9943) );
  AND U10483 ( .A(o[39]), .B(\stack[1][9] ), .Z(n9940) );
  OR U10484 ( .A(n9881), .B(n9880), .Z(n9885) );
  OR U10485 ( .A(n9883), .B(n9882), .Z(n9884) );
  NAND U10486 ( .A(n9885), .B(n9884), .Z(n9941) );
  XNOR U10487 ( .A(n9940), .B(n9941), .Z(n9942) );
  XOR U10488 ( .A(n9943), .B(n9942), .Z(n10171) );
  XNOR U10489 ( .A(n10172), .B(n10171), .Z(n10173) );
  XNOR U10490 ( .A(n10174), .B(n10173), .Z(n9936) );
  NANDN U10491 ( .A(n17219), .B(o[41]), .Z(n9934) );
  OR U10492 ( .A(n9887), .B(n9886), .Z(n9891) );
  OR U10493 ( .A(n9889), .B(n9888), .Z(n9890) );
  NAND U10494 ( .A(n9891), .B(n9890), .Z(n9935) );
  XOR U10495 ( .A(n9934), .B(n9935), .Z(n9937) );
  XNOR U10496 ( .A(n9936), .B(n9937), .Z(n10177) );
  XNOR U10497 ( .A(n10178), .B(n10177), .Z(n10179) );
  XNOR U10498 ( .A(n10180), .B(n10179), .Z(n9930) );
  NANDN U10499 ( .A(n17296), .B(o[43]), .Z(n9928) );
  OR U10500 ( .A(n9893), .B(n9892), .Z(n9897) );
  OR U10501 ( .A(n9895), .B(n9894), .Z(n9896) );
  NAND U10502 ( .A(n9897), .B(n9896), .Z(n9929) );
  XOR U10503 ( .A(n9928), .B(n9929), .Z(n9931) );
  XNOR U10504 ( .A(n9930), .B(n9931), .Z(n10183) );
  XNOR U10505 ( .A(n10184), .B(n10183), .Z(n10185) );
  XNOR U10506 ( .A(n10186), .B(n10185), .Z(n9924) );
  NANDN U10507 ( .A(n17375), .B(o[45]), .Z(n9922) );
  OR U10508 ( .A(n9899), .B(n9898), .Z(n9903) );
  OR U10509 ( .A(n9901), .B(n9900), .Z(n9902) );
  NAND U10510 ( .A(n9903), .B(n9902), .Z(n9923) );
  XOR U10511 ( .A(n9922), .B(n9923), .Z(n9925) );
  XNOR U10512 ( .A(n9924), .B(n9925), .Z(n10189) );
  XNOR U10513 ( .A(n10190), .B(n10189), .Z(n10191) );
  AND U10514 ( .A(o[47]), .B(\stack[1][1] ), .Z(n9916) );
  OR U10515 ( .A(n9905), .B(n9904), .Z(n9909) );
  OR U10516 ( .A(n9907), .B(n9906), .Z(n9908) );
  NAND U10517 ( .A(n9909), .B(n9908), .Z(n9917) );
  XNOR U10518 ( .A(n9916), .B(n9917), .Z(n9919) );
  XOR U10519 ( .A(n9918), .B(n9919), .Z(n9910) );
  NANDN U10520 ( .A(n9911), .B(n9910), .Z(n9913) );
  XOR U10521 ( .A(n9911), .B(n9910), .Z(n15626) );
  AND U10522 ( .A(o[48]), .B(\stack[1][0] ), .Z(n15627) );
  OR U10523 ( .A(n15626), .B(n15627), .Z(n9912) );
  AND U10524 ( .A(n9913), .B(n9912), .Z(n9915) );
  OR U10525 ( .A(n9914), .B(n9915), .Z(n10196) );
  XNOR U10526 ( .A(n9915), .B(n9914), .Z(n15587) );
  NANDN U10527 ( .A(n2969), .B(o[48]), .Z(n10480) );
  OR U10528 ( .A(n9917), .B(n9916), .Z(n9921) );
  OR U10529 ( .A(n9919), .B(n9918), .Z(n9920) );
  NAND U10530 ( .A(n9921), .B(n9920), .Z(n10478) );
  NANDN U10531 ( .A(n17375), .B(o[46]), .Z(n10474) );
  NANDN U10532 ( .A(n9923), .B(n9922), .Z(n9927) );
  NANDN U10533 ( .A(n9925), .B(n9924), .Z(n9926) );
  NAND U10534 ( .A(n9927), .B(n9926), .Z(n10472) );
  NANDN U10535 ( .A(n17296), .B(o[44]), .Z(n10468) );
  NANDN U10536 ( .A(n9929), .B(n9928), .Z(n9933) );
  NANDN U10537 ( .A(n9931), .B(n9930), .Z(n9932) );
  NAND U10538 ( .A(n9933), .B(n9932), .Z(n10466) );
  NANDN U10539 ( .A(n17219), .B(o[42]), .Z(n10462) );
  NANDN U10540 ( .A(n9935), .B(n9934), .Z(n9939) );
  NANDN U10541 ( .A(n9937), .B(n9936), .Z(n9938) );
  NAND U10542 ( .A(n9939), .B(n9938), .Z(n10460) );
  AND U10543 ( .A(o[40]), .B(\stack[1][9] ), .Z(n10456) );
  OR U10544 ( .A(n9941), .B(n9940), .Z(n9945) );
  OR U10545 ( .A(n9943), .B(n9942), .Z(n9944) );
  AND U10546 ( .A(n9945), .B(n9944), .Z(n10453) );
  OR U10547 ( .A(n9947), .B(n9946), .Z(n9951) );
  NANDN U10548 ( .A(n9949), .B(n9948), .Z(n9950) );
  AND U10549 ( .A(n9951), .B(n9950), .Z(n10221) );
  AND U10550 ( .A(o[39]), .B(\stack[1][10] ), .Z(n10222) );
  XNOR U10551 ( .A(n10221), .B(n10222), .Z(n10224) );
  NANDN U10552 ( .A(n9953), .B(n9952), .Z(n9957) );
  OR U10553 ( .A(n9955), .B(n9954), .Z(n9956) );
  NAND U10554 ( .A(n9957), .B(n9956), .Z(n10228) );
  ANDN U10555 ( .B(o[37]), .A(n2973), .Z(n10227) );
  XNOR U10556 ( .A(n10228), .B(n10227), .Z(n10229) );
  NANDN U10557 ( .A(n2974), .B(o[36]), .Z(n10444) );
  NANDN U10558 ( .A(n9959), .B(n9958), .Z(n9963) );
  NANDN U10559 ( .A(n9961), .B(n9960), .Z(n9962) );
  AND U10560 ( .A(n9963), .B(n9962), .Z(n10441) );
  NANDN U10561 ( .A(n2976), .B(o[34]), .Z(n10438) );
  NANDN U10562 ( .A(n9965), .B(n9964), .Z(n9969) );
  NANDN U10563 ( .A(n9967), .B(n9966), .Z(n9968) );
  NAND U10564 ( .A(n9969), .B(n9968), .Z(n10436) );
  NANDN U10565 ( .A(n16826), .B(o[32]), .Z(n10432) );
  NANDN U10566 ( .A(n9971), .B(n9970), .Z(n9975) );
  NANDN U10567 ( .A(n9973), .B(n9972), .Z(n9974) );
  NAND U10568 ( .A(n9975), .B(n9974), .Z(n10430) );
  NANDN U10569 ( .A(n16746), .B(o[30]), .Z(n10426) );
  NANDN U10570 ( .A(n9977), .B(n9976), .Z(n9981) );
  NANDN U10571 ( .A(n9979), .B(n9978), .Z(n9980) );
  NAND U10572 ( .A(n9981), .B(n9980), .Z(n10424) );
  NANDN U10573 ( .A(n2978), .B(o[28]), .Z(n10420) );
  NANDN U10574 ( .A(n9983), .B(n9982), .Z(n9987) );
  NANDN U10575 ( .A(n9985), .B(n9984), .Z(n9986) );
  NAND U10576 ( .A(n9987), .B(n9986), .Z(n10418) );
  NANDN U10577 ( .A(n2980), .B(o[26]), .Z(n10414) );
  OR U10578 ( .A(n9989), .B(n9988), .Z(n9993) );
  OR U10579 ( .A(n9991), .B(n9990), .Z(n9992) );
  NAND U10580 ( .A(n9993), .B(n9992), .Z(n10412) );
  NANDN U10581 ( .A(n3018), .B(\stack[1][25] ), .Z(n10408) );
  OR U10582 ( .A(n9995), .B(n9994), .Z(n9999) );
  OR U10583 ( .A(n9997), .B(n9996), .Z(n9998) );
  AND U10584 ( .A(n9999), .B(n9998), .Z(n10405) );
  NANDN U10585 ( .A(n3016), .B(\stack[1][27] ), .Z(n10402) );
  OR U10586 ( .A(n10001), .B(n10000), .Z(n10005) );
  OR U10587 ( .A(n10003), .B(n10002), .Z(n10004) );
  NAND U10588 ( .A(n10005), .B(n10004), .Z(n10400) );
  NANDN U10589 ( .A(n3014), .B(\stack[1][29] ), .Z(n10396) );
  OR U10590 ( .A(n10007), .B(n10006), .Z(n10011) );
  OR U10591 ( .A(n10009), .B(n10008), .Z(n10010) );
  NAND U10592 ( .A(n10011), .B(n10010), .Z(n10394) );
  NANDN U10593 ( .A(n3012), .B(\stack[1][31] ), .Z(n10290) );
  OR U10594 ( .A(n10013), .B(n10012), .Z(n10017) );
  OR U10595 ( .A(n10015), .B(n10014), .Z(n10016) );
  NAND U10596 ( .A(n10017), .B(n10016), .Z(n10288) );
  OR U10597 ( .A(n10019), .B(n10018), .Z(n10023) );
  NANDN U10598 ( .A(n10021), .B(n10020), .Z(n10022) );
  AND U10599 ( .A(n10023), .B(n10022), .Z(n10387) );
  AND U10600 ( .A(\stack[1][32] ), .B(o[17]), .Z(n10388) );
  XNOR U10601 ( .A(n10387), .B(n10388), .Z(n10390) );
  OR U10602 ( .A(n10025), .B(n10024), .Z(n10029) );
  OR U10603 ( .A(n10027), .B(n10026), .Z(n10028) );
  AND U10604 ( .A(n10029), .B(n10028), .Z(n10293) );
  NANDN U10605 ( .A(n10031), .B(n10030), .Z(n10035) );
  OR U10606 ( .A(n10033), .B(n10032), .Z(n10034) );
  NAND U10607 ( .A(n10035), .B(n10034), .Z(n10382) );
  ANDN U10608 ( .B(\stack[1][38] ), .A(n3005), .Z(n10314) );
  NANDN U10609 ( .A(n10037), .B(n10036), .Z(n10041) );
  NANDN U10610 ( .A(n10039), .B(n10038), .Z(n10040) );
  AND U10611 ( .A(n10041), .B(n10040), .Z(n10311) );
  AND U10612 ( .A(\stack[1][39] ), .B(o[10]), .Z(n10320) );
  AND U10613 ( .A(\stack[1][40] ), .B(o[9]), .Z(n10371) );
  NANDN U10614 ( .A(n10043), .B(n10042), .Z(n10047) );
  NAND U10615 ( .A(n10045), .B(n10044), .Z(n10046) );
  AND U10616 ( .A(n10047), .B(n10046), .Z(n10360) );
  AND U10617 ( .A(\stack[1][44] ), .B(o[5]), .Z(n10354) );
  OR U10618 ( .A(n10049), .B(n10048), .Z(n10053) );
  NANDN U10619 ( .A(n10051), .B(n10050), .Z(n10052) );
  AND U10620 ( .A(n10053), .B(n10052), .Z(n10351) );
  AND U10621 ( .A(\stack[1][45] ), .B(o[4]), .Z(n10332) );
  AND U10622 ( .A(\stack[1][46] ), .B(o[3]), .Z(n10348) );
  NANDN U10623 ( .A(n10054), .B(n10335), .Z(n10055) );
  AND U10624 ( .A(n10056), .B(n10055), .Z(n10060) );
  OR U10625 ( .A(n10058), .B(n10057), .Z(n10059) );
  AND U10626 ( .A(n10060), .B(n10059), .Z(n10345) );
  AND U10627 ( .A(\stack[1][49] ), .B(o[1]), .Z(n10343) );
  ANDN U10628 ( .B(n10343), .A(n10061), .Z(n10638) );
  XNOR U10629 ( .A(n10638), .B(n10335), .Z(n10063) );
  NAND U10630 ( .A(o[0]), .B(\stack[1][49] ), .Z(n10342) );
  NANDN U10631 ( .A(n10062), .B(n10342), .Z(n10337) );
  NAND U10632 ( .A(n10063), .B(n10337), .Z(n10339) );
  AND U10633 ( .A(\stack[1][47] ), .B(o[2]), .Z(n10338) );
  XNOR U10634 ( .A(n10339), .B(n10338), .Z(n10346) );
  XOR U10635 ( .A(n10345), .B(n10346), .Z(n10347) );
  XOR U10636 ( .A(n10348), .B(n10347), .Z(n10330) );
  OR U10637 ( .A(n10065), .B(n10064), .Z(n10069) );
  NANDN U10638 ( .A(n10067), .B(n10066), .Z(n10068) );
  AND U10639 ( .A(n10069), .B(n10068), .Z(n10329) );
  XOR U10640 ( .A(n10330), .B(n10329), .Z(n10331) );
  XOR U10641 ( .A(n10332), .B(n10331), .Z(n10352) );
  XNOR U10642 ( .A(n10351), .B(n10352), .Z(n10353) );
  OR U10643 ( .A(n10071), .B(n10070), .Z(n10075) );
  OR U10644 ( .A(n10073), .B(n10072), .Z(n10074) );
  NAND U10645 ( .A(n10075), .B(n10074), .Z(n10324) );
  IV U10646 ( .A(\stack[1][43] ), .Z(n15818) );
  ANDN U10647 ( .B(o[6]), .A(n15818), .Z(n10323) );
  XNOR U10648 ( .A(n10324), .B(n10323), .Z(n10326) );
  XNOR U10649 ( .A(n10325), .B(n10326), .Z(n10358) );
  ANDN U10650 ( .B(o[7]), .A(n15857), .Z(n10357) );
  XOR U10651 ( .A(n10358), .B(n10357), .Z(n10359) );
  NANDN U10652 ( .A(n10077), .B(n10076), .Z(n10081) );
  OR U10653 ( .A(n10079), .B(n10078), .Z(n10080) );
  AND U10654 ( .A(n10081), .B(n10080), .Z(n10363) );
  XNOR U10655 ( .A(n10364), .B(n10363), .Z(n10366) );
  AND U10656 ( .A(\stack[1][41] ), .B(o[8]), .Z(n10365) );
  XNOR U10657 ( .A(n10366), .B(n10365), .Z(n10369) );
  OR U10658 ( .A(n10083), .B(n10082), .Z(n10087) );
  NANDN U10659 ( .A(n10085), .B(n10084), .Z(n10086) );
  NAND U10660 ( .A(n10087), .B(n10086), .Z(n10370) );
  XNOR U10661 ( .A(n10369), .B(n10370), .Z(n10372) );
  XNOR U10662 ( .A(n10371), .B(n10372), .Z(n10318) );
  NANDN U10663 ( .A(n10089), .B(n10088), .Z(n10093) );
  NANDN U10664 ( .A(n10091), .B(n10090), .Z(n10092) );
  AND U10665 ( .A(n10093), .B(n10092), .Z(n10317) );
  XOR U10666 ( .A(n10318), .B(n10317), .Z(n10319) );
  XOR U10667 ( .A(n10320), .B(n10319), .Z(n10312) );
  XNOR U10668 ( .A(n10311), .B(n10312), .Z(n10313) );
  OR U10669 ( .A(n10095), .B(n10094), .Z(n10099) );
  NANDN U10670 ( .A(n10097), .B(n10096), .Z(n10098) );
  NAND U10671 ( .A(n10099), .B(n10098), .Z(n10376) );
  ANDN U10672 ( .B(\stack[1][37] ), .A(n3006), .Z(n10375) );
  XOR U10673 ( .A(n10376), .B(n10375), .Z(n10378) );
  OR U10674 ( .A(n10101), .B(n10100), .Z(n10105) );
  NANDN U10675 ( .A(n10103), .B(n10102), .Z(n10104) );
  AND U10676 ( .A(n10105), .B(n10104), .Z(n10305) );
  AND U10677 ( .A(\stack[1][36] ), .B(o[13]), .Z(n10306) );
  XNOR U10678 ( .A(n10305), .B(n10306), .Z(n10308) );
  XOR U10679 ( .A(n10307), .B(n10308), .Z(n10381) );
  XOR U10680 ( .A(n10382), .B(n10381), .Z(n10384) );
  AND U10681 ( .A(\stack[1][35] ), .B(o[14]), .Z(n10383) );
  XNOR U10682 ( .A(n10384), .B(n10383), .Z(n10301) );
  AND U10683 ( .A(\stack[1][34] ), .B(o[15]), .Z(n10299) );
  NANDN U10684 ( .A(n10107), .B(n10106), .Z(n10111) );
  NANDN U10685 ( .A(n10109), .B(n10108), .Z(n10110) );
  NAND U10686 ( .A(n10111), .B(n10110), .Z(n10300) );
  XNOR U10687 ( .A(n10299), .B(n10300), .Z(n10302) );
  XNOR U10688 ( .A(n10301), .B(n10302), .Z(n10294) );
  XOR U10689 ( .A(n10293), .B(n10294), .Z(n10295) );
  AND U10690 ( .A(\stack[1][33] ), .B(o[16]), .Z(n10296) );
  XOR U10691 ( .A(n10295), .B(n10296), .Z(n10389) );
  XOR U10692 ( .A(n10390), .B(n10389), .Z(n10287) );
  XNOR U10693 ( .A(n10288), .B(n10287), .Z(n10289) );
  XNOR U10694 ( .A(n10290), .B(n10289), .Z(n10283) );
  NANDN U10695 ( .A(n2987), .B(o[19]), .Z(n10281) );
  OR U10696 ( .A(n10113), .B(n10112), .Z(n10117) );
  OR U10697 ( .A(n10115), .B(n10114), .Z(n10116) );
  NAND U10698 ( .A(n10117), .B(n10116), .Z(n10282) );
  XOR U10699 ( .A(n10281), .B(n10282), .Z(n10284) );
  XNOR U10700 ( .A(n10283), .B(n10284), .Z(n10393) );
  XNOR U10701 ( .A(n10394), .B(n10393), .Z(n10395) );
  XNOR U10702 ( .A(n10396), .B(n10395), .Z(n10277) );
  NANDN U10703 ( .A(n2985), .B(o[21]), .Z(n10275) );
  OR U10704 ( .A(n10119), .B(n10118), .Z(n10123) );
  OR U10705 ( .A(n10121), .B(n10120), .Z(n10122) );
  NAND U10706 ( .A(n10123), .B(n10122), .Z(n10276) );
  XOR U10707 ( .A(n10275), .B(n10276), .Z(n10278) );
  XNOR U10708 ( .A(n10277), .B(n10278), .Z(n10399) );
  XNOR U10709 ( .A(n10400), .B(n10399), .Z(n10401) );
  XOR U10710 ( .A(n10402), .B(n10401), .Z(n10271) );
  AND U10711 ( .A(\stack[1][26] ), .B(o[23]), .Z(n10269) );
  NANDN U10712 ( .A(n10125), .B(n10124), .Z(n10129) );
  OR U10713 ( .A(n10127), .B(n10126), .Z(n10128) );
  NAND U10714 ( .A(n10129), .B(n10128), .Z(n10270) );
  XNOR U10715 ( .A(n10269), .B(n10270), .Z(n10272) );
  XNOR U10716 ( .A(n10405), .B(n10406), .Z(n10407) );
  XNOR U10717 ( .A(n10408), .B(n10407), .Z(n10265) );
  OR U10718 ( .A(n10131), .B(n10130), .Z(n10134) );
  OR U10719 ( .A(n10132), .B(n16555), .Z(n10133) );
  AND U10720 ( .A(n10134), .B(n10133), .Z(n10264) );
  NANDN U10721 ( .A(n3019), .B(\stack[1][24] ), .Z(n10263) );
  XOR U10722 ( .A(n10264), .B(n10263), .Z(n10266) );
  XNOR U10723 ( .A(n10265), .B(n10266), .Z(n10411) );
  XNOR U10724 ( .A(n10412), .B(n10411), .Z(n10413) );
  XNOR U10725 ( .A(n10414), .B(n10413), .Z(n10259) );
  NANDN U10726 ( .A(n2979), .B(o[27]), .Z(n10257) );
  OR U10727 ( .A(n10136), .B(n10135), .Z(n10140) );
  OR U10728 ( .A(n10138), .B(n10137), .Z(n10139) );
  NAND U10729 ( .A(n10140), .B(n10139), .Z(n10258) );
  XOR U10730 ( .A(n10257), .B(n10258), .Z(n10260) );
  XNOR U10731 ( .A(n10259), .B(n10260), .Z(n10417) );
  XNOR U10732 ( .A(n10418), .B(n10417), .Z(n10419) );
  XNOR U10733 ( .A(n10420), .B(n10419), .Z(n10253) );
  NANDN U10734 ( .A(n16712), .B(o[29]), .Z(n10251) );
  OR U10735 ( .A(n10142), .B(n10141), .Z(n10146) );
  OR U10736 ( .A(n10144), .B(n10143), .Z(n10145) );
  NAND U10737 ( .A(n10146), .B(n10145), .Z(n10252) );
  XOR U10738 ( .A(n10251), .B(n10252), .Z(n10254) );
  XNOR U10739 ( .A(n10253), .B(n10254), .Z(n10423) );
  XNOR U10740 ( .A(n10424), .B(n10423), .Z(n10425) );
  XNOR U10741 ( .A(n10426), .B(n10425), .Z(n10247) );
  NANDN U10742 ( .A(n16786), .B(o[31]), .Z(n10245) );
  OR U10743 ( .A(n10148), .B(n10147), .Z(n10152) );
  OR U10744 ( .A(n10150), .B(n10149), .Z(n10151) );
  NAND U10745 ( .A(n10152), .B(n10151), .Z(n10246) );
  XOR U10746 ( .A(n10245), .B(n10246), .Z(n10248) );
  XNOR U10747 ( .A(n10247), .B(n10248), .Z(n10429) );
  XNOR U10748 ( .A(n10430), .B(n10429), .Z(n10431) );
  XNOR U10749 ( .A(n10432), .B(n10431), .Z(n10241) );
  NANDN U10750 ( .A(n2977), .B(o[33]), .Z(n10239) );
  OR U10751 ( .A(n10154), .B(n10153), .Z(n10158) );
  OR U10752 ( .A(n10156), .B(n10155), .Z(n10157) );
  NAND U10753 ( .A(n10158), .B(n10157), .Z(n10240) );
  XOR U10754 ( .A(n10239), .B(n10240), .Z(n10242) );
  XNOR U10755 ( .A(n10241), .B(n10242), .Z(n10435) );
  XNOR U10756 ( .A(n10436), .B(n10435), .Z(n10437) );
  XNOR U10757 ( .A(n10438), .B(n10437), .Z(n10235) );
  NANDN U10758 ( .A(n2975), .B(o[35]), .Z(n10233) );
  OR U10759 ( .A(n10160), .B(n10159), .Z(n10164) );
  OR U10760 ( .A(n10162), .B(n10161), .Z(n10163) );
  NAND U10761 ( .A(n10164), .B(n10163), .Z(n10234) );
  XOR U10762 ( .A(n10233), .B(n10234), .Z(n10236) );
  XNOR U10763 ( .A(n10235), .B(n10236), .Z(n10442) );
  XNOR U10764 ( .A(n10441), .B(n10442), .Z(n10443) );
  XOR U10765 ( .A(n10229), .B(n10230), .Z(n10447) );
  OR U10766 ( .A(n10166), .B(n10165), .Z(n10170) );
  NANDN U10767 ( .A(n10168), .B(n10167), .Z(n10169) );
  AND U10768 ( .A(n10170), .B(n10169), .Z(n10448) );
  XOR U10769 ( .A(n10447), .B(n10448), .Z(n10450) );
  AND U10770 ( .A(o[38]), .B(\stack[1][11] ), .Z(n10449) );
  XOR U10771 ( .A(n10450), .B(n10449), .Z(n10223) );
  XOR U10772 ( .A(n10224), .B(n10223), .Z(n10454) );
  XOR U10773 ( .A(n10453), .B(n10454), .Z(n10455) );
  XOR U10774 ( .A(n10456), .B(n10455), .Z(n10218) );
  AND U10775 ( .A(o[41]), .B(\stack[1][8] ), .Z(n10215) );
  OR U10776 ( .A(n10172), .B(n10171), .Z(n10176) );
  OR U10777 ( .A(n10174), .B(n10173), .Z(n10175) );
  NAND U10778 ( .A(n10176), .B(n10175), .Z(n10216) );
  XNOR U10779 ( .A(n10215), .B(n10216), .Z(n10217) );
  XOR U10780 ( .A(n10218), .B(n10217), .Z(n10459) );
  XNOR U10781 ( .A(n10460), .B(n10459), .Z(n10461) );
  XNOR U10782 ( .A(n10462), .B(n10461), .Z(n10211) );
  NANDN U10783 ( .A(n17256), .B(o[43]), .Z(n10209) );
  OR U10784 ( .A(n10178), .B(n10177), .Z(n10182) );
  OR U10785 ( .A(n10180), .B(n10179), .Z(n10181) );
  NAND U10786 ( .A(n10182), .B(n10181), .Z(n10210) );
  XOR U10787 ( .A(n10209), .B(n10210), .Z(n10212) );
  XNOR U10788 ( .A(n10211), .B(n10212), .Z(n10465) );
  XNOR U10789 ( .A(n10466), .B(n10465), .Z(n10467) );
  XNOR U10790 ( .A(n10468), .B(n10467), .Z(n10205) );
  AND U10791 ( .A(o[45]), .B(\stack[1][4] ), .Z(n10203) );
  OR U10792 ( .A(n10184), .B(n10183), .Z(n10188) );
  OR U10793 ( .A(n10186), .B(n10185), .Z(n10187) );
  NAND U10794 ( .A(n10188), .B(n10187), .Z(n10204) );
  XNOR U10795 ( .A(n10203), .B(n10204), .Z(n10206) );
  XNOR U10796 ( .A(n10205), .B(n10206), .Z(n10471) );
  XNOR U10797 ( .A(n10472), .B(n10471), .Z(n10473) );
  XOR U10798 ( .A(n10474), .B(n10473), .Z(n10200) );
  AND U10799 ( .A(o[47]), .B(\stack[1][2] ), .Z(n10197) );
  OR U10800 ( .A(n10190), .B(n10189), .Z(n10194) );
  OR U10801 ( .A(n10192), .B(n10191), .Z(n10193) );
  NAND U10802 ( .A(n10194), .B(n10193), .Z(n10198) );
  XOR U10803 ( .A(n10197), .B(n10198), .Z(n10199) );
  XNOR U10804 ( .A(n10200), .B(n10199), .Z(n10477) );
  XNOR U10805 ( .A(n10478), .B(n10477), .Z(n10479) );
  XOR U10806 ( .A(n10480), .B(n10479), .Z(n15588) );
  OR U10807 ( .A(n15587), .B(n15588), .Z(n10195) );
  AND U10808 ( .A(n10196), .B(n10195), .Z(n10484) );
  NANDN U10809 ( .A(n2970), .B(o[48]), .Z(n10777) );
  OR U10810 ( .A(n10198), .B(n10197), .Z(n10202) );
  NANDN U10811 ( .A(n10200), .B(n10199), .Z(n10201) );
  NAND U10812 ( .A(n10202), .B(n10201), .Z(n10775) );
  NANDN U10813 ( .A(n2971), .B(o[46]), .Z(n10771) );
  OR U10814 ( .A(n10204), .B(n10203), .Z(n10208) );
  NANDN U10815 ( .A(n10206), .B(n10205), .Z(n10207) );
  NAND U10816 ( .A(n10208), .B(n10207), .Z(n10769) );
  NANDN U10817 ( .A(n17256), .B(o[44]), .Z(n10765) );
  NANDN U10818 ( .A(n10210), .B(n10209), .Z(n10214) );
  NANDN U10819 ( .A(n10212), .B(n10211), .Z(n10213) );
  NAND U10820 ( .A(n10214), .B(n10213), .Z(n10763) );
  NANDN U10821 ( .A(n17179), .B(o[42]), .Z(n10759) );
  OR U10822 ( .A(n10216), .B(n10215), .Z(n10220) );
  OR U10823 ( .A(n10218), .B(n10217), .Z(n10219) );
  NAND U10824 ( .A(n10220), .B(n10219), .Z(n10757) );
  NANDN U10825 ( .A(n17101), .B(o[40]), .Z(n10753) );
  OR U10826 ( .A(n10222), .B(n10221), .Z(n10226) );
  NANDN U10827 ( .A(n10224), .B(n10223), .Z(n10225) );
  NAND U10828 ( .A(n10226), .B(n10225), .Z(n10751) );
  NANDN U10829 ( .A(n2973), .B(o[38]), .Z(n10747) );
  NANDN U10830 ( .A(n10228), .B(n10227), .Z(n10232) );
  NANDN U10831 ( .A(n10230), .B(n10229), .Z(n10231) );
  AND U10832 ( .A(n10232), .B(n10231), .Z(n10744) );
  NANDN U10833 ( .A(n2975), .B(o[36]), .Z(n10741) );
  NANDN U10834 ( .A(n10234), .B(n10233), .Z(n10238) );
  NANDN U10835 ( .A(n10236), .B(n10235), .Z(n10237) );
  NAND U10836 ( .A(n10238), .B(n10237), .Z(n10739) );
  NANDN U10837 ( .A(n2977), .B(o[34]), .Z(n10735) );
  NANDN U10838 ( .A(n10240), .B(n10239), .Z(n10244) );
  NANDN U10839 ( .A(n10242), .B(n10241), .Z(n10243) );
  NAND U10840 ( .A(n10244), .B(n10243), .Z(n10733) );
  NANDN U10841 ( .A(n16786), .B(o[32]), .Z(n10729) );
  NANDN U10842 ( .A(n10246), .B(n10245), .Z(n10250) );
  NANDN U10843 ( .A(n10248), .B(n10247), .Z(n10249) );
  NAND U10844 ( .A(n10250), .B(n10249), .Z(n10727) );
  NANDN U10845 ( .A(n16712), .B(o[30]), .Z(n10723) );
  NANDN U10846 ( .A(n10252), .B(n10251), .Z(n10256) );
  NANDN U10847 ( .A(n10254), .B(n10253), .Z(n10255) );
  NAND U10848 ( .A(n10256), .B(n10255), .Z(n10721) );
  NANDN U10849 ( .A(n2979), .B(o[28]), .Z(n10717) );
  NANDN U10850 ( .A(n10258), .B(n10257), .Z(n10262) );
  NANDN U10851 ( .A(n10260), .B(n10259), .Z(n10261) );
  NAND U10852 ( .A(n10262), .B(n10261), .Z(n10715) );
  NANDN U10853 ( .A(n2981), .B(o[26]), .Z(n10711) );
  NANDN U10854 ( .A(n10264), .B(n10263), .Z(n10268) );
  NANDN U10855 ( .A(n10266), .B(n10265), .Z(n10267) );
  NAND U10856 ( .A(n10268), .B(n10267), .Z(n10709) );
  NANDN U10857 ( .A(n3018), .B(\stack[1][26] ), .Z(n10705) );
  OR U10858 ( .A(n10270), .B(n10269), .Z(n10274) );
  OR U10859 ( .A(n10272), .B(n10271), .Z(n10273) );
  NAND U10860 ( .A(n10274), .B(n10273), .Z(n10703) );
  NANDN U10861 ( .A(n3016), .B(\stack[1][28] ), .Z(n10699) );
  NANDN U10862 ( .A(n10276), .B(n10275), .Z(n10280) );
  NANDN U10863 ( .A(n10278), .B(n10277), .Z(n10279) );
  NAND U10864 ( .A(n10280), .B(n10279), .Z(n10697) );
  AND U10865 ( .A(\stack[1][30] ), .B(o[20]), .Z(n10693) );
  NANDN U10866 ( .A(n10282), .B(n10281), .Z(n10286) );
  NANDN U10867 ( .A(n10284), .B(n10283), .Z(n10285) );
  AND U10868 ( .A(n10286), .B(n10285), .Z(n10690) );
  AND U10869 ( .A(\stack[1][31] ), .B(o[19]), .Z(n10578) );
  OR U10870 ( .A(n10288), .B(n10287), .Z(n10292) );
  OR U10871 ( .A(n10290), .B(n10289), .Z(n10291) );
  NAND U10872 ( .A(n10292), .B(n10291), .Z(n10579) );
  XNOR U10873 ( .A(n10578), .B(n10579), .Z(n10581) );
  OR U10874 ( .A(n10294), .B(n10293), .Z(n10298) );
  NANDN U10875 ( .A(n10296), .B(n10295), .Z(n10297) );
  NAND U10876 ( .A(n10298), .B(n10297), .Z(n10585) );
  ANDN U10877 ( .B(o[17]), .A(n2990), .Z(n10584) );
  XOR U10878 ( .A(n10585), .B(n10584), .Z(n10586) );
  NANDN U10879 ( .A(n3010), .B(\stack[1][34] ), .Z(n10593) );
  OR U10880 ( .A(n10300), .B(n10299), .Z(n10304) );
  OR U10881 ( .A(n10302), .B(n10301), .Z(n10303) );
  NAND U10882 ( .A(n10304), .B(n10303), .Z(n10591) );
  NANDN U10883 ( .A(n3008), .B(\stack[1][36] ), .Z(n10681) );
  OR U10884 ( .A(n10306), .B(n10305), .Z(n10310) );
  NANDN U10885 ( .A(n10308), .B(n10307), .Z(n10309) );
  NAND U10886 ( .A(n10310), .B(n10309), .Z(n10679) );
  ANDN U10887 ( .B(\stack[1][38] ), .A(n3006), .Z(n10611) );
  OR U10888 ( .A(n10312), .B(n10311), .Z(n10316) );
  OR U10889 ( .A(n10314), .B(n10313), .Z(n10315) );
  AND U10890 ( .A(n10316), .B(n10315), .Z(n10608) );
  AND U10891 ( .A(\stack[1][39] ), .B(o[11]), .Z(n10617) );
  OR U10892 ( .A(n10318), .B(n10317), .Z(n10322) );
  NANDN U10893 ( .A(n10320), .B(n10319), .Z(n10321) );
  AND U10894 ( .A(n10322), .B(n10321), .Z(n10614) );
  AND U10895 ( .A(\stack[1][40] ), .B(o[10]), .Z(n10623) );
  AND U10896 ( .A(\stack[1][41] ), .B(o[9]), .Z(n10674) );
  NANDN U10897 ( .A(n10324), .B(n10323), .Z(n10328) );
  NAND U10898 ( .A(n10326), .B(n10325), .Z(n10327) );
  AND U10899 ( .A(n10328), .B(n10327), .Z(n10663) );
  AND U10900 ( .A(\stack[1][45] ), .B(o[5]), .Z(n10657) );
  OR U10901 ( .A(n10330), .B(n10329), .Z(n10334) );
  NANDN U10902 ( .A(n10332), .B(n10331), .Z(n10333) );
  AND U10903 ( .A(n10334), .B(n10333), .Z(n10654) );
  AND U10904 ( .A(\stack[1][46] ), .B(o[4]), .Z(n10635) );
  AND U10905 ( .A(\stack[1][47] ), .B(o[3]), .Z(n10651) );
  NANDN U10906 ( .A(n10335), .B(n10638), .Z(n10336) );
  AND U10907 ( .A(n10337), .B(n10336), .Z(n10341) );
  OR U10908 ( .A(n10339), .B(n10338), .Z(n10340) );
  AND U10909 ( .A(n10341), .B(n10340), .Z(n10648) );
  AND U10910 ( .A(\stack[1][50] ), .B(o[1]), .Z(n10646) );
  ANDN U10911 ( .B(n10646), .A(n10342), .Z(n10932) );
  XNOR U10912 ( .A(n10932), .B(n10638), .Z(n10344) );
  NAND U10913 ( .A(\stack[1][50] ), .B(o[0]), .Z(n10645) );
  NANDN U10914 ( .A(n10343), .B(n10645), .Z(n10640) );
  NAND U10915 ( .A(n10344), .B(n10640), .Z(n10642) );
  AND U10916 ( .A(\stack[1][48] ), .B(o[2]), .Z(n10641) );
  XNOR U10917 ( .A(n10642), .B(n10641), .Z(n10649) );
  XOR U10918 ( .A(n10648), .B(n10649), .Z(n10650) );
  XOR U10919 ( .A(n10651), .B(n10650), .Z(n10633) );
  OR U10920 ( .A(n10346), .B(n10345), .Z(n10350) );
  NANDN U10921 ( .A(n10348), .B(n10347), .Z(n10349) );
  AND U10922 ( .A(n10350), .B(n10349), .Z(n10632) );
  XOR U10923 ( .A(n10633), .B(n10632), .Z(n10634) );
  XOR U10924 ( .A(n10635), .B(n10634), .Z(n10655) );
  XNOR U10925 ( .A(n10654), .B(n10655), .Z(n10656) );
  OR U10926 ( .A(n10352), .B(n10351), .Z(n10356) );
  OR U10927 ( .A(n10354), .B(n10353), .Z(n10355) );
  NAND U10928 ( .A(n10356), .B(n10355), .Z(n10627) );
  IV U10929 ( .A(\stack[1][44] ), .Z(n15779) );
  ANDN U10930 ( .B(o[6]), .A(n15779), .Z(n10626) );
  XNOR U10931 ( .A(n10627), .B(n10626), .Z(n10629) );
  XNOR U10932 ( .A(n10628), .B(n10629), .Z(n10661) );
  ANDN U10933 ( .B(o[7]), .A(n15818), .Z(n10660) );
  XOR U10934 ( .A(n10661), .B(n10660), .Z(n10662) );
  NANDN U10935 ( .A(n10358), .B(n10357), .Z(n10362) );
  OR U10936 ( .A(n10360), .B(n10359), .Z(n10361) );
  AND U10937 ( .A(n10362), .B(n10361), .Z(n10666) );
  XNOR U10938 ( .A(n10667), .B(n10666), .Z(n10669) );
  AND U10939 ( .A(\stack[1][42] ), .B(o[8]), .Z(n10668) );
  XNOR U10940 ( .A(n10669), .B(n10668), .Z(n10672) );
  OR U10941 ( .A(n10364), .B(n10363), .Z(n10368) );
  NANDN U10942 ( .A(n10366), .B(n10365), .Z(n10367) );
  NAND U10943 ( .A(n10368), .B(n10367), .Z(n10673) );
  XNOR U10944 ( .A(n10672), .B(n10673), .Z(n10675) );
  XNOR U10945 ( .A(n10674), .B(n10675), .Z(n10621) );
  OR U10946 ( .A(n10370), .B(n10369), .Z(n10374) );
  OR U10947 ( .A(n10372), .B(n10371), .Z(n10373) );
  AND U10948 ( .A(n10374), .B(n10373), .Z(n10620) );
  XOR U10949 ( .A(n10621), .B(n10620), .Z(n10622) );
  XOR U10950 ( .A(n10623), .B(n10622), .Z(n10615) );
  XOR U10951 ( .A(n10614), .B(n10615), .Z(n10616) );
  XOR U10952 ( .A(n10617), .B(n10616), .Z(n10609) );
  XOR U10953 ( .A(n10608), .B(n10609), .Z(n10610) );
  XOR U10954 ( .A(n10611), .B(n10610), .Z(n10605) );
  AND U10955 ( .A(\stack[1][37] ), .B(o[13]), .Z(n10602) );
  NANDN U10956 ( .A(n10376), .B(n10375), .Z(n10380) );
  NANDN U10957 ( .A(n10378), .B(n10377), .Z(n10379) );
  NAND U10958 ( .A(n10380), .B(n10379), .Z(n10603) );
  XNOR U10959 ( .A(n10602), .B(n10603), .Z(n10604) );
  XOR U10960 ( .A(n10605), .B(n10604), .Z(n10678) );
  XNOR U10961 ( .A(n10679), .B(n10678), .Z(n10680) );
  XNOR U10962 ( .A(n10681), .B(n10680), .Z(n10598) );
  AND U10963 ( .A(\stack[1][35] ), .B(o[15]), .Z(n10596) );
  NANDN U10964 ( .A(n10382), .B(n10381), .Z(n10386) );
  NANDN U10965 ( .A(n10384), .B(n10383), .Z(n10385) );
  NAND U10966 ( .A(n10386), .B(n10385), .Z(n10597) );
  XNOR U10967 ( .A(n10596), .B(n10597), .Z(n10599) );
  XNOR U10968 ( .A(n10598), .B(n10599), .Z(n10590) );
  XNOR U10969 ( .A(n10591), .B(n10590), .Z(n10592) );
  XNOR U10970 ( .A(n10593), .B(n10592), .Z(n10587) );
  OR U10971 ( .A(n10388), .B(n10387), .Z(n10392) );
  OR U10972 ( .A(n10390), .B(n10389), .Z(n10391) );
  AND U10973 ( .A(n10392), .B(n10391), .Z(n10685) );
  XNOR U10974 ( .A(n10684), .B(n10685), .Z(n10687) );
  AND U10975 ( .A(\stack[1][32] ), .B(o[18]), .Z(n10686) );
  XOR U10976 ( .A(n10687), .B(n10686), .Z(n10580) );
  XOR U10977 ( .A(n10581), .B(n10580), .Z(n10691) );
  XOR U10978 ( .A(n10690), .B(n10691), .Z(n10692) );
  XOR U10979 ( .A(n10693), .B(n10692), .Z(n10575) );
  AND U10980 ( .A(\stack[1][29] ), .B(o[21]), .Z(n10572) );
  OR U10981 ( .A(n10394), .B(n10393), .Z(n10398) );
  OR U10982 ( .A(n10396), .B(n10395), .Z(n10397) );
  NAND U10983 ( .A(n10398), .B(n10397), .Z(n10573) );
  XNOR U10984 ( .A(n10572), .B(n10573), .Z(n10574) );
  XOR U10985 ( .A(n10575), .B(n10574), .Z(n10696) );
  XNOR U10986 ( .A(n10697), .B(n10696), .Z(n10698) );
  XNOR U10987 ( .A(n10699), .B(n10698), .Z(n10568) );
  NANDN U10988 ( .A(n2984), .B(o[23]), .Z(n10566) );
  OR U10989 ( .A(n10400), .B(n10399), .Z(n10404) );
  OR U10990 ( .A(n10402), .B(n10401), .Z(n10403) );
  NAND U10991 ( .A(n10404), .B(n10403), .Z(n10567) );
  XOR U10992 ( .A(n10566), .B(n10567), .Z(n10569) );
  XNOR U10993 ( .A(n10568), .B(n10569), .Z(n10702) );
  XNOR U10994 ( .A(n10703), .B(n10702), .Z(n10704) );
  XNOR U10995 ( .A(n10705), .B(n10704), .Z(n10562) );
  AND U10996 ( .A(o[25]), .B(\stack[1][25] ), .Z(n16514) );
  OR U10997 ( .A(n10406), .B(n10405), .Z(n10410) );
  OR U10998 ( .A(n10408), .B(n10407), .Z(n10409) );
  NAND U10999 ( .A(n10410), .B(n10409), .Z(n10561) );
  XNOR U11000 ( .A(n16514), .B(n10561), .Z(n10563) );
  XNOR U11001 ( .A(n10562), .B(n10563), .Z(n10708) );
  XNOR U11002 ( .A(n10709), .B(n10708), .Z(n10710) );
  XNOR U11003 ( .A(n10711), .B(n10710), .Z(n10557) );
  NANDN U11004 ( .A(n2980), .B(o[27]), .Z(n10555) );
  OR U11005 ( .A(n10412), .B(n10411), .Z(n10416) );
  OR U11006 ( .A(n10414), .B(n10413), .Z(n10415) );
  NAND U11007 ( .A(n10416), .B(n10415), .Z(n10556) );
  XOR U11008 ( .A(n10555), .B(n10556), .Z(n10558) );
  XNOR U11009 ( .A(n10557), .B(n10558), .Z(n10714) );
  XNOR U11010 ( .A(n10715), .B(n10714), .Z(n10716) );
  XNOR U11011 ( .A(n10717), .B(n10716), .Z(n10551) );
  NANDN U11012 ( .A(n2978), .B(o[29]), .Z(n10549) );
  OR U11013 ( .A(n10418), .B(n10417), .Z(n10422) );
  OR U11014 ( .A(n10420), .B(n10419), .Z(n10421) );
  NAND U11015 ( .A(n10422), .B(n10421), .Z(n10550) );
  XOR U11016 ( .A(n10549), .B(n10550), .Z(n10552) );
  XNOR U11017 ( .A(n10551), .B(n10552), .Z(n10720) );
  XNOR U11018 ( .A(n10721), .B(n10720), .Z(n10722) );
  XNOR U11019 ( .A(n10723), .B(n10722), .Z(n10545) );
  NANDN U11020 ( .A(n16746), .B(o[31]), .Z(n10543) );
  OR U11021 ( .A(n10424), .B(n10423), .Z(n10428) );
  OR U11022 ( .A(n10426), .B(n10425), .Z(n10427) );
  NAND U11023 ( .A(n10428), .B(n10427), .Z(n10544) );
  XOR U11024 ( .A(n10543), .B(n10544), .Z(n10546) );
  XNOR U11025 ( .A(n10545), .B(n10546), .Z(n10726) );
  XNOR U11026 ( .A(n10727), .B(n10726), .Z(n10728) );
  XNOR U11027 ( .A(n10729), .B(n10728), .Z(n10539) );
  NANDN U11028 ( .A(n16826), .B(o[33]), .Z(n10537) );
  OR U11029 ( .A(n10430), .B(n10429), .Z(n10434) );
  OR U11030 ( .A(n10432), .B(n10431), .Z(n10433) );
  NAND U11031 ( .A(n10434), .B(n10433), .Z(n10538) );
  XOR U11032 ( .A(n10537), .B(n10538), .Z(n10540) );
  XNOR U11033 ( .A(n10539), .B(n10540), .Z(n10732) );
  XNOR U11034 ( .A(n10733), .B(n10732), .Z(n10734) );
  XNOR U11035 ( .A(n10735), .B(n10734), .Z(n10533) );
  NANDN U11036 ( .A(n2976), .B(o[35]), .Z(n10531) );
  OR U11037 ( .A(n10436), .B(n10435), .Z(n10440) );
  OR U11038 ( .A(n10438), .B(n10437), .Z(n10439) );
  NAND U11039 ( .A(n10440), .B(n10439), .Z(n10532) );
  XOR U11040 ( .A(n10531), .B(n10532), .Z(n10534) );
  XNOR U11041 ( .A(n10533), .B(n10534), .Z(n10738) );
  XNOR U11042 ( .A(n10739), .B(n10738), .Z(n10740) );
  XOR U11043 ( .A(n10741), .B(n10740), .Z(n10527) );
  AND U11044 ( .A(o[37]), .B(\stack[1][13] ), .Z(n10525) );
  OR U11045 ( .A(n10442), .B(n10441), .Z(n10446) );
  OR U11046 ( .A(n10444), .B(n10443), .Z(n10445) );
  NAND U11047 ( .A(n10446), .B(n10445), .Z(n10526) );
  XNOR U11048 ( .A(n10525), .B(n10526), .Z(n10528) );
  XNOR U11049 ( .A(n10744), .B(n10745), .Z(n10746) );
  XNOR U11050 ( .A(n10747), .B(n10746), .Z(n10521) );
  NANDN U11051 ( .A(n10448), .B(n10447), .Z(n10452) );
  OR U11052 ( .A(n10450), .B(n10449), .Z(n10451) );
  AND U11053 ( .A(n10452), .B(n10451), .Z(n10520) );
  NANDN U11054 ( .A(n2972), .B(o[39]), .Z(n10519) );
  XOR U11055 ( .A(n10520), .B(n10519), .Z(n10522) );
  XNOR U11056 ( .A(n10521), .B(n10522), .Z(n10750) );
  XNOR U11057 ( .A(n10751), .B(n10750), .Z(n10752) );
  XNOR U11058 ( .A(n10753), .B(n10752), .Z(n10515) );
  OR U11059 ( .A(n10454), .B(n10453), .Z(n10458) );
  NANDN U11060 ( .A(n10456), .B(n10455), .Z(n10457) );
  AND U11061 ( .A(n10458), .B(n10457), .Z(n10514) );
  NANDN U11062 ( .A(n17145), .B(o[41]), .Z(n10513) );
  XOR U11063 ( .A(n10514), .B(n10513), .Z(n10516) );
  XNOR U11064 ( .A(n10515), .B(n10516), .Z(n10756) );
  XNOR U11065 ( .A(n10757), .B(n10756), .Z(n10758) );
  XNOR U11066 ( .A(n10759), .B(n10758), .Z(n10509) );
  NANDN U11067 ( .A(n17219), .B(o[43]), .Z(n10507) );
  OR U11068 ( .A(n10460), .B(n10459), .Z(n10464) );
  OR U11069 ( .A(n10462), .B(n10461), .Z(n10463) );
  NAND U11070 ( .A(n10464), .B(n10463), .Z(n10508) );
  XOR U11071 ( .A(n10507), .B(n10508), .Z(n10510) );
  XNOR U11072 ( .A(n10509), .B(n10510), .Z(n10762) );
  XNOR U11073 ( .A(n10763), .B(n10762), .Z(n10764) );
  XNOR U11074 ( .A(n10765), .B(n10764), .Z(n10503) );
  NANDN U11075 ( .A(n17296), .B(o[45]), .Z(n10501) );
  OR U11076 ( .A(n10466), .B(n10465), .Z(n10470) );
  OR U11077 ( .A(n10468), .B(n10467), .Z(n10469) );
  NAND U11078 ( .A(n10470), .B(n10469), .Z(n10502) );
  XOR U11079 ( .A(n10501), .B(n10502), .Z(n10504) );
  XNOR U11080 ( .A(n10503), .B(n10504), .Z(n10768) );
  XNOR U11081 ( .A(n10769), .B(n10768), .Z(n10770) );
  XNOR U11082 ( .A(n10771), .B(n10770), .Z(n10497) );
  NANDN U11083 ( .A(n17375), .B(o[47]), .Z(n10495) );
  OR U11084 ( .A(n10472), .B(n10471), .Z(n10476) );
  OR U11085 ( .A(n10474), .B(n10473), .Z(n10475) );
  NAND U11086 ( .A(n10476), .B(n10475), .Z(n10496) );
  XOR U11087 ( .A(n10495), .B(n10496), .Z(n10498) );
  XNOR U11088 ( .A(n10497), .B(n10498), .Z(n10774) );
  XNOR U11089 ( .A(n10775), .B(n10774), .Z(n10776) );
  AND U11090 ( .A(o[49]), .B(\stack[1][1] ), .Z(n10489) );
  OR U11091 ( .A(n10478), .B(n10477), .Z(n10482) );
  OR U11092 ( .A(n10480), .B(n10479), .Z(n10481) );
  NAND U11093 ( .A(n10482), .B(n10481), .Z(n10490) );
  XNOR U11094 ( .A(n10489), .B(n10490), .Z(n10492) );
  XOR U11095 ( .A(n10491), .B(n10492), .Z(n10483) );
  NANDN U11096 ( .A(n10484), .B(n10483), .Z(n10486) );
  XOR U11097 ( .A(n10484), .B(n10483), .Z(n15549) );
  AND U11098 ( .A(o[50]), .B(\stack[1][0] ), .Z(n15550) );
  OR U11099 ( .A(n15549), .B(n15550), .Z(n10485) );
  AND U11100 ( .A(n10486), .B(n10485), .Z(n10488) );
  OR U11101 ( .A(n10487), .B(n10488), .Z(n10781) );
  XNOR U11102 ( .A(n10488), .B(n10487), .Z(n15510) );
  NANDN U11103 ( .A(n2969), .B(o[50]), .Z(n11077) );
  OR U11104 ( .A(n10490), .B(n10489), .Z(n10494) );
  OR U11105 ( .A(n10492), .B(n10491), .Z(n10493) );
  NAND U11106 ( .A(n10494), .B(n10493), .Z(n11075) );
  NANDN U11107 ( .A(n17375), .B(o[48]), .Z(n11071) );
  NANDN U11108 ( .A(n10496), .B(n10495), .Z(n10500) );
  NANDN U11109 ( .A(n10498), .B(n10497), .Z(n10499) );
  NAND U11110 ( .A(n10500), .B(n10499), .Z(n11069) );
  NANDN U11111 ( .A(n17296), .B(o[46]), .Z(n11065) );
  NANDN U11112 ( .A(n10502), .B(n10501), .Z(n10506) );
  NANDN U11113 ( .A(n10504), .B(n10503), .Z(n10505) );
  NAND U11114 ( .A(n10506), .B(n10505), .Z(n11063) );
  NANDN U11115 ( .A(n17219), .B(o[44]), .Z(n11059) );
  NANDN U11116 ( .A(n10508), .B(n10507), .Z(n10512) );
  NANDN U11117 ( .A(n10510), .B(n10509), .Z(n10511) );
  NAND U11118 ( .A(n10512), .B(n10511), .Z(n11057) );
  NANDN U11119 ( .A(n17145), .B(o[42]), .Z(n11053) );
  NANDN U11120 ( .A(n10514), .B(n10513), .Z(n10518) );
  NANDN U11121 ( .A(n10516), .B(n10515), .Z(n10517) );
  NAND U11122 ( .A(n10518), .B(n10517), .Z(n11051) );
  NANDN U11123 ( .A(n2972), .B(o[40]), .Z(n11047) );
  NANDN U11124 ( .A(n10520), .B(n10519), .Z(n10524) );
  NANDN U11125 ( .A(n10522), .B(n10521), .Z(n10523) );
  NAND U11126 ( .A(n10524), .B(n10523), .Z(n11045) );
  NANDN U11127 ( .A(n2974), .B(o[38]), .Z(n11041) );
  OR U11128 ( .A(n10526), .B(n10525), .Z(n10530) );
  OR U11129 ( .A(n10528), .B(n10527), .Z(n10529) );
  NAND U11130 ( .A(n10530), .B(n10529), .Z(n11039) );
  NANDN U11131 ( .A(n2976), .B(o[36]), .Z(n11035) );
  NANDN U11132 ( .A(n10532), .B(n10531), .Z(n10536) );
  NANDN U11133 ( .A(n10534), .B(n10533), .Z(n10535) );
  NAND U11134 ( .A(n10536), .B(n10535), .Z(n11033) );
  NANDN U11135 ( .A(n16826), .B(o[34]), .Z(n11029) );
  NANDN U11136 ( .A(n10538), .B(n10537), .Z(n10542) );
  NANDN U11137 ( .A(n10540), .B(n10539), .Z(n10541) );
  NAND U11138 ( .A(n10542), .B(n10541), .Z(n11027) );
  NANDN U11139 ( .A(n16746), .B(o[32]), .Z(n11023) );
  NANDN U11140 ( .A(n10544), .B(n10543), .Z(n10548) );
  NANDN U11141 ( .A(n10546), .B(n10545), .Z(n10547) );
  NAND U11142 ( .A(n10548), .B(n10547), .Z(n11021) );
  NANDN U11143 ( .A(n2978), .B(o[30]), .Z(n11017) );
  NANDN U11144 ( .A(n10550), .B(n10549), .Z(n10554) );
  NANDN U11145 ( .A(n10552), .B(n10551), .Z(n10553) );
  NAND U11146 ( .A(n10554), .B(n10553), .Z(n11015) );
  NANDN U11147 ( .A(n2980), .B(o[28]), .Z(n11011) );
  NANDN U11148 ( .A(n10556), .B(n10555), .Z(n10560) );
  NANDN U11149 ( .A(n10558), .B(n10557), .Z(n10559) );
  NAND U11150 ( .A(n10560), .B(n10559), .Z(n11009) );
  NANDN U11151 ( .A(n2982), .B(o[26]), .Z(n11005) );
  OR U11152 ( .A(n10561), .B(n16514), .Z(n10565) );
  NANDN U11153 ( .A(n10563), .B(n10562), .Z(n10564) );
  NAND U11154 ( .A(n10565), .B(n10564), .Z(n11003) );
  NANDN U11155 ( .A(n3018), .B(\stack[1][27] ), .Z(n10999) );
  NANDN U11156 ( .A(n10567), .B(n10566), .Z(n10571) );
  NANDN U11157 ( .A(n10569), .B(n10568), .Z(n10570) );
  NAND U11158 ( .A(n10571), .B(n10570), .Z(n10997) );
  NANDN U11159 ( .A(n3016), .B(\stack[1][29] ), .Z(n10993) );
  OR U11160 ( .A(n10573), .B(n10572), .Z(n10577) );
  OR U11161 ( .A(n10575), .B(n10574), .Z(n10576) );
  NAND U11162 ( .A(n10577), .B(n10576), .Z(n10991) );
  NANDN U11163 ( .A(n3014), .B(\stack[1][31] ), .Z(n10987) );
  OR U11164 ( .A(n10579), .B(n10578), .Z(n10583) );
  NANDN U11165 ( .A(n10581), .B(n10580), .Z(n10582) );
  NAND U11166 ( .A(n10583), .B(n10582), .Z(n10985) );
  NANDN U11167 ( .A(n3012), .B(\stack[1][33] ), .Z(n10981) );
  NANDN U11168 ( .A(n10585), .B(n10584), .Z(n10589) );
  OR U11169 ( .A(n10587), .B(n10586), .Z(n10588) );
  AND U11170 ( .A(n10589), .B(n10588), .Z(n10978) );
  AND U11171 ( .A(\stack[1][34] ), .B(o[17]), .Z(n10878) );
  OR U11172 ( .A(n10591), .B(n10590), .Z(n10595) );
  OR U11173 ( .A(n10593), .B(n10592), .Z(n10594) );
  NAND U11174 ( .A(n10595), .B(n10594), .Z(n10879) );
  XNOR U11175 ( .A(n10878), .B(n10879), .Z(n10881) );
  OR U11176 ( .A(n10597), .B(n10596), .Z(n10601) );
  NANDN U11177 ( .A(n10599), .B(n10598), .Z(n10600) );
  AND U11178 ( .A(n10601), .B(n10600), .Z(n10972) );
  OR U11179 ( .A(n10603), .B(n10602), .Z(n10607) );
  OR U11180 ( .A(n10605), .B(n10604), .Z(n10606) );
  NAND U11181 ( .A(n10607), .B(n10606), .Z(n10891) );
  ANDN U11182 ( .B(\stack[1][38] ), .A(n3007), .Z(n10899) );
  OR U11183 ( .A(n10609), .B(n10608), .Z(n10613) );
  NANDN U11184 ( .A(n10611), .B(n10610), .Z(n10612) );
  AND U11185 ( .A(n10613), .B(n10612), .Z(n10896) );
  OR U11186 ( .A(n10615), .B(n10614), .Z(n10619) );
  NANDN U11187 ( .A(n10617), .B(n10616), .Z(n10618) );
  NAND U11188 ( .A(n10619), .B(n10618), .Z(n10905) );
  AND U11189 ( .A(\stack[1][40] ), .B(o[11]), .Z(n10911) );
  OR U11190 ( .A(n10621), .B(n10620), .Z(n10625) );
  NANDN U11191 ( .A(n10623), .B(n10622), .Z(n10624) );
  AND U11192 ( .A(n10625), .B(n10624), .Z(n10908) );
  AND U11193 ( .A(\stack[1][41] ), .B(o[10]), .Z(n10917) );
  AND U11194 ( .A(\stack[1][42] ), .B(o[9]), .Z(n10968) );
  NANDN U11195 ( .A(n10627), .B(n10626), .Z(n10631) );
  NAND U11196 ( .A(n10629), .B(n10628), .Z(n10630) );
  AND U11197 ( .A(n10631), .B(n10630), .Z(n10957) );
  AND U11198 ( .A(\stack[1][46] ), .B(o[5]), .Z(n10951) );
  OR U11199 ( .A(n10633), .B(n10632), .Z(n10637) );
  NANDN U11200 ( .A(n10635), .B(n10634), .Z(n10636) );
  AND U11201 ( .A(n10637), .B(n10636), .Z(n10948) );
  AND U11202 ( .A(\stack[1][47] ), .B(o[4]), .Z(n10929) );
  AND U11203 ( .A(\stack[1][48] ), .B(o[3]), .Z(n10945) );
  NANDN U11204 ( .A(n10638), .B(n10932), .Z(n10639) );
  AND U11205 ( .A(n10640), .B(n10639), .Z(n10644) );
  OR U11206 ( .A(n10642), .B(n10641), .Z(n10643) );
  AND U11207 ( .A(n10644), .B(n10643), .Z(n10942) );
  AND U11208 ( .A(\stack[1][51] ), .B(o[1]), .Z(n10940) );
  ANDN U11209 ( .B(n10940), .A(n10645), .Z(n11242) );
  XNOR U11210 ( .A(n11242), .B(n10932), .Z(n10647) );
  NAND U11211 ( .A(\stack[1][51] ), .B(o[0]), .Z(n10939) );
  NANDN U11212 ( .A(n10646), .B(n10939), .Z(n10934) );
  NAND U11213 ( .A(n10647), .B(n10934), .Z(n10936) );
  ANDN U11214 ( .B(\stack[1][49] ), .A(n2996), .Z(n10935) );
  XNOR U11215 ( .A(n10936), .B(n10935), .Z(n10943) );
  XOR U11216 ( .A(n10942), .B(n10943), .Z(n10944) );
  XOR U11217 ( .A(n10945), .B(n10944), .Z(n10927) );
  OR U11218 ( .A(n10649), .B(n10648), .Z(n10653) );
  NANDN U11219 ( .A(n10651), .B(n10650), .Z(n10652) );
  AND U11220 ( .A(n10653), .B(n10652), .Z(n10926) );
  XOR U11221 ( .A(n10927), .B(n10926), .Z(n10928) );
  XOR U11222 ( .A(n10929), .B(n10928), .Z(n10949) );
  XNOR U11223 ( .A(n10948), .B(n10949), .Z(n10950) );
  OR U11224 ( .A(n10655), .B(n10654), .Z(n10659) );
  OR U11225 ( .A(n10657), .B(n10656), .Z(n10658) );
  NAND U11226 ( .A(n10659), .B(n10658), .Z(n10921) );
  IV U11227 ( .A(\stack[1][45] ), .Z(n15740) );
  ANDN U11228 ( .B(o[6]), .A(n15740), .Z(n10920) );
  XNOR U11229 ( .A(n10921), .B(n10920), .Z(n10923) );
  XNOR U11230 ( .A(n10922), .B(n10923), .Z(n10955) );
  ANDN U11231 ( .B(o[7]), .A(n15779), .Z(n10954) );
  XOR U11232 ( .A(n10955), .B(n10954), .Z(n10956) );
  NANDN U11233 ( .A(n10661), .B(n10660), .Z(n10665) );
  OR U11234 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U11235 ( .A(n10665), .B(n10664), .Z(n10960) );
  XNOR U11236 ( .A(n10961), .B(n10960), .Z(n10963) );
  AND U11237 ( .A(\stack[1][43] ), .B(o[8]), .Z(n10962) );
  XNOR U11238 ( .A(n10963), .B(n10962), .Z(n10966) );
  OR U11239 ( .A(n10667), .B(n10666), .Z(n10671) );
  NANDN U11240 ( .A(n10669), .B(n10668), .Z(n10670) );
  NAND U11241 ( .A(n10671), .B(n10670), .Z(n10967) );
  XNOR U11242 ( .A(n10966), .B(n10967), .Z(n10969) );
  XNOR U11243 ( .A(n10968), .B(n10969), .Z(n10915) );
  OR U11244 ( .A(n10673), .B(n10672), .Z(n10677) );
  OR U11245 ( .A(n10675), .B(n10674), .Z(n10676) );
  AND U11246 ( .A(n10677), .B(n10676), .Z(n10914) );
  XOR U11247 ( .A(n10915), .B(n10914), .Z(n10916) );
  XOR U11248 ( .A(n10917), .B(n10916), .Z(n10909) );
  XNOR U11249 ( .A(n10908), .B(n10909), .Z(n10910) );
  NANDN U11250 ( .A(n3006), .B(\stack[1][39] ), .Z(n10903) );
  XOR U11251 ( .A(n10902), .B(n10903), .Z(n10904) );
  XOR U11252 ( .A(n10905), .B(n10904), .Z(n10897) );
  XNOR U11253 ( .A(n10896), .B(n10897), .Z(n10898) );
  XOR U11254 ( .A(n10891), .B(n10890), .Z(n10893) );
  AND U11255 ( .A(\stack[1][37] ), .B(o[14]), .Z(n10892) );
  XNOR U11256 ( .A(n10893), .B(n10892), .Z(n10886) );
  AND U11257 ( .A(\stack[1][36] ), .B(o[15]), .Z(n10884) );
  OR U11258 ( .A(n10679), .B(n10678), .Z(n10683) );
  OR U11259 ( .A(n10681), .B(n10680), .Z(n10682) );
  NAND U11260 ( .A(n10683), .B(n10682), .Z(n10885) );
  XNOR U11261 ( .A(n10884), .B(n10885), .Z(n10887) );
  XNOR U11262 ( .A(n10886), .B(n10887), .Z(n10973) );
  XNOR U11263 ( .A(n10972), .B(n10973), .Z(n10974) );
  AND U11264 ( .A(\stack[1][35] ), .B(o[16]), .Z(n10975) );
  XOR U11265 ( .A(n10881), .B(n10880), .Z(n10979) );
  XNOR U11266 ( .A(n10978), .B(n10979), .Z(n10980) );
  XNOR U11267 ( .A(n10981), .B(n10980), .Z(n10874) );
  OR U11268 ( .A(n10685), .B(n10684), .Z(n10689) );
  OR U11269 ( .A(n10687), .B(n10686), .Z(n10688) );
  AND U11270 ( .A(n10689), .B(n10688), .Z(n10873) );
  NANDN U11271 ( .A(n2989), .B(o[19]), .Z(n10872) );
  XOR U11272 ( .A(n10873), .B(n10872), .Z(n10875) );
  XNOR U11273 ( .A(n10874), .B(n10875), .Z(n10984) );
  XNOR U11274 ( .A(n10985), .B(n10984), .Z(n10986) );
  XNOR U11275 ( .A(n10987), .B(n10986), .Z(n10868) );
  OR U11276 ( .A(n10691), .B(n10690), .Z(n10695) );
  NANDN U11277 ( .A(n10693), .B(n10692), .Z(n10694) );
  AND U11278 ( .A(n10695), .B(n10694), .Z(n10867) );
  NANDN U11279 ( .A(n2987), .B(o[21]), .Z(n10866) );
  XOR U11280 ( .A(n10867), .B(n10866), .Z(n10869) );
  XNOR U11281 ( .A(n10868), .B(n10869), .Z(n10990) );
  XNOR U11282 ( .A(n10991), .B(n10990), .Z(n10992) );
  XNOR U11283 ( .A(n10993), .B(n10992), .Z(n10862) );
  NANDN U11284 ( .A(n2985), .B(o[23]), .Z(n10860) );
  OR U11285 ( .A(n10697), .B(n10696), .Z(n10701) );
  OR U11286 ( .A(n10699), .B(n10698), .Z(n10700) );
  NAND U11287 ( .A(n10701), .B(n10700), .Z(n10861) );
  XOR U11288 ( .A(n10860), .B(n10861), .Z(n10863) );
  XNOR U11289 ( .A(n10862), .B(n10863), .Z(n10996) );
  XNOR U11290 ( .A(n10997), .B(n10996), .Z(n10998) );
  XNOR U11291 ( .A(n10999), .B(n10998), .Z(n10856) );
  NANDN U11292 ( .A(n2983), .B(o[25]), .Z(n10854) );
  OR U11293 ( .A(n10703), .B(n10702), .Z(n10707) );
  OR U11294 ( .A(n10705), .B(n10704), .Z(n10706) );
  NAND U11295 ( .A(n10707), .B(n10706), .Z(n10855) );
  XOR U11296 ( .A(n10854), .B(n10855), .Z(n10857) );
  XNOR U11297 ( .A(n10856), .B(n10857), .Z(n11002) );
  XNOR U11298 ( .A(n11003), .B(n11002), .Z(n11004) );
  XNOR U11299 ( .A(n11005), .B(n11004), .Z(n10850) );
  NANDN U11300 ( .A(n2981), .B(o[27]), .Z(n10848) );
  OR U11301 ( .A(n10709), .B(n10708), .Z(n10713) );
  OR U11302 ( .A(n10711), .B(n10710), .Z(n10712) );
  NAND U11303 ( .A(n10713), .B(n10712), .Z(n10849) );
  XOR U11304 ( .A(n10848), .B(n10849), .Z(n10851) );
  XNOR U11305 ( .A(n10850), .B(n10851), .Z(n11008) );
  XNOR U11306 ( .A(n11009), .B(n11008), .Z(n11010) );
  XNOR U11307 ( .A(n11011), .B(n11010), .Z(n10844) );
  NANDN U11308 ( .A(n2979), .B(o[29]), .Z(n10842) );
  OR U11309 ( .A(n10715), .B(n10714), .Z(n10719) );
  OR U11310 ( .A(n10717), .B(n10716), .Z(n10718) );
  NAND U11311 ( .A(n10719), .B(n10718), .Z(n10843) );
  XOR U11312 ( .A(n10842), .B(n10843), .Z(n10845) );
  XNOR U11313 ( .A(n10844), .B(n10845), .Z(n11014) );
  XNOR U11314 ( .A(n11015), .B(n11014), .Z(n11016) );
  XNOR U11315 ( .A(n11017), .B(n11016), .Z(n10838) );
  NANDN U11316 ( .A(n16712), .B(o[31]), .Z(n10836) );
  OR U11317 ( .A(n10721), .B(n10720), .Z(n10725) );
  OR U11318 ( .A(n10723), .B(n10722), .Z(n10724) );
  NAND U11319 ( .A(n10725), .B(n10724), .Z(n10837) );
  XOR U11320 ( .A(n10836), .B(n10837), .Z(n10839) );
  XNOR U11321 ( .A(n10838), .B(n10839), .Z(n11020) );
  XNOR U11322 ( .A(n11021), .B(n11020), .Z(n11022) );
  XNOR U11323 ( .A(n11023), .B(n11022), .Z(n10832) );
  NANDN U11324 ( .A(n16786), .B(o[33]), .Z(n10830) );
  OR U11325 ( .A(n10727), .B(n10726), .Z(n10731) );
  OR U11326 ( .A(n10729), .B(n10728), .Z(n10730) );
  NAND U11327 ( .A(n10731), .B(n10730), .Z(n10831) );
  XOR U11328 ( .A(n10830), .B(n10831), .Z(n10833) );
  XNOR U11329 ( .A(n10832), .B(n10833), .Z(n11026) );
  XNOR U11330 ( .A(n11027), .B(n11026), .Z(n11028) );
  XNOR U11331 ( .A(n11029), .B(n11028), .Z(n10826) );
  NANDN U11332 ( .A(n2977), .B(o[35]), .Z(n10824) );
  OR U11333 ( .A(n10733), .B(n10732), .Z(n10737) );
  OR U11334 ( .A(n10735), .B(n10734), .Z(n10736) );
  NAND U11335 ( .A(n10737), .B(n10736), .Z(n10825) );
  XOR U11336 ( .A(n10824), .B(n10825), .Z(n10827) );
  XNOR U11337 ( .A(n10826), .B(n10827), .Z(n11032) );
  XNOR U11338 ( .A(n11033), .B(n11032), .Z(n11034) );
  XNOR U11339 ( .A(n11035), .B(n11034), .Z(n10820) );
  NANDN U11340 ( .A(n2975), .B(o[37]), .Z(n10818) );
  OR U11341 ( .A(n10739), .B(n10738), .Z(n10743) );
  OR U11342 ( .A(n10741), .B(n10740), .Z(n10742) );
  NAND U11343 ( .A(n10743), .B(n10742), .Z(n10819) );
  XOR U11344 ( .A(n10818), .B(n10819), .Z(n10821) );
  XNOR U11345 ( .A(n10820), .B(n10821), .Z(n11038) );
  XNOR U11346 ( .A(n11039), .B(n11038), .Z(n11040) );
  XNOR U11347 ( .A(n11041), .B(n11040), .Z(n10814) );
  NANDN U11348 ( .A(n2973), .B(o[39]), .Z(n10812) );
  OR U11349 ( .A(n10745), .B(n10744), .Z(n10749) );
  OR U11350 ( .A(n10747), .B(n10746), .Z(n10748) );
  NAND U11351 ( .A(n10749), .B(n10748), .Z(n10813) );
  XOR U11352 ( .A(n10812), .B(n10813), .Z(n10815) );
  XNOR U11353 ( .A(n10814), .B(n10815), .Z(n11044) );
  XNOR U11354 ( .A(n11045), .B(n11044), .Z(n11046) );
  XNOR U11355 ( .A(n11047), .B(n11046), .Z(n10808) );
  NANDN U11356 ( .A(n17101), .B(o[41]), .Z(n10806) );
  OR U11357 ( .A(n10751), .B(n10750), .Z(n10755) );
  OR U11358 ( .A(n10753), .B(n10752), .Z(n10754) );
  NAND U11359 ( .A(n10755), .B(n10754), .Z(n10807) );
  XOR U11360 ( .A(n10806), .B(n10807), .Z(n10809) );
  XNOR U11361 ( .A(n10808), .B(n10809), .Z(n11050) );
  XNOR U11362 ( .A(n11051), .B(n11050), .Z(n11052) );
  XNOR U11363 ( .A(n11053), .B(n11052), .Z(n10802) );
  NANDN U11364 ( .A(n17179), .B(o[43]), .Z(n10800) );
  OR U11365 ( .A(n10757), .B(n10756), .Z(n10761) );
  OR U11366 ( .A(n10759), .B(n10758), .Z(n10760) );
  NAND U11367 ( .A(n10761), .B(n10760), .Z(n10801) );
  XOR U11368 ( .A(n10800), .B(n10801), .Z(n10803) );
  XNOR U11369 ( .A(n10802), .B(n10803), .Z(n11056) );
  XNOR U11370 ( .A(n11057), .B(n11056), .Z(n11058) );
  XNOR U11371 ( .A(n11059), .B(n11058), .Z(n10796) );
  NANDN U11372 ( .A(n17256), .B(o[45]), .Z(n10794) );
  OR U11373 ( .A(n10763), .B(n10762), .Z(n10767) );
  OR U11374 ( .A(n10765), .B(n10764), .Z(n10766) );
  NAND U11375 ( .A(n10767), .B(n10766), .Z(n10795) );
  XOR U11376 ( .A(n10794), .B(n10795), .Z(n10797) );
  XNOR U11377 ( .A(n10796), .B(n10797), .Z(n11062) );
  XNOR U11378 ( .A(n11063), .B(n11062), .Z(n11064) );
  XNOR U11379 ( .A(n11065), .B(n11064), .Z(n10790) );
  AND U11380 ( .A(o[47]), .B(\stack[1][4] ), .Z(n10788) );
  OR U11381 ( .A(n10769), .B(n10768), .Z(n10773) );
  OR U11382 ( .A(n10771), .B(n10770), .Z(n10772) );
  NAND U11383 ( .A(n10773), .B(n10772), .Z(n10789) );
  XNOR U11384 ( .A(n10788), .B(n10789), .Z(n10791) );
  XNOR U11385 ( .A(n10790), .B(n10791), .Z(n11068) );
  XNOR U11386 ( .A(n11069), .B(n11068), .Z(n11070) );
  XOR U11387 ( .A(n11071), .B(n11070), .Z(n10785) );
  AND U11388 ( .A(o[49]), .B(\stack[1][2] ), .Z(n10782) );
  OR U11389 ( .A(n10775), .B(n10774), .Z(n10779) );
  OR U11390 ( .A(n10777), .B(n10776), .Z(n10778) );
  NAND U11391 ( .A(n10779), .B(n10778), .Z(n10783) );
  XOR U11392 ( .A(n10782), .B(n10783), .Z(n10784) );
  XNOR U11393 ( .A(n10785), .B(n10784), .Z(n11074) );
  XNOR U11394 ( .A(n11075), .B(n11074), .Z(n11076) );
  XOR U11395 ( .A(n11077), .B(n11076), .Z(n15511) );
  OR U11396 ( .A(n15510), .B(n15511), .Z(n10780) );
  AND U11397 ( .A(n10781), .B(n10780), .Z(n11081) );
  NANDN U11398 ( .A(n2970), .B(o[50]), .Z(n11387) );
  OR U11399 ( .A(n10783), .B(n10782), .Z(n10787) );
  NANDN U11400 ( .A(n10785), .B(n10784), .Z(n10786) );
  NAND U11401 ( .A(n10787), .B(n10786), .Z(n11385) );
  NANDN U11402 ( .A(n2971), .B(o[48]), .Z(n11381) );
  OR U11403 ( .A(n10789), .B(n10788), .Z(n10793) );
  NANDN U11404 ( .A(n10791), .B(n10790), .Z(n10792) );
  NAND U11405 ( .A(n10793), .B(n10792), .Z(n11379) );
  NANDN U11406 ( .A(n17256), .B(o[46]), .Z(n11375) );
  NANDN U11407 ( .A(n10795), .B(n10794), .Z(n10799) );
  NANDN U11408 ( .A(n10797), .B(n10796), .Z(n10798) );
  NAND U11409 ( .A(n10799), .B(n10798), .Z(n11373) );
  NANDN U11410 ( .A(n17179), .B(o[44]), .Z(n11369) );
  NANDN U11411 ( .A(n10801), .B(n10800), .Z(n10805) );
  NANDN U11412 ( .A(n10803), .B(n10802), .Z(n10804) );
  NAND U11413 ( .A(n10805), .B(n10804), .Z(n11367) );
  NANDN U11414 ( .A(n17101), .B(o[42]), .Z(n11363) );
  NANDN U11415 ( .A(n10807), .B(n10806), .Z(n10811) );
  NANDN U11416 ( .A(n10809), .B(n10808), .Z(n10810) );
  NAND U11417 ( .A(n10811), .B(n10810), .Z(n11361) );
  NANDN U11418 ( .A(n2973), .B(o[40]), .Z(n11357) );
  NANDN U11419 ( .A(n10813), .B(n10812), .Z(n10817) );
  NANDN U11420 ( .A(n10815), .B(n10814), .Z(n10816) );
  NAND U11421 ( .A(n10817), .B(n10816), .Z(n11355) );
  NANDN U11422 ( .A(n2975), .B(o[38]), .Z(n11351) );
  NANDN U11423 ( .A(n10819), .B(n10818), .Z(n10823) );
  NANDN U11424 ( .A(n10821), .B(n10820), .Z(n10822) );
  NAND U11425 ( .A(n10823), .B(n10822), .Z(n11349) );
  NANDN U11426 ( .A(n2977), .B(o[36]), .Z(n11345) );
  NANDN U11427 ( .A(n10825), .B(n10824), .Z(n10829) );
  NANDN U11428 ( .A(n10827), .B(n10826), .Z(n10828) );
  NAND U11429 ( .A(n10829), .B(n10828), .Z(n11343) );
  NANDN U11430 ( .A(n16786), .B(o[34]), .Z(n11339) );
  NANDN U11431 ( .A(n10831), .B(n10830), .Z(n10835) );
  NANDN U11432 ( .A(n10833), .B(n10832), .Z(n10834) );
  NAND U11433 ( .A(n10835), .B(n10834), .Z(n11337) );
  NANDN U11434 ( .A(n16712), .B(o[32]), .Z(n11333) );
  NANDN U11435 ( .A(n10837), .B(n10836), .Z(n10841) );
  NANDN U11436 ( .A(n10839), .B(n10838), .Z(n10840) );
  NAND U11437 ( .A(n10841), .B(n10840), .Z(n11331) );
  NANDN U11438 ( .A(n2979), .B(o[30]), .Z(n11327) );
  NANDN U11439 ( .A(n10843), .B(n10842), .Z(n10847) );
  NANDN U11440 ( .A(n10845), .B(n10844), .Z(n10846) );
  NAND U11441 ( .A(n10847), .B(n10846), .Z(n11325) );
  NANDN U11442 ( .A(n2981), .B(o[28]), .Z(n11321) );
  NANDN U11443 ( .A(n10849), .B(n10848), .Z(n10853) );
  NANDN U11444 ( .A(n10851), .B(n10850), .Z(n10852) );
  NAND U11445 ( .A(n10853), .B(n10852), .Z(n11319) );
  NOR U11446 ( .A(n3020), .B(n2983), .Z(n11314) );
  NANDN U11447 ( .A(n10855), .B(n10854), .Z(n10859) );
  NANDN U11448 ( .A(n10857), .B(n10856), .Z(n10858) );
  NAND U11449 ( .A(n10859), .B(n10858), .Z(n11313) );
  NANDN U11450 ( .A(n3018), .B(\stack[1][28] ), .Z(n11309) );
  NANDN U11451 ( .A(n10861), .B(n10860), .Z(n10865) );
  NANDN U11452 ( .A(n10863), .B(n10862), .Z(n10864) );
  NAND U11453 ( .A(n10865), .B(n10864), .Z(n11307) );
  NANDN U11454 ( .A(n3016), .B(\stack[1][30] ), .Z(n11303) );
  NANDN U11455 ( .A(n10867), .B(n10866), .Z(n10871) );
  NANDN U11456 ( .A(n10869), .B(n10868), .Z(n10870) );
  NAND U11457 ( .A(n10871), .B(n10870), .Z(n11301) );
  NANDN U11458 ( .A(n3014), .B(\stack[1][32] ), .Z(n11297) );
  NANDN U11459 ( .A(n10873), .B(n10872), .Z(n10877) );
  NANDN U11460 ( .A(n10875), .B(n10874), .Z(n10876) );
  NAND U11461 ( .A(n10877), .B(n10876), .Z(n11295) );
  NANDN U11462 ( .A(n3012), .B(\stack[1][34] ), .Z(n11191) );
  OR U11463 ( .A(n10879), .B(n10878), .Z(n10883) );
  OR U11464 ( .A(n10881), .B(n10880), .Z(n10882) );
  NAND U11465 ( .A(n10883), .B(n10882), .Z(n11189) );
  AND U11466 ( .A(\stack[1][36] ), .B(o[16]), .Z(n11197) );
  OR U11467 ( .A(n10885), .B(n10884), .Z(n10889) );
  OR U11468 ( .A(n10887), .B(n10886), .Z(n10888) );
  AND U11469 ( .A(n10889), .B(n10888), .Z(n11194) );
  AND U11470 ( .A(\stack[1][37] ), .B(o[15]), .Z(n11200) );
  NANDN U11471 ( .A(n10891), .B(n10890), .Z(n10895) );
  NANDN U11472 ( .A(n10893), .B(n10892), .Z(n10894) );
  NAND U11473 ( .A(n10895), .B(n10894), .Z(n11201) );
  XNOR U11474 ( .A(n11200), .B(n11201), .Z(n11203) );
  NANDN U11475 ( .A(n3008), .B(\stack[1][38] ), .Z(n11208) );
  OR U11476 ( .A(n10897), .B(n10896), .Z(n10901) );
  OR U11477 ( .A(n10899), .B(n10898), .Z(n10900) );
  AND U11478 ( .A(n10901), .B(n10900), .Z(n11207) );
  NANDN U11479 ( .A(n10903), .B(n10902), .Z(n10907) );
  OR U11480 ( .A(n10905), .B(n10904), .Z(n10906) );
  AND U11481 ( .A(n10907), .B(n10906), .Z(n11285) );
  OR U11482 ( .A(n10909), .B(n10908), .Z(n10913) );
  OR U11483 ( .A(n10911), .B(n10910), .Z(n10912) );
  NAND U11484 ( .A(n10913), .B(n10912), .Z(n11215) );
  AND U11485 ( .A(\stack[1][41] ), .B(o[11]), .Z(n11221) );
  OR U11486 ( .A(n10915), .B(n10914), .Z(n10919) );
  NANDN U11487 ( .A(n10917), .B(n10916), .Z(n10918) );
  AND U11488 ( .A(n10919), .B(n10918), .Z(n11218) );
  AND U11489 ( .A(\stack[1][42] ), .B(o[10]), .Z(n11227) );
  AND U11490 ( .A(\stack[1][43] ), .B(o[9]), .Z(n11278) );
  NANDN U11491 ( .A(n10921), .B(n10920), .Z(n10925) );
  NAND U11492 ( .A(n10923), .B(n10922), .Z(n10924) );
  AND U11493 ( .A(n10925), .B(n10924), .Z(n11267) );
  AND U11494 ( .A(\stack[1][47] ), .B(o[5]), .Z(n11261) );
  OR U11495 ( .A(n10927), .B(n10926), .Z(n10931) );
  NANDN U11496 ( .A(n10929), .B(n10928), .Z(n10930) );
  AND U11497 ( .A(n10931), .B(n10930), .Z(n11258) );
  AND U11498 ( .A(\stack[1][48] ), .B(o[4]), .Z(n11239) );
  ANDN U11499 ( .B(\stack[1][49] ), .A(n2997), .Z(n11255) );
  NANDN U11500 ( .A(n10932), .B(n11242), .Z(n10933) );
  AND U11501 ( .A(n10934), .B(n10933), .Z(n10938) );
  OR U11502 ( .A(n10936), .B(n10935), .Z(n10937) );
  AND U11503 ( .A(n10938), .B(n10937), .Z(n11252) );
  AND U11504 ( .A(\stack[1][52] ), .B(o[1]), .Z(n11250) );
  ANDN U11505 ( .B(n11250), .A(n10939), .Z(n11542) );
  XNOR U11506 ( .A(n11542), .B(n11242), .Z(n10941) );
  NAND U11507 ( .A(\stack[1][52] ), .B(o[0]), .Z(n11249) );
  NANDN U11508 ( .A(n10940), .B(n11249), .Z(n11244) );
  NAND U11509 ( .A(n10941), .B(n11244), .Z(n11246) );
  AND U11510 ( .A(\stack[1][50] ), .B(o[2]), .Z(n11245) );
  XNOR U11511 ( .A(n11246), .B(n11245), .Z(n11253) );
  XOR U11512 ( .A(n11252), .B(n11253), .Z(n11254) );
  XOR U11513 ( .A(n11255), .B(n11254), .Z(n11237) );
  OR U11514 ( .A(n10943), .B(n10942), .Z(n10947) );
  NANDN U11515 ( .A(n10945), .B(n10944), .Z(n10946) );
  AND U11516 ( .A(n10947), .B(n10946), .Z(n11236) );
  XOR U11517 ( .A(n11237), .B(n11236), .Z(n11238) );
  XOR U11518 ( .A(n11239), .B(n11238), .Z(n11259) );
  XNOR U11519 ( .A(n11258), .B(n11259), .Z(n11260) );
  OR U11520 ( .A(n10949), .B(n10948), .Z(n10953) );
  OR U11521 ( .A(n10951), .B(n10950), .Z(n10952) );
  NAND U11522 ( .A(n10953), .B(n10952), .Z(n11231) );
  IV U11523 ( .A(\stack[1][46] ), .Z(n15701) );
  ANDN U11524 ( .B(o[6]), .A(n15701), .Z(n11230) );
  XNOR U11525 ( .A(n11231), .B(n11230), .Z(n11233) );
  XNOR U11526 ( .A(n11232), .B(n11233), .Z(n11265) );
  ANDN U11527 ( .B(o[7]), .A(n15740), .Z(n11264) );
  XOR U11528 ( .A(n11265), .B(n11264), .Z(n11266) );
  NANDN U11529 ( .A(n10955), .B(n10954), .Z(n10959) );
  OR U11530 ( .A(n10957), .B(n10956), .Z(n10958) );
  AND U11531 ( .A(n10959), .B(n10958), .Z(n11270) );
  XNOR U11532 ( .A(n11271), .B(n11270), .Z(n11273) );
  AND U11533 ( .A(\stack[1][44] ), .B(o[8]), .Z(n11272) );
  XNOR U11534 ( .A(n11273), .B(n11272), .Z(n11276) );
  OR U11535 ( .A(n10961), .B(n10960), .Z(n10965) );
  NANDN U11536 ( .A(n10963), .B(n10962), .Z(n10964) );
  NAND U11537 ( .A(n10965), .B(n10964), .Z(n11277) );
  XNOR U11538 ( .A(n11276), .B(n11277), .Z(n11279) );
  XNOR U11539 ( .A(n11278), .B(n11279), .Z(n11225) );
  OR U11540 ( .A(n10967), .B(n10966), .Z(n10971) );
  OR U11541 ( .A(n10969), .B(n10968), .Z(n10970) );
  AND U11542 ( .A(n10971), .B(n10970), .Z(n11224) );
  XOR U11543 ( .A(n11225), .B(n11224), .Z(n11226) );
  XOR U11544 ( .A(n11227), .B(n11226), .Z(n11219) );
  XOR U11545 ( .A(n11218), .B(n11219), .Z(n11220) );
  XOR U11546 ( .A(n11221), .B(n11220), .Z(n11213) );
  AND U11547 ( .A(\stack[1][40] ), .B(o[12]), .Z(n11212) );
  XNOR U11548 ( .A(n11213), .B(n11212), .Z(n11214) );
  XNOR U11549 ( .A(n11215), .B(n11214), .Z(n11283) );
  ANDN U11550 ( .B(\stack[1][39] ), .A(n3007), .Z(n11282) );
  XOR U11551 ( .A(n11283), .B(n11282), .Z(n11284) );
  XOR U11552 ( .A(n11207), .B(n11206), .Z(n11209) );
  XNOR U11553 ( .A(n11208), .B(n11209), .Z(n11202) );
  XOR U11554 ( .A(n11203), .B(n11202), .Z(n11195) );
  XOR U11555 ( .A(n11194), .B(n11195), .Z(n11196) );
  XOR U11556 ( .A(n11197), .B(n11196), .Z(n11291) );
  OR U11557 ( .A(n10973), .B(n10972), .Z(n10977) );
  OR U11558 ( .A(n10975), .B(n10974), .Z(n10976) );
  AND U11559 ( .A(n10977), .B(n10976), .Z(n11288) );
  AND U11560 ( .A(\stack[1][35] ), .B(o[17]), .Z(n11289) );
  XNOR U11561 ( .A(n11288), .B(n11289), .Z(n11290) );
  XOR U11562 ( .A(n11291), .B(n11290), .Z(n11188) );
  XNOR U11563 ( .A(n11189), .B(n11188), .Z(n11190) );
  XNOR U11564 ( .A(n11191), .B(n11190), .Z(n11184) );
  NANDN U11565 ( .A(n2990), .B(o[19]), .Z(n11182) );
  OR U11566 ( .A(n10979), .B(n10978), .Z(n10983) );
  OR U11567 ( .A(n10981), .B(n10980), .Z(n10982) );
  NAND U11568 ( .A(n10983), .B(n10982), .Z(n11183) );
  XOR U11569 ( .A(n11182), .B(n11183), .Z(n11185) );
  XNOR U11570 ( .A(n11184), .B(n11185), .Z(n11294) );
  XNOR U11571 ( .A(n11295), .B(n11294), .Z(n11296) );
  XNOR U11572 ( .A(n11297), .B(n11296), .Z(n11178) );
  NANDN U11573 ( .A(n2988), .B(o[21]), .Z(n11176) );
  OR U11574 ( .A(n10985), .B(n10984), .Z(n10989) );
  OR U11575 ( .A(n10987), .B(n10986), .Z(n10988) );
  NAND U11576 ( .A(n10989), .B(n10988), .Z(n11177) );
  XOR U11577 ( .A(n11176), .B(n11177), .Z(n11179) );
  XNOR U11578 ( .A(n11178), .B(n11179), .Z(n11300) );
  XNOR U11579 ( .A(n11301), .B(n11300), .Z(n11302) );
  XNOR U11580 ( .A(n11303), .B(n11302), .Z(n11172) );
  NANDN U11581 ( .A(n2986), .B(o[23]), .Z(n11170) );
  OR U11582 ( .A(n10991), .B(n10990), .Z(n10995) );
  OR U11583 ( .A(n10993), .B(n10992), .Z(n10994) );
  NAND U11584 ( .A(n10995), .B(n10994), .Z(n11171) );
  XOR U11585 ( .A(n11170), .B(n11171), .Z(n11173) );
  XNOR U11586 ( .A(n11172), .B(n11173), .Z(n11306) );
  XNOR U11587 ( .A(n11307), .B(n11306), .Z(n11308) );
  XNOR U11588 ( .A(n11309), .B(n11308), .Z(n11166) );
  NANDN U11589 ( .A(n2984), .B(o[25]), .Z(n11164) );
  OR U11590 ( .A(n10997), .B(n10996), .Z(n11001) );
  OR U11591 ( .A(n10999), .B(n10998), .Z(n11000) );
  NAND U11592 ( .A(n11001), .B(n11000), .Z(n11165) );
  XOR U11593 ( .A(n11164), .B(n11165), .Z(n11167) );
  XNOR U11594 ( .A(n11166), .B(n11167), .Z(n11312) );
  XNOR U11595 ( .A(n11313), .B(n11312), .Z(n11315) );
  XOR U11596 ( .A(n11314), .B(n11315), .Z(n11160) );
  NANDN U11597 ( .A(n2982), .B(o[27]), .Z(n11158) );
  OR U11598 ( .A(n11003), .B(n11002), .Z(n11007) );
  OR U11599 ( .A(n11005), .B(n11004), .Z(n11006) );
  NAND U11600 ( .A(n11007), .B(n11006), .Z(n11159) );
  XOR U11601 ( .A(n11158), .B(n11159), .Z(n11161) );
  XNOR U11602 ( .A(n11160), .B(n11161), .Z(n11318) );
  XNOR U11603 ( .A(n11319), .B(n11318), .Z(n11320) );
  XNOR U11604 ( .A(n11321), .B(n11320), .Z(n11154) );
  NANDN U11605 ( .A(n2980), .B(o[29]), .Z(n11152) );
  OR U11606 ( .A(n11009), .B(n11008), .Z(n11013) );
  OR U11607 ( .A(n11011), .B(n11010), .Z(n11012) );
  NAND U11608 ( .A(n11013), .B(n11012), .Z(n11153) );
  XOR U11609 ( .A(n11152), .B(n11153), .Z(n11155) );
  XNOR U11610 ( .A(n11154), .B(n11155), .Z(n11324) );
  XNOR U11611 ( .A(n11325), .B(n11324), .Z(n11326) );
  XNOR U11612 ( .A(n11327), .B(n11326), .Z(n11148) );
  NANDN U11613 ( .A(n2978), .B(o[31]), .Z(n11146) );
  OR U11614 ( .A(n11015), .B(n11014), .Z(n11019) );
  OR U11615 ( .A(n11017), .B(n11016), .Z(n11018) );
  NAND U11616 ( .A(n11019), .B(n11018), .Z(n11147) );
  XOR U11617 ( .A(n11146), .B(n11147), .Z(n11149) );
  XNOR U11618 ( .A(n11148), .B(n11149), .Z(n11330) );
  XNOR U11619 ( .A(n11331), .B(n11330), .Z(n11332) );
  XNOR U11620 ( .A(n11333), .B(n11332), .Z(n11142) );
  NANDN U11621 ( .A(n16746), .B(o[33]), .Z(n11140) );
  OR U11622 ( .A(n11021), .B(n11020), .Z(n11025) );
  OR U11623 ( .A(n11023), .B(n11022), .Z(n11024) );
  NAND U11624 ( .A(n11025), .B(n11024), .Z(n11141) );
  XOR U11625 ( .A(n11140), .B(n11141), .Z(n11143) );
  XNOR U11626 ( .A(n11142), .B(n11143), .Z(n11336) );
  XNOR U11627 ( .A(n11337), .B(n11336), .Z(n11338) );
  XNOR U11628 ( .A(n11339), .B(n11338), .Z(n11136) );
  NANDN U11629 ( .A(n16826), .B(o[35]), .Z(n11134) );
  OR U11630 ( .A(n11027), .B(n11026), .Z(n11031) );
  OR U11631 ( .A(n11029), .B(n11028), .Z(n11030) );
  NAND U11632 ( .A(n11031), .B(n11030), .Z(n11135) );
  XOR U11633 ( .A(n11134), .B(n11135), .Z(n11137) );
  XNOR U11634 ( .A(n11136), .B(n11137), .Z(n11342) );
  XNOR U11635 ( .A(n11343), .B(n11342), .Z(n11344) );
  XNOR U11636 ( .A(n11345), .B(n11344), .Z(n11130) );
  NANDN U11637 ( .A(n2976), .B(o[37]), .Z(n11128) );
  OR U11638 ( .A(n11033), .B(n11032), .Z(n11037) );
  OR U11639 ( .A(n11035), .B(n11034), .Z(n11036) );
  NAND U11640 ( .A(n11037), .B(n11036), .Z(n11129) );
  XOR U11641 ( .A(n11128), .B(n11129), .Z(n11131) );
  XNOR U11642 ( .A(n11130), .B(n11131), .Z(n11348) );
  XNOR U11643 ( .A(n11349), .B(n11348), .Z(n11350) );
  XNOR U11644 ( .A(n11351), .B(n11350), .Z(n11124) );
  NANDN U11645 ( .A(n2974), .B(o[39]), .Z(n11122) );
  OR U11646 ( .A(n11039), .B(n11038), .Z(n11043) );
  OR U11647 ( .A(n11041), .B(n11040), .Z(n11042) );
  NAND U11648 ( .A(n11043), .B(n11042), .Z(n11123) );
  XOR U11649 ( .A(n11122), .B(n11123), .Z(n11125) );
  XNOR U11650 ( .A(n11124), .B(n11125), .Z(n11354) );
  XNOR U11651 ( .A(n11355), .B(n11354), .Z(n11356) );
  XNOR U11652 ( .A(n11357), .B(n11356), .Z(n11118) );
  NANDN U11653 ( .A(n2972), .B(o[41]), .Z(n11116) );
  OR U11654 ( .A(n11045), .B(n11044), .Z(n11049) );
  OR U11655 ( .A(n11047), .B(n11046), .Z(n11048) );
  NAND U11656 ( .A(n11049), .B(n11048), .Z(n11117) );
  XOR U11657 ( .A(n11116), .B(n11117), .Z(n11119) );
  XNOR U11658 ( .A(n11118), .B(n11119), .Z(n11360) );
  XNOR U11659 ( .A(n11361), .B(n11360), .Z(n11362) );
  XNOR U11660 ( .A(n11363), .B(n11362), .Z(n11112) );
  NANDN U11661 ( .A(n17145), .B(o[43]), .Z(n11110) );
  OR U11662 ( .A(n11051), .B(n11050), .Z(n11055) );
  OR U11663 ( .A(n11053), .B(n11052), .Z(n11054) );
  NAND U11664 ( .A(n11055), .B(n11054), .Z(n11111) );
  XOR U11665 ( .A(n11110), .B(n11111), .Z(n11113) );
  XNOR U11666 ( .A(n11112), .B(n11113), .Z(n11366) );
  XNOR U11667 ( .A(n11367), .B(n11366), .Z(n11368) );
  XNOR U11668 ( .A(n11369), .B(n11368), .Z(n11106) );
  NANDN U11669 ( .A(n17219), .B(o[45]), .Z(n11104) );
  OR U11670 ( .A(n11057), .B(n11056), .Z(n11061) );
  OR U11671 ( .A(n11059), .B(n11058), .Z(n11060) );
  NAND U11672 ( .A(n11061), .B(n11060), .Z(n11105) );
  XOR U11673 ( .A(n11104), .B(n11105), .Z(n11107) );
  XNOR U11674 ( .A(n11106), .B(n11107), .Z(n11372) );
  XNOR U11675 ( .A(n11373), .B(n11372), .Z(n11374) );
  XNOR U11676 ( .A(n11375), .B(n11374), .Z(n11100) );
  NANDN U11677 ( .A(n17296), .B(o[47]), .Z(n11098) );
  OR U11678 ( .A(n11063), .B(n11062), .Z(n11067) );
  OR U11679 ( .A(n11065), .B(n11064), .Z(n11066) );
  NAND U11680 ( .A(n11067), .B(n11066), .Z(n11099) );
  XOR U11681 ( .A(n11098), .B(n11099), .Z(n11101) );
  XNOR U11682 ( .A(n11100), .B(n11101), .Z(n11378) );
  XNOR U11683 ( .A(n11379), .B(n11378), .Z(n11380) );
  XNOR U11684 ( .A(n11381), .B(n11380), .Z(n11094) );
  NANDN U11685 ( .A(n17375), .B(o[49]), .Z(n11092) );
  OR U11686 ( .A(n11069), .B(n11068), .Z(n11073) );
  OR U11687 ( .A(n11071), .B(n11070), .Z(n11072) );
  NAND U11688 ( .A(n11073), .B(n11072), .Z(n11093) );
  XOR U11689 ( .A(n11092), .B(n11093), .Z(n11095) );
  XNOR U11690 ( .A(n11094), .B(n11095), .Z(n11384) );
  XNOR U11691 ( .A(n11385), .B(n11384), .Z(n11386) );
  AND U11692 ( .A(o[51]), .B(\stack[1][1] ), .Z(n11086) );
  OR U11693 ( .A(n11075), .B(n11074), .Z(n11079) );
  OR U11694 ( .A(n11077), .B(n11076), .Z(n11078) );
  NAND U11695 ( .A(n11079), .B(n11078), .Z(n11087) );
  XNOR U11696 ( .A(n11086), .B(n11087), .Z(n11089) );
  XOR U11697 ( .A(n11088), .B(n11089), .Z(n11080) );
  NANDN U11698 ( .A(n11081), .B(n11080), .Z(n11083) );
  XOR U11699 ( .A(n11081), .B(n11080), .Z(n15471) );
  AND U11700 ( .A(o[52]), .B(\stack[1][0] ), .Z(n15472) );
  OR U11701 ( .A(n15471), .B(n15472), .Z(n11082) );
  AND U11702 ( .A(n11083), .B(n11082), .Z(n11085) );
  OR U11703 ( .A(n11084), .B(n11085), .Z(n11391) );
  XNOR U11704 ( .A(n11085), .B(n11084), .Z(n15432) );
  NANDN U11705 ( .A(n2969), .B(o[52]), .Z(n11699) );
  OR U11706 ( .A(n11087), .B(n11086), .Z(n11091) );
  OR U11707 ( .A(n11089), .B(n11088), .Z(n11090) );
  NAND U11708 ( .A(n11091), .B(n11090), .Z(n11697) );
  NANDN U11709 ( .A(n17375), .B(o[50]), .Z(n11693) );
  NANDN U11710 ( .A(n11093), .B(n11092), .Z(n11097) );
  NANDN U11711 ( .A(n11095), .B(n11094), .Z(n11096) );
  NAND U11712 ( .A(n11097), .B(n11096), .Z(n11691) );
  NANDN U11713 ( .A(n17296), .B(o[48]), .Z(n11687) );
  NANDN U11714 ( .A(n11099), .B(n11098), .Z(n11103) );
  NANDN U11715 ( .A(n11101), .B(n11100), .Z(n11102) );
  NAND U11716 ( .A(n11103), .B(n11102), .Z(n11685) );
  NANDN U11717 ( .A(n17219), .B(o[46]), .Z(n11681) );
  NANDN U11718 ( .A(n11105), .B(n11104), .Z(n11109) );
  NANDN U11719 ( .A(n11107), .B(n11106), .Z(n11108) );
  NAND U11720 ( .A(n11109), .B(n11108), .Z(n11679) );
  NANDN U11721 ( .A(n17145), .B(o[44]), .Z(n11675) );
  NANDN U11722 ( .A(n11111), .B(n11110), .Z(n11115) );
  NANDN U11723 ( .A(n11113), .B(n11112), .Z(n11114) );
  NAND U11724 ( .A(n11115), .B(n11114), .Z(n11673) );
  NANDN U11725 ( .A(n2972), .B(o[42]), .Z(n11669) );
  NANDN U11726 ( .A(n11117), .B(n11116), .Z(n11121) );
  NANDN U11727 ( .A(n11119), .B(n11118), .Z(n11120) );
  NAND U11728 ( .A(n11121), .B(n11120), .Z(n11667) );
  NANDN U11729 ( .A(n2974), .B(o[40]), .Z(n11663) );
  NANDN U11730 ( .A(n11123), .B(n11122), .Z(n11127) );
  NANDN U11731 ( .A(n11125), .B(n11124), .Z(n11126) );
  NAND U11732 ( .A(n11127), .B(n11126), .Z(n11661) );
  NANDN U11733 ( .A(n2976), .B(o[38]), .Z(n11657) );
  NANDN U11734 ( .A(n11129), .B(n11128), .Z(n11133) );
  NANDN U11735 ( .A(n11131), .B(n11130), .Z(n11132) );
  NAND U11736 ( .A(n11133), .B(n11132), .Z(n11655) );
  NANDN U11737 ( .A(n16826), .B(o[36]), .Z(n11651) );
  NANDN U11738 ( .A(n11135), .B(n11134), .Z(n11139) );
  NANDN U11739 ( .A(n11137), .B(n11136), .Z(n11138) );
  NAND U11740 ( .A(n11139), .B(n11138), .Z(n11649) );
  NANDN U11741 ( .A(n16746), .B(o[34]), .Z(n11645) );
  NANDN U11742 ( .A(n11141), .B(n11140), .Z(n11145) );
  NANDN U11743 ( .A(n11143), .B(n11142), .Z(n11144) );
  NAND U11744 ( .A(n11145), .B(n11144), .Z(n11643) );
  NANDN U11745 ( .A(n2978), .B(o[32]), .Z(n11639) );
  NANDN U11746 ( .A(n11147), .B(n11146), .Z(n11151) );
  NANDN U11747 ( .A(n11149), .B(n11148), .Z(n11150) );
  NAND U11748 ( .A(n11151), .B(n11150), .Z(n11637) );
  NANDN U11749 ( .A(n2980), .B(o[30]), .Z(n11633) );
  NANDN U11750 ( .A(n11153), .B(n11152), .Z(n11157) );
  NANDN U11751 ( .A(n11155), .B(n11154), .Z(n11156) );
  NAND U11752 ( .A(n11157), .B(n11156), .Z(n11631) );
  NANDN U11753 ( .A(n2982), .B(o[28]), .Z(n11627) );
  NANDN U11754 ( .A(n11159), .B(n11158), .Z(n11163) );
  NANDN U11755 ( .A(n11161), .B(n11160), .Z(n11162) );
  NAND U11756 ( .A(n11163), .B(n11162), .Z(n11625) );
  NANDN U11757 ( .A(n3020), .B(\stack[1][27] ), .Z(n11621) );
  NANDN U11758 ( .A(n11165), .B(n11164), .Z(n11169) );
  NANDN U11759 ( .A(n11167), .B(n11166), .Z(n11168) );
  NAND U11760 ( .A(n11169), .B(n11168), .Z(n11619) );
  NANDN U11761 ( .A(n3018), .B(\stack[1][29] ), .Z(n11615) );
  NANDN U11762 ( .A(n11171), .B(n11170), .Z(n11175) );
  NANDN U11763 ( .A(n11173), .B(n11172), .Z(n11174) );
  NAND U11764 ( .A(n11175), .B(n11174), .Z(n11613) );
  NANDN U11765 ( .A(n3016), .B(\stack[1][31] ), .Z(n11609) );
  NANDN U11766 ( .A(n11177), .B(n11176), .Z(n11181) );
  NANDN U11767 ( .A(n11179), .B(n11178), .Z(n11180) );
  NAND U11768 ( .A(n11181), .B(n11180), .Z(n11607) );
  AND U11769 ( .A(\stack[1][33] ), .B(o[20]), .Z(n11603) );
  NANDN U11770 ( .A(n11183), .B(n11182), .Z(n11187) );
  NANDN U11771 ( .A(n11185), .B(n11184), .Z(n11186) );
  AND U11772 ( .A(n11187), .B(n11186), .Z(n11600) );
  AND U11773 ( .A(\stack[1][34] ), .B(o[19]), .Z(n11488) );
  OR U11774 ( .A(n11189), .B(n11188), .Z(n11193) );
  OR U11775 ( .A(n11191), .B(n11190), .Z(n11192) );
  NAND U11776 ( .A(n11193), .B(n11192), .Z(n11489) );
  XNOR U11777 ( .A(n11488), .B(n11489), .Z(n11491) );
  OR U11778 ( .A(n11195), .B(n11194), .Z(n11199) );
  NANDN U11779 ( .A(n11197), .B(n11196), .Z(n11198) );
  NAND U11780 ( .A(n11199), .B(n11198), .Z(n11495) );
  ANDN U11781 ( .B(o[17]), .A(n2993), .Z(n11494) );
  XOR U11782 ( .A(n11495), .B(n11494), .Z(n11496) );
  NANDN U11783 ( .A(n3010), .B(\stack[1][37] ), .Z(n11503) );
  OR U11784 ( .A(n11201), .B(n11200), .Z(n11205) );
  NANDN U11785 ( .A(n11203), .B(n11202), .Z(n11204) );
  NAND U11786 ( .A(n11205), .B(n11204), .Z(n11501) );
  ANDN U11787 ( .B(\stack[1][38] ), .A(n3009), .Z(n11509) );
  NANDN U11788 ( .A(n11207), .B(n11206), .Z(n11211) );
  NANDN U11789 ( .A(n11209), .B(n11208), .Z(n11210) );
  AND U11790 ( .A(n11211), .B(n11210), .Z(n11506) );
  NAND U11791 ( .A(n11213), .B(n11212), .Z(n11217) );
  OR U11792 ( .A(n11215), .B(n11214), .Z(n11216) );
  AND U11793 ( .A(n11217), .B(n11216), .Z(n11585) );
  OR U11794 ( .A(n11219), .B(n11218), .Z(n11223) );
  NANDN U11795 ( .A(n11221), .B(n11220), .Z(n11222) );
  NAND U11796 ( .A(n11223), .B(n11222), .Z(n11515) );
  AND U11797 ( .A(\stack[1][42] ), .B(o[11]), .Z(n11521) );
  OR U11798 ( .A(n11225), .B(n11224), .Z(n11229) );
  NANDN U11799 ( .A(n11227), .B(n11226), .Z(n11228) );
  AND U11800 ( .A(n11229), .B(n11228), .Z(n11518) );
  AND U11801 ( .A(\stack[1][43] ), .B(o[10]), .Z(n11527) );
  AND U11802 ( .A(\stack[1][44] ), .B(o[9]), .Z(n11578) );
  NANDN U11803 ( .A(n11231), .B(n11230), .Z(n11235) );
  NAND U11804 ( .A(n11233), .B(n11232), .Z(n11234) );
  AND U11805 ( .A(n11235), .B(n11234), .Z(n11567) );
  AND U11806 ( .A(\stack[1][48] ), .B(o[5]), .Z(n11561) );
  OR U11807 ( .A(n11237), .B(n11236), .Z(n11241) );
  NANDN U11808 ( .A(n11239), .B(n11238), .Z(n11240) );
  AND U11809 ( .A(n11241), .B(n11240), .Z(n11558) );
  ANDN U11810 ( .B(\stack[1][49] ), .A(n2998), .Z(n11539) );
  AND U11811 ( .A(\stack[1][50] ), .B(o[3]), .Z(n11555) );
  NANDN U11812 ( .A(n11242), .B(n11542), .Z(n11243) );
  AND U11813 ( .A(n11244), .B(n11243), .Z(n11248) );
  OR U11814 ( .A(n11246), .B(n11245), .Z(n11247) );
  AND U11815 ( .A(n11248), .B(n11247), .Z(n11552) );
  AND U11816 ( .A(\stack[1][53] ), .B(o[1]), .Z(n11550) );
  ANDN U11817 ( .B(n11550), .A(n11249), .Z(n11863) );
  XNOR U11818 ( .A(n11863), .B(n11542), .Z(n11251) );
  NAND U11819 ( .A(o[0]), .B(\stack[1][53] ), .Z(n11549) );
  NANDN U11820 ( .A(n11250), .B(n11549), .Z(n11544) );
  NAND U11821 ( .A(n11251), .B(n11544), .Z(n11546) );
  AND U11822 ( .A(\stack[1][51] ), .B(o[2]), .Z(n11545) );
  XNOR U11823 ( .A(n11546), .B(n11545), .Z(n11553) );
  XOR U11824 ( .A(n11552), .B(n11553), .Z(n11554) );
  XOR U11825 ( .A(n11555), .B(n11554), .Z(n11537) );
  OR U11826 ( .A(n11253), .B(n11252), .Z(n11257) );
  NANDN U11827 ( .A(n11255), .B(n11254), .Z(n11256) );
  AND U11828 ( .A(n11257), .B(n11256), .Z(n11536) );
  XOR U11829 ( .A(n11537), .B(n11536), .Z(n11538) );
  XOR U11830 ( .A(n11539), .B(n11538), .Z(n11559) );
  XNOR U11831 ( .A(n11558), .B(n11559), .Z(n11560) );
  OR U11832 ( .A(n11259), .B(n11258), .Z(n11263) );
  OR U11833 ( .A(n11261), .B(n11260), .Z(n11262) );
  NAND U11834 ( .A(n11263), .B(n11262), .Z(n11531) );
  IV U11835 ( .A(\stack[1][47] ), .Z(n15662) );
  ANDN U11836 ( .B(o[6]), .A(n15662), .Z(n11530) );
  XNOR U11837 ( .A(n11531), .B(n11530), .Z(n11533) );
  XNOR U11838 ( .A(n11532), .B(n11533), .Z(n11565) );
  ANDN U11839 ( .B(o[7]), .A(n15701), .Z(n11564) );
  XOR U11840 ( .A(n11565), .B(n11564), .Z(n11566) );
  NANDN U11841 ( .A(n11265), .B(n11264), .Z(n11269) );
  OR U11842 ( .A(n11267), .B(n11266), .Z(n11268) );
  AND U11843 ( .A(n11269), .B(n11268), .Z(n11570) );
  XNOR U11844 ( .A(n11571), .B(n11570), .Z(n11573) );
  AND U11845 ( .A(\stack[1][45] ), .B(o[8]), .Z(n11572) );
  XNOR U11846 ( .A(n11573), .B(n11572), .Z(n11576) );
  OR U11847 ( .A(n11271), .B(n11270), .Z(n11275) );
  NANDN U11848 ( .A(n11273), .B(n11272), .Z(n11274) );
  NAND U11849 ( .A(n11275), .B(n11274), .Z(n11577) );
  XNOR U11850 ( .A(n11576), .B(n11577), .Z(n11579) );
  XNOR U11851 ( .A(n11578), .B(n11579), .Z(n11525) );
  OR U11852 ( .A(n11277), .B(n11276), .Z(n11281) );
  OR U11853 ( .A(n11279), .B(n11278), .Z(n11280) );
  AND U11854 ( .A(n11281), .B(n11280), .Z(n11524) );
  XOR U11855 ( .A(n11525), .B(n11524), .Z(n11526) );
  XOR U11856 ( .A(n11527), .B(n11526), .Z(n11519) );
  XOR U11857 ( .A(n11518), .B(n11519), .Z(n11520) );
  XOR U11858 ( .A(n11521), .B(n11520), .Z(n11513) );
  AND U11859 ( .A(\stack[1][41] ), .B(o[12]), .Z(n11512) );
  XNOR U11860 ( .A(n11513), .B(n11512), .Z(n11514) );
  XNOR U11861 ( .A(n11515), .B(n11514), .Z(n11583) );
  ANDN U11862 ( .B(o[13]), .A(n15935), .Z(n11582) );
  XOR U11863 ( .A(n11583), .B(n11582), .Z(n11584) );
  NANDN U11864 ( .A(n11283), .B(n11282), .Z(n11287) );
  OR U11865 ( .A(n11285), .B(n11284), .Z(n11286) );
  AND U11866 ( .A(n11287), .B(n11286), .Z(n11588) );
  XNOR U11867 ( .A(n11589), .B(n11588), .Z(n11591) );
  NANDN U11868 ( .A(n3008), .B(\stack[1][39] ), .Z(n11590) );
  XOR U11869 ( .A(n11591), .B(n11590), .Z(n11507) );
  XNOR U11870 ( .A(n11506), .B(n11507), .Z(n11508) );
  XOR U11871 ( .A(n11501), .B(n11500), .Z(n11502) );
  XNOR U11872 ( .A(n11503), .B(n11502), .Z(n11497) );
  OR U11873 ( .A(n11289), .B(n11288), .Z(n11293) );
  OR U11874 ( .A(n11291), .B(n11290), .Z(n11292) );
  AND U11875 ( .A(n11293), .B(n11292), .Z(n11595) );
  XNOR U11876 ( .A(n11594), .B(n11595), .Z(n11597) );
  AND U11877 ( .A(\stack[1][35] ), .B(o[18]), .Z(n11596) );
  XOR U11878 ( .A(n11597), .B(n11596), .Z(n11490) );
  XOR U11879 ( .A(n11491), .B(n11490), .Z(n11601) );
  XOR U11880 ( .A(n11600), .B(n11601), .Z(n11602) );
  XOR U11881 ( .A(n11603), .B(n11602), .Z(n11485) );
  AND U11882 ( .A(\stack[1][32] ), .B(o[21]), .Z(n11482) );
  OR U11883 ( .A(n11295), .B(n11294), .Z(n11299) );
  OR U11884 ( .A(n11297), .B(n11296), .Z(n11298) );
  NAND U11885 ( .A(n11299), .B(n11298), .Z(n11483) );
  XNOR U11886 ( .A(n11482), .B(n11483), .Z(n11484) );
  XOR U11887 ( .A(n11485), .B(n11484), .Z(n11606) );
  XNOR U11888 ( .A(n11607), .B(n11606), .Z(n11608) );
  XNOR U11889 ( .A(n11609), .B(n11608), .Z(n11478) );
  NANDN U11890 ( .A(n2987), .B(o[23]), .Z(n11476) );
  OR U11891 ( .A(n11301), .B(n11300), .Z(n11305) );
  OR U11892 ( .A(n11303), .B(n11302), .Z(n11304) );
  NAND U11893 ( .A(n11305), .B(n11304), .Z(n11477) );
  XOR U11894 ( .A(n11476), .B(n11477), .Z(n11479) );
  XNOR U11895 ( .A(n11478), .B(n11479), .Z(n11612) );
  XNOR U11896 ( .A(n11613), .B(n11612), .Z(n11614) );
  XNOR U11897 ( .A(n11615), .B(n11614), .Z(n11472) );
  NANDN U11898 ( .A(n2985), .B(o[25]), .Z(n11470) );
  OR U11899 ( .A(n11307), .B(n11306), .Z(n11311) );
  OR U11900 ( .A(n11309), .B(n11308), .Z(n11310) );
  NAND U11901 ( .A(n11311), .B(n11310), .Z(n11471) );
  XOR U11902 ( .A(n11470), .B(n11471), .Z(n11473) );
  XNOR U11903 ( .A(n11472), .B(n11473), .Z(n11618) );
  XNOR U11904 ( .A(n11619), .B(n11618), .Z(n11620) );
  XNOR U11905 ( .A(n11621), .B(n11620), .Z(n11466) );
  NANDN U11906 ( .A(n2983), .B(o[27]), .Z(n11464) );
  OR U11907 ( .A(n11313), .B(n11312), .Z(n11317) );
  IV U11908 ( .A(n11314), .Z(n16472) );
  OR U11909 ( .A(n11315), .B(n16472), .Z(n11316) );
  NAND U11910 ( .A(n11317), .B(n11316), .Z(n11465) );
  XOR U11911 ( .A(n11464), .B(n11465), .Z(n11467) );
  XNOR U11912 ( .A(n11466), .B(n11467), .Z(n11624) );
  XNOR U11913 ( .A(n11625), .B(n11624), .Z(n11626) );
  XNOR U11914 ( .A(n11627), .B(n11626), .Z(n11460) );
  NANDN U11915 ( .A(n2981), .B(o[29]), .Z(n11458) );
  OR U11916 ( .A(n11319), .B(n11318), .Z(n11323) );
  OR U11917 ( .A(n11321), .B(n11320), .Z(n11322) );
  NAND U11918 ( .A(n11323), .B(n11322), .Z(n11459) );
  XOR U11919 ( .A(n11458), .B(n11459), .Z(n11461) );
  XNOR U11920 ( .A(n11460), .B(n11461), .Z(n11630) );
  XNOR U11921 ( .A(n11631), .B(n11630), .Z(n11632) );
  XNOR U11922 ( .A(n11633), .B(n11632), .Z(n11454) );
  NANDN U11923 ( .A(n2979), .B(o[31]), .Z(n11452) );
  OR U11924 ( .A(n11325), .B(n11324), .Z(n11329) );
  OR U11925 ( .A(n11327), .B(n11326), .Z(n11328) );
  NAND U11926 ( .A(n11329), .B(n11328), .Z(n11453) );
  XOR U11927 ( .A(n11452), .B(n11453), .Z(n11455) );
  XNOR U11928 ( .A(n11454), .B(n11455), .Z(n11636) );
  XNOR U11929 ( .A(n11637), .B(n11636), .Z(n11638) );
  XNOR U11930 ( .A(n11639), .B(n11638), .Z(n11448) );
  NANDN U11931 ( .A(n16712), .B(o[33]), .Z(n11446) );
  OR U11932 ( .A(n11331), .B(n11330), .Z(n11335) );
  OR U11933 ( .A(n11333), .B(n11332), .Z(n11334) );
  NAND U11934 ( .A(n11335), .B(n11334), .Z(n11447) );
  XOR U11935 ( .A(n11446), .B(n11447), .Z(n11449) );
  XNOR U11936 ( .A(n11448), .B(n11449), .Z(n11642) );
  XNOR U11937 ( .A(n11643), .B(n11642), .Z(n11644) );
  XNOR U11938 ( .A(n11645), .B(n11644), .Z(n11442) );
  NANDN U11939 ( .A(n16786), .B(o[35]), .Z(n11440) );
  OR U11940 ( .A(n11337), .B(n11336), .Z(n11341) );
  OR U11941 ( .A(n11339), .B(n11338), .Z(n11340) );
  NAND U11942 ( .A(n11341), .B(n11340), .Z(n11441) );
  XOR U11943 ( .A(n11440), .B(n11441), .Z(n11443) );
  XNOR U11944 ( .A(n11442), .B(n11443), .Z(n11648) );
  XNOR U11945 ( .A(n11649), .B(n11648), .Z(n11650) );
  XNOR U11946 ( .A(n11651), .B(n11650), .Z(n11436) );
  NANDN U11947 ( .A(n2977), .B(o[37]), .Z(n11434) );
  OR U11948 ( .A(n11343), .B(n11342), .Z(n11347) );
  OR U11949 ( .A(n11345), .B(n11344), .Z(n11346) );
  NAND U11950 ( .A(n11347), .B(n11346), .Z(n11435) );
  XOR U11951 ( .A(n11434), .B(n11435), .Z(n11437) );
  XNOR U11952 ( .A(n11436), .B(n11437), .Z(n11654) );
  XNOR U11953 ( .A(n11655), .B(n11654), .Z(n11656) );
  XNOR U11954 ( .A(n11657), .B(n11656), .Z(n11430) );
  NANDN U11955 ( .A(n2975), .B(o[39]), .Z(n11428) );
  OR U11956 ( .A(n11349), .B(n11348), .Z(n11353) );
  OR U11957 ( .A(n11351), .B(n11350), .Z(n11352) );
  NAND U11958 ( .A(n11353), .B(n11352), .Z(n11429) );
  XOR U11959 ( .A(n11428), .B(n11429), .Z(n11431) );
  XNOR U11960 ( .A(n11430), .B(n11431), .Z(n11660) );
  XNOR U11961 ( .A(n11661), .B(n11660), .Z(n11662) );
  XNOR U11962 ( .A(n11663), .B(n11662), .Z(n11424) );
  NANDN U11963 ( .A(n2973), .B(o[41]), .Z(n11422) );
  OR U11964 ( .A(n11355), .B(n11354), .Z(n11359) );
  OR U11965 ( .A(n11357), .B(n11356), .Z(n11358) );
  NAND U11966 ( .A(n11359), .B(n11358), .Z(n11423) );
  XOR U11967 ( .A(n11422), .B(n11423), .Z(n11425) );
  XNOR U11968 ( .A(n11424), .B(n11425), .Z(n11666) );
  XNOR U11969 ( .A(n11667), .B(n11666), .Z(n11668) );
  XNOR U11970 ( .A(n11669), .B(n11668), .Z(n11418) );
  NANDN U11971 ( .A(n17101), .B(o[43]), .Z(n11416) );
  OR U11972 ( .A(n11361), .B(n11360), .Z(n11365) );
  OR U11973 ( .A(n11363), .B(n11362), .Z(n11364) );
  NAND U11974 ( .A(n11365), .B(n11364), .Z(n11417) );
  XOR U11975 ( .A(n11416), .B(n11417), .Z(n11419) );
  XNOR U11976 ( .A(n11418), .B(n11419), .Z(n11672) );
  XNOR U11977 ( .A(n11673), .B(n11672), .Z(n11674) );
  XNOR U11978 ( .A(n11675), .B(n11674), .Z(n11412) );
  NANDN U11979 ( .A(n17179), .B(o[45]), .Z(n11410) );
  OR U11980 ( .A(n11367), .B(n11366), .Z(n11371) );
  OR U11981 ( .A(n11369), .B(n11368), .Z(n11370) );
  NAND U11982 ( .A(n11371), .B(n11370), .Z(n11411) );
  XOR U11983 ( .A(n11410), .B(n11411), .Z(n11413) );
  XNOR U11984 ( .A(n11412), .B(n11413), .Z(n11678) );
  XNOR U11985 ( .A(n11679), .B(n11678), .Z(n11680) );
  XNOR U11986 ( .A(n11681), .B(n11680), .Z(n11406) );
  NANDN U11987 ( .A(n17256), .B(o[47]), .Z(n11404) );
  OR U11988 ( .A(n11373), .B(n11372), .Z(n11377) );
  OR U11989 ( .A(n11375), .B(n11374), .Z(n11376) );
  NAND U11990 ( .A(n11377), .B(n11376), .Z(n11405) );
  XOR U11991 ( .A(n11404), .B(n11405), .Z(n11407) );
  XNOR U11992 ( .A(n11406), .B(n11407), .Z(n11684) );
  XNOR U11993 ( .A(n11685), .B(n11684), .Z(n11686) );
  XNOR U11994 ( .A(n11687), .B(n11686), .Z(n11400) );
  AND U11995 ( .A(o[49]), .B(\stack[1][4] ), .Z(n11398) );
  OR U11996 ( .A(n11379), .B(n11378), .Z(n11383) );
  OR U11997 ( .A(n11381), .B(n11380), .Z(n11382) );
  NAND U11998 ( .A(n11383), .B(n11382), .Z(n11399) );
  XNOR U11999 ( .A(n11398), .B(n11399), .Z(n11401) );
  XNOR U12000 ( .A(n11400), .B(n11401), .Z(n11690) );
  XNOR U12001 ( .A(n11691), .B(n11690), .Z(n11692) );
  XOR U12002 ( .A(n11693), .B(n11692), .Z(n11395) );
  AND U12003 ( .A(o[51]), .B(\stack[1][2] ), .Z(n11392) );
  OR U12004 ( .A(n11385), .B(n11384), .Z(n11389) );
  OR U12005 ( .A(n11387), .B(n11386), .Z(n11388) );
  NAND U12006 ( .A(n11389), .B(n11388), .Z(n11393) );
  XOR U12007 ( .A(n11392), .B(n11393), .Z(n11394) );
  XNOR U12008 ( .A(n11395), .B(n11394), .Z(n11696) );
  XNOR U12009 ( .A(n11697), .B(n11696), .Z(n11698) );
  XOR U12010 ( .A(n11699), .B(n11698), .Z(n15433) );
  OR U12011 ( .A(n15432), .B(n15433), .Z(n11390) );
  AND U12012 ( .A(n11391), .B(n11390), .Z(n11703) );
  NANDN U12013 ( .A(n2970), .B(o[52]), .Z(n12020) );
  OR U12014 ( .A(n11393), .B(n11392), .Z(n11397) );
  NANDN U12015 ( .A(n11395), .B(n11394), .Z(n11396) );
  NAND U12016 ( .A(n11397), .B(n11396), .Z(n12018) );
  NANDN U12017 ( .A(n2971), .B(o[50]), .Z(n12014) );
  OR U12018 ( .A(n11399), .B(n11398), .Z(n11403) );
  NANDN U12019 ( .A(n11401), .B(n11400), .Z(n11402) );
  NAND U12020 ( .A(n11403), .B(n11402), .Z(n12012) );
  NANDN U12021 ( .A(n17256), .B(o[48]), .Z(n12008) );
  NANDN U12022 ( .A(n11405), .B(n11404), .Z(n11409) );
  NANDN U12023 ( .A(n11407), .B(n11406), .Z(n11408) );
  NAND U12024 ( .A(n11409), .B(n11408), .Z(n12006) );
  NANDN U12025 ( .A(n17179), .B(o[46]), .Z(n12002) );
  NANDN U12026 ( .A(n11411), .B(n11410), .Z(n11415) );
  NANDN U12027 ( .A(n11413), .B(n11412), .Z(n11414) );
  NAND U12028 ( .A(n11415), .B(n11414), .Z(n12000) );
  NANDN U12029 ( .A(n17101), .B(o[44]), .Z(n11996) );
  NANDN U12030 ( .A(n11417), .B(n11416), .Z(n11421) );
  NANDN U12031 ( .A(n11419), .B(n11418), .Z(n11420) );
  NAND U12032 ( .A(n11421), .B(n11420), .Z(n11994) );
  NANDN U12033 ( .A(n2973), .B(o[42]), .Z(n11990) );
  NANDN U12034 ( .A(n11423), .B(n11422), .Z(n11427) );
  NANDN U12035 ( .A(n11425), .B(n11424), .Z(n11426) );
  NAND U12036 ( .A(n11427), .B(n11426), .Z(n11988) );
  NANDN U12037 ( .A(n2975), .B(o[40]), .Z(n11984) );
  NANDN U12038 ( .A(n11429), .B(n11428), .Z(n11433) );
  NANDN U12039 ( .A(n11431), .B(n11430), .Z(n11432) );
  NAND U12040 ( .A(n11433), .B(n11432), .Z(n11982) );
  NANDN U12041 ( .A(n2977), .B(o[38]), .Z(n11978) );
  NANDN U12042 ( .A(n11435), .B(n11434), .Z(n11439) );
  NANDN U12043 ( .A(n11437), .B(n11436), .Z(n11438) );
  NAND U12044 ( .A(n11439), .B(n11438), .Z(n11976) );
  NANDN U12045 ( .A(n16786), .B(o[36]), .Z(n11972) );
  NANDN U12046 ( .A(n11441), .B(n11440), .Z(n11445) );
  NANDN U12047 ( .A(n11443), .B(n11442), .Z(n11444) );
  NAND U12048 ( .A(n11445), .B(n11444), .Z(n11970) );
  NANDN U12049 ( .A(n16712), .B(o[34]), .Z(n11966) );
  NANDN U12050 ( .A(n11447), .B(n11446), .Z(n11451) );
  NANDN U12051 ( .A(n11449), .B(n11448), .Z(n11450) );
  NAND U12052 ( .A(n11451), .B(n11450), .Z(n11964) );
  NANDN U12053 ( .A(n2979), .B(o[32]), .Z(n11960) );
  NANDN U12054 ( .A(n11453), .B(n11452), .Z(n11457) );
  NANDN U12055 ( .A(n11455), .B(n11454), .Z(n11456) );
  NAND U12056 ( .A(n11457), .B(n11456), .Z(n11958) );
  NANDN U12057 ( .A(n2981), .B(o[30]), .Z(n11954) );
  NANDN U12058 ( .A(n11459), .B(n11458), .Z(n11463) );
  NANDN U12059 ( .A(n11461), .B(n11460), .Z(n11462) );
  NAND U12060 ( .A(n11463), .B(n11462), .Z(n11952) );
  NANDN U12061 ( .A(n2983), .B(o[28]), .Z(n11948) );
  NANDN U12062 ( .A(n11465), .B(n11464), .Z(n11469) );
  NANDN U12063 ( .A(n11467), .B(n11466), .Z(n11468) );
  NAND U12064 ( .A(n11469), .B(n11468), .Z(n11946) );
  NANDN U12065 ( .A(n3020), .B(\stack[1][28] ), .Z(n11942) );
  NANDN U12066 ( .A(n11471), .B(n11470), .Z(n11475) );
  NANDN U12067 ( .A(n11473), .B(n11472), .Z(n11474) );
  NAND U12068 ( .A(n11475), .B(n11474), .Z(n11940) );
  NANDN U12069 ( .A(n3018), .B(\stack[1][30] ), .Z(n11936) );
  NANDN U12070 ( .A(n11477), .B(n11476), .Z(n11481) );
  NANDN U12071 ( .A(n11479), .B(n11478), .Z(n11480) );
  NAND U12072 ( .A(n11481), .B(n11480), .Z(n11934) );
  NANDN U12073 ( .A(n3016), .B(\stack[1][32] ), .Z(n11930) );
  OR U12074 ( .A(n11483), .B(n11482), .Z(n11487) );
  OR U12075 ( .A(n11485), .B(n11484), .Z(n11486) );
  NAND U12076 ( .A(n11487), .B(n11486), .Z(n11928) );
  NANDN U12077 ( .A(n3014), .B(\stack[1][34] ), .Z(n11812) );
  OR U12078 ( .A(n11489), .B(n11488), .Z(n11493) );
  NANDN U12079 ( .A(n11491), .B(n11490), .Z(n11492) );
  NAND U12080 ( .A(n11493), .B(n11492), .Z(n11810) );
  NANDN U12081 ( .A(n11495), .B(n11494), .Z(n11499) );
  OR U12082 ( .A(n11497), .B(n11496), .Z(n11498) );
  AND U12083 ( .A(n11499), .B(n11498), .Z(n11815) );
  AND U12084 ( .A(\stack[1][37] ), .B(o[17]), .Z(n11821) );
  NANDN U12085 ( .A(n11501), .B(n11500), .Z(n11505) );
  OR U12086 ( .A(n11503), .B(n11502), .Z(n11504) );
  NAND U12087 ( .A(n11505), .B(n11504), .Z(n11822) );
  XNOR U12088 ( .A(n11821), .B(n11822), .Z(n11824) );
  ANDN U12089 ( .B(\stack[1][38] ), .A(n3010), .Z(n11830) );
  OR U12090 ( .A(n11507), .B(n11506), .Z(n11511) );
  OR U12091 ( .A(n11509), .B(n11508), .Z(n11510) );
  AND U12092 ( .A(n11511), .B(n11510), .Z(n11827) );
  NANDN U12093 ( .A(n3009), .B(\stack[1][39] ), .Z(n11836) );
  NAND U12094 ( .A(n11513), .B(n11512), .Z(n11517) );
  OR U12095 ( .A(n11515), .B(n11514), .Z(n11516) );
  AND U12096 ( .A(n11517), .B(n11516), .Z(n11912) );
  OR U12097 ( .A(n11519), .B(n11518), .Z(n11523) );
  NANDN U12098 ( .A(n11521), .B(n11520), .Z(n11522) );
  NAND U12099 ( .A(n11523), .B(n11522), .Z(n11842) );
  NANDN U12100 ( .A(n3006), .B(\stack[1][42] ), .Z(n11840) );
  NANDN U12101 ( .A(n15818), .B(o[11]), .Z(n11905) );
  OR U12102 ( .A(n11525), .B(n11524), .Z(n11529) );
  NANDN U12103 ( .A(n11527), .B(n11526), .Z(n11528) );
  AND U12104 ( .A(n11529), .B(n11528), .Z(n11904) );
  NANDN U12105 ( .A(n15779), .B(o[10]), .Z(n11847) );
  AND U12106 ( .A(\stack[1][45] ), .B(o[9]), .Z(n11899) );
  NANDN U12107 ( .A(n11531), .B(n11530), .Z(n11535) );
  NAND U12108 ( .A(n11533), .B(n11532), .Z(n11534) );
  AND U12109 ( .A(n11535), .B(n11534), .Z(n11888) );
  ANDN U12110 ( .B(\stack[1][49] ), .A(n2999), .Z(n11882) );
  OR U12111 ( .A(n11537), .B(n11536), .Z(n11541) );
  NANDN U12112 ( .A(n11539), .B(n11538), .Z(n11540) );
  AND U12113 ( .A(n11541), .B(n11540), .Z(n11879) );
  AND U12114 ( .A(\stack[1][50] ), .B(o[4]), .Z(n11860) );
  AND U12115 ( .A(\stack[1][51] ), .B(o[3]), .Z(n11876) );
  NANDN U12116 ( .A(n11542), .B(n11863), .Z(n11543) );
  AND U12117 ( .A(n11544), .B(n11543), .Z(n11548) );
  OR U12118 ( .A(n11546), .B(n11545), .Z(n11547) );
  AND U12119 ( .A(n11548), .B(n11547), .Z(n11873) );
  AND U12120 ( .A(\stack[1][54] ), .B(o[1]), .Z(n11871) );
  ANDN U12121 ( .B(n11871), .A(n11549), .Z(n12193) );
  XNOR U12122 ( .A(n12193), .B(n11863), .Z(n11551) );
  NAND U12123 ( .A(o[0]), .B(\stack[1][54] ), .Z(n11870) );
  NANDN U12124 ( .A(n11550), .B(n11870), .Z(n11865) );
  NAND U12125 ( .A(n11551), .B(n11865), .Z(n11867) );
  AND U12126 ( .A(\stack[1][52] ), .B(o[2]), .Z(n11866) );
  XNOR U12127 ( .A(n11867), .B(n11866), .Z(n11874) );
  XOR U12128 ( .A(n11873), .B(n11874), .Z(n11875) );
  XOR U12129 ( .A(n11876), .B(n11875), .Z(n11858) );
  OR U12130 ( .A(n11553), .B(n11552), .Z(n11557) );
  NANDN U12131 ( .A(n11555), .B(n11554), .Z(n11556) );
  AND U12132 ( .A(n11557), .B(n11556), .Z(n11857) );
  XOR U12133 ( .A(n11858), .B(n11857), .Z(n11859) );
  XOR U12134 ( .A(n11860), .B(n11859), .Z(n11880) );
  XNOR U12135 ( .A(n11879), .B(n11880), .Z(n11881) );
  OR U12136 ( .A(n11559), .B(n11558), .Z(n11563) );
  OR U12137 ( .A(n11561), .B(n11560), .Z(n11562) );
  NAND U12138 ( .A(n11563), .B(n11562), .Z(n11852) );
  IV U12139 ( .A(\stack[1][48] ), .Z(n15623) );
  ANDN U12140 ( .B(o[6]), .A(n15623), .Z(n11851) );
  XNOR U12141 ( .A(n11852), .B(n11851), .Z(n11854) );
  XNOR U12142 ( .A(n11853), .B(n11854), .Z(n11886) );
  ANDN U12143 ( .B(o[7]), .A(n15662), .Z(n11885) );
  XOR U12144 ( .A(n11886), .B(n11885), .Z(n11887) );
  NANDN U12145 ( .A(n11565), .B(n11564), .Z(n11569) );
  OR U12146 ( .A(n11567), .B(n11566), .Z(n11568) );
  AND U12147 ( .A(n11569), .B(n11568), .Z(n11891) );
  XNOR U12148 ( .A(n11892), .B(n11891), .Z(n11894) );
  AND U12149 ( .A(\stack[1][46] ), .B(o[8]), .Z(n11893) );
  XNOR U12150 ( .A(n11894), .B(n11893), .Z(n11897) );
  OR U12151 ( .A(n11571), .B(n11570), .Z(n11575) );
  NANDN U12152 ( .A(n11573), .B(n11572), .Z(n11574) );
  NAND U12153 ( .A(n11575), .B(n11574), .Z(n11898) );
  XNOR U12154 ( .A(n11897), .B(n11898), .Z(n11900) );
  XNOR U12155 ( .A(n11899), .B(n11900), .Z(n11846) );
  OR U12156 ( .A(n11577), .B(n11576), .Z(n11581) );
  OR U12157 ( .A(n11579), .B(n11578), .Z(n11580) );
  AND U12158 ( .A(n11581), .B(n11580), .Z(n11845) );
  XNOR U12159 ( .A(n11846), .B(n11845), .Z(n11848) );
  XNOR U12160 ( .A(n11847), .B(n11848), .Z(n11903) );
  XOR U12161 ( .A(n11904), .B(n11903), .Z(n11906) );
  XNOR U12162 ( .A(n11905), .B(n11906), .Z(n11839) );
  XNOR U12163 ( .A(n11840), .B(n11839), .Z(n11841) );
  XNOR U12164 ( .A(n11842), .B(n11841), .Z(n11910) );
  ANDN U12165 ( .B(o[13]), .A(n15896), .Z(n11909) );
  XOR U12166 ( .A(n11910), .B(n11909), .Z(n11911) );
  NANDN U12167 ( .A(n11583), .B(n11582), .Z(n11587) );
  OR U12168 ( .A(n11585), .B(n11584), .Z(n11586) );
  AND U12169 ( .A(n11587), .B(n11586), .Z(n11915) );
  XNOR U12170 ( .A(n11916), .B(n11915), .Z(n11918) );
  ANDN U12171 ( .B(o[14]), .A(n15935), .Z(n11917) );
  XOR U12172 ( .A(n11918), .B(n11917), .Z(n11834) );
  OR U12173 ( .A(n11589), .B(n11588), .Z(n11593) );
  OR U12174 ( .A(n11591), .B(n11590), .Z(n11592) );
  AND U12175 ( .A(n11593), .B(n11592), .Z(n11833) );
  XNOR U12176 ( .A(n11834), .B(n11833), .Z(n11835) );
  XOR U12177 ( .A(n11836), .B(n11835), .Z(n11828) );
  XOR U12178 ( .A(n11827), .B(n11828), .Z(n11829) );
  XOR U12179 ( .A(n11830), .B(n11829), .Z(n11823) );
  XOR U12180 ( .A(n11824), .B(n11823), .Z(n11816) );
  XNOR U12181 ( .A(n11815), .B(n11816), .Z(n11818) );
  ANDN U12182 ( .B(o[18]), .A(n2993), .Z(n11817) );
  XOR U12183 ( .A(n11818), .B(n11817), .Z(n11923) );
  OR U12184 ( .A(n11595), .B(n11594), .Z(n11599) );
  OR U12185 ( .A(n11597), .B(n11596), .Z(n11598) );
  AND U12186 ( .A(n11599), .B(n11598), .Z(n11922) );
  NANDN U12187 ( .A(n2992), .B(o[19]), .Z(n11921) );
  XOR U12188 ( .A(n11922), .B(n11921), .Z(n11924) );
  XNOR U12189 ( .A(n11923), .B(n11924), .Z(n11809) );
  XNOR U12190 ( .A(n11810), .B(n11809), .Z(n11811) );
  XNOR U12191 ( .A(n11812), .B(n11811), .Z(n11805) );
  OR U12192 ( .A(n11601), .B(n11600), .Z(n11605) );
  NANDN U12193 ( .A(n11603), .B(n11602), .Z(n11604) );
  AND U12194 ( .A(n11605), .B(n11604), .Z(n11804) );
  NANDN U12195 ( .A(n2990), .B(o[21]), .Z(n11803) );
  XOR U12196 ( .A(n11804), .B(n11803), .Z(n11806) );
  XNOR U12197 ( .A(n11805), .B(n11806), .Z(n11927) );
  XNOR U12198 ( .A(n11928), .B(n11927), .Z(n11929) );
  XNOR U12199 ( .A(n11930), .B(n11929), .Z(n11799) );
  NANDN U12200 ( .A(n2988), .B(o[23]), .Z(n11797) );
  OR U12201 ( .A(n11607), .B(n11606), .Z(n11611) );
  OR U12202 ( .A(n11609), .B(n11608), .Z(n11610) );
  NAND U12203 ( .A(n11611), .B(n11610), .Z(n11798) );
  XOR U12204 ( .A(n11797), .B(n11798), .Z(n11800) );
  XNOR U12205 ( .A(n11799), .B(n11800), .Z(n11933) );
  XNOR U12206 ( .A(n11934), .B(n11933), .Z(n11935) );
  XNOR U12207 ( .A(n11936), .B(n11935), .Z(n11793) );
  NANDN U12208 ( .A(n2986), .B(o[25]), .Z(n11791) );
  OR U12209 ( .A(n11613), .B(n11612), .Z(n11617) );
  OR U12210 ( .A(n11615), .B(n11614), .Z(n11616) );
  NAND U12211 ( .A(n11617), .B(n11616), .Z(n11792) );
  XOR U12212 ( .A(n11791), .B(n11792), .Z(n11794) );
  XNOR U12213 ( .A(n11793), .B(n11794), .Z(n11939) );
  XNOR U12214 ( .A(n11940), .B(n11939), .Z(n11941) );
  XNOR U12215 ( .A(n11942), .B(n11941), .Z(n11787) );
  AND U12216 ( .A(o[27]), .B(\stack[1][27] ), .Z(n16433) );
  OR U12217 ( .A(n11619), .B(n11618), .Z(n11623) );
  OR U12218 ( .A(n11621), .B(n11620), .Z(n11622) );
  NAND U12219 ( .A(n11623), .B(n11622), .Z(n11786) );
  XNOR U12220 ( .A(n16433), .B(n11786), .Z(n11788) );
  XNOR U12221 ( .A(n11787), .B(n11788), .Z(n11945) );
  XNOR U12222 ( .A(n11946), .B(n11945), .Z(n11947) );
  XNOR U12223 ( .A(n11948), .B(n11947), .Z(n11782) );
  NANDN U12224 ( .A(n2982), .B(o[29]), .Z(n11780) );
  OR U12225 ( .A(n11625), .B(n11624), .Z(n11629) );
  OR U12226 ( .A(n11627), .B(n11626), .Z(n11628) );
  NAND U12227 ( .A(n11629), .B(n11628), .Z(n11781) );
  XOR U12228 ( .A(n11780), .B(n11781), .Z(n11783) );
  XNOR U12229 ( .A(n11782), .B(n11783), .Z(n11951) );
  XNOR U12230 ( .A(n11952), .B(n11951), .Z(n11953) );
  XNOR U12231 ( .A(n11954), .B(n11953), .Z(n11776) );
  NANDN U12232 ( .A(n2980), .B(o[31]), .Z(n11774) );
  OR U12233 ( .A(n11631), .B(n11630), .Z(n11635) );
  OR U12234 ( .A(n11633), .B(n11632), .Z(n11634) );
  NAND U12235 ( .A(n11635), .B(n11634), .Z(n11775) );
  XOR U12236 ( .A(n11774), .B(n11775), .Z(n11777) );
  XNOR U12237 ( .A(n11776), .B(n11777), .Z(n11957) );
  XNOR U12238 ( .A(n11958), .B(n11957), .Z(n11959) );
  XNOR U12239 ( .A(n11960), .B(n11959), .Z(n11770) );
  NANDN U12240 ( .A(n2978), .B(o[33]), .Z(n11768) );
  OR U12241 ( .A(n11637), .B(n11636), .Z(n11641) );
  OR U12242 ( .A(n11639), .B(n11638), .Z(n11640) );
  NAND U12243 ( .A(n11641), .B(n11640), .Z(n11769) );
  XOR U12244 ( .A(n11768), .B(n11769), .Z(n11771) );
  XNOR U12245 ( .A(n11770), .B(n11771), .Z(n11963) );
  XNOR U12246 ( .A(n11964), .B(n11963), .Z(n11965) );
  XNOR U12247 ( .A(n11966), .B(n11965), .Z(n11764) );
  NANDN U12248 ( .A(n16746), .B(o[35]), .Z(n11762) );
  OR U12249 ( .A(n11643), .B(n11642), .Z(n11647) );
  OR U12250 ( .A(n11645), .B(n11644), .Z(n11646) );
  NAND U12251 ( .A(n11647), .B(n11646), .Z(n11763) );
  XOR U12252 ( .A(n11762), .B(n11763), .Z(n11765) );
  XNOR U12253 ( .A(n11764), .B(n11765), .Z(n11969) );
  XNOR U12254 ( .A(n11970), .B(n11969), .Z(n11971) );
  XNOR U12255 ( .A(n11972), .B(n11971), .Z(n11758) );
  NANDN U12256 ( .A(n16826), .B(o[37]), .Z(n11756) );
  OR U12257 ( .A(n11649), .B(n11648), .Z(n11653) );
  OR U12258 ( .A(n11651), .B(n11650), .Z(n11652) );
  NAND U12259 ( .A(n11653), .B(n11652), .Z(n11757) );
  XOR U12260 ( .A(n11756), .B(n11757), .Z(n11759) );
  XNOR U12261 ( .A(n11758), .B(n11759), .Z(n11975) );
  XNOR U12262 ( .A(n11976), .B(n11975), .Z(n11977) );
  XNOR U12263 ( .A(n11978), .B(n11977), .Z(n11752) );
  NANDN U12264 ( .A(n2976), .B(o[39]), .Z(n11750) );
  OR U12265 ( .A(n11655), .B(n11654), .Z(n11659) );
  OR U12266 ( .A(n11657), .B(n11656), .Z(n11658) );
  NAND U12267 ( .A(n11659), .B(n11658), .Z(n11751) );
  XOR U12268 ( .A(n11750), .B(n11751), .Z(n11753) );
  XNOR U12269 ( .A(n11752), .B(n11753), .Z(n11981) );
  XNOR U12270 ( .A(n11982), .B(n11981), .Z(n11983) );
  XNOR U12271 ( .A(n11984), .B(n11983), .Z(n11746) );
  NANDN U12272 ( .A(n2974), .B(o[41]), .Z(n11744) );
  OR U12273 ( .A(n11661), .B(n11660), .Z(n11665) );
  OR U12274 ( .A(n11663), .B(n11662), .Z(n11664) );
  NAND U12275 ( .A(n11665), .B(n11664), .Z(n11745) );
  XOR U12276 ( .A(n11744), .B(n11745), .Z(n11747) );
  XNOR U12277 ( .A(n11746), .B(n11747), .Z(n11987) );
  XNOR U12278 ( .A(n11988), .B(n11987), .Z(n11989) );
  XNOR U12279 ( .A(n11990), .B(n11989), .Z(n11740) );
  NANDN U12280 ( .A(n2972), .B(o[43]), .Z(n11738) );
  OR U12281 ( .A(n11667), .B(n11666), .Z(n11671) );
  OR U12282 ( .A(n11669), .B(n11668), .Z(n11670) );
  NAND U12283 ( .A(n11671), .B(n11670), .Z(n11739) );
  XOR U12284 ( .A(n11738), .B(n11739), .Z(n11741) );
  XNOR U12285 ( .A(n11740), .B(n11741), .Z(n11993) );
  XNOR U12286 ( .A(n11994), .B(n11993), .Z(n11995) );
  XNOR U12287 ( .A(n11996), .B(n11995), .Z(n11734) );
  NANDN U12288 ( .A(n17145), .B(o[45]), .Z(n11732) );
  OR U12289 ( .A(n11673), .B(n11672), .Z(n11677) );
  OR U12290 ( .A(n11675), .B(n11674), .Z(n11676) );
  NAND U12291 ( .A(n11677), .B(n11676), .Z(n11733) );
  XOR U12292 ( .A(n11732), .B(n11733), .Z(n11735) );
  XNOR U12293 ( .A(n11734), .B(n11735), .Z(n11999) );
  XNOR U12294 ( .A(n12000), .B(n11999), .Z(n12001) );
  XNOR U12295 ( .A(n12002), .B(n12001), .Z(n11728) );
  NANDN U12296 ( .A(n17219), .B(o[47]), .Z(n11726) );
  OR U12297 ( .A(n11679), .B(n11678), .Z(n11683) );
  OR U12298 ( .A(n11681), .B(n11680), .Z(n11682) );
  NAND U12299 ( .A(n11683), .B(n11682), .Z(n11727) );
  XOR U12300 ( .A(n11726), .B(n11727), .Z(n11729) );
  XNOR U12301 ( .A(n11728), .B(n11729), .Z(n12005) );
  XNOR U12302 ( .A(n12006), .B(n12005), .Z(n12007) );
  XNOR U12303 ( .A(n12008), .B(n12007), .Z(n11722) );
  NANDN U12304 ( .A(n17296), .B(o[49]), .Z(n11720) );
  OR U12305 ( .A(n11685), .B(n11684), .Z(n11689) );
  OR U12306 ( .A(n11687), .B(n11686), .Z(n11688) );
  NAND U12307 ( .A(n11689), .B(n11688), .Z(n11721) );
  XOR U12308 ( .A(n11720), .B(n11721), .Z(n11723) );
  XNOR U12309 ( .A(n11722), .B(n11723), .Z(n12011) );
  XNOR U12310 ( .A(n12012), .B(n12011), .Z(n12013) );
  XNOR U12311 ( .A(n12014), .B(n12013), .Z(n11716) );
  NANDN U12312 ( .A(n17375), .B(o[51]), .Z(n11714) );
  OR U12313 ( .A(n11691), .B(n11690), .Z(n11695) );
  OR U12314 ( .A(n11693), .B(n11692), .Z(n11694) );
  NAND U12315 ( .A(n11695), .B(n11694), .Z(n11715) );
  XOR U12316 ( .A(n11714), .B(n11715), .Z(n11717) );
  XNOR U12317 ( .A(n11716), .B(n11717), .Z(n12017) );
  XNOR U12318 ( .A(n12018), .B(n12017), .Z(n12019) );
  AND U12319 ( .A(o[53]), .B(\stack[1][1] ), .Z(n11708) );
  OR U12320 ( .A(n11697), .B(n11696), .Z(n11701) );
  OR U12321 ( .A(n11699), .B(n11698), .Z(n11700) );
  NAND U12322 ( .A(n11701), .B(n11700), .Z(n11709) );
  XNOR U12323 ( .A(n11708), .B(n11709), .Z(n11711) );
  XOR U12324 ( .A(n11710), .B(n11711), .Z(n11702) );
  NANDN U12325 ( .A(n11703), .B(n11702), .Z(n11705) );
  XOR U12326 ( .A(n11703), .B(n11702), .Z(n15394) );
  AND U12327 ( .A(o[54]), .B(\stack[1][0] ), .Z(n15395) );
  OR U12328 ( .A(n15394), .B(n15395), .Z(n11704) );
  AND U12329 ( .A(n11705), .B(n11704), .Z(n11707) );
  OR U12330 ( .A(n11706), .B(n11707), .Z(n12024) );
  XNOR U12331 ( .A(n11707), .B(n11706), .Z(n15356) );
  NANDN U12332 ( .A(n2969), .B(o[54]), .Z(n12344) );
  OR U12333 ( .A(n11709), .B(n11708), .Z(n11713) );
  OR U12334 ( .A(n11711), .B(n11710), .Z(n11712) );
  NAND U12335 ( .A(n11713), .B(n11712), .Z(n12342) );
  NANDN U12336 ( .A(n17375), .B(o[52]), .Z(n12338) );
  NANDN U12337 ( .A(n11715), .B(n11714), .Z(n11719) );
  NANDN U12338 ( .A(n11717), .B(n11716), .Z(n11718) );
  NAND U12339 ( .A(n11719), .B(n11718), .Z(n12336) );
  NANDN U12340 ( .A(n17296), .B(o[50]), .Z(n12332) );
  NANDN U12341 ( .A(n11721), .B(n11720), .Z(n11725) );
  NANDN U12342 ( .A(n11723), .B(n11722), .Z(n11724) );
  NAND U12343 ( .A(n11725), .B(n11724), .Z(n12330) );
  NANDN U12344 ( .A(n17219), .B(o[48]), .Z(n12326) );
  NANDN U12345 ( .A(n11727), .B(n11726), .Z(n11731) );
  NANDN U12346 ( .A(n11729), .B(n11728), .Z(n11730) );
  NAND U12347 ( .A(n11731), .B(n11730), .Z(n12324) );
  NANDN U12348 ( .A(n17145), .B(o[46]), .Z(n12320) );
  NANDN U12349 ( .A(n11733), .B(n11732), .Z(n11737) );
  NANDN U12350 ( .A(n11735), .B(n11734), .Z(n11736) );
  NAND U12351 ( .A(n11737), .B(n11736), .Z(n12318) );
  NANDN U12352 ( .A(n2972), .B(o[44]), .Z(n12314) );
  NANDN U12353 ( .A(n11739), .B(n11738), .Z(n11743) );
  NANDN U12354 ( .A(n11741), .B(n11740), .Z(n11742) );
  NAND U12355 ( .A(n11743), .B(n11742), .Z(n12312) );
  NANDN U12356 ( .A(n2974), .B(o[42]), .Z(n12308) );
  NANDN U12357 ( .A(n11745), .B(n11744), .Z(n11749) );
  NANDN U12358 ( .A(n11747), .B(n11746), .Z(n11748) );
  NAND U12359 ( .A(n11749), .B(n11748), .Z(n12306) );
  NANDN U12360 ( .A(n2976), .B(o[40]), .Z(n12302) );
  NANDN U12361 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U12362 ( .A(n11753), .B(n11752), .Z(n11754) );
  NAND U12363 ( .A(n11755), .B(n11754), .Z(n12300) );
  NANDN U12364 ( .A(n16826), .B(o[38]), .Z(n12296) );
  NANDN U12365 ( .A(n11757), .B(n11756), .Z(n11761) );
  NANDN U12366 ( .A(n11759), .B(n11758), .Z(n11760) );
  NAND U12367 ( .A(n11761), .B(n11760), .Z(n12294) );
  NANDN U12368 ( .A(n16746), .B(o[36]), .Z(n12290) );
  NANDN U12369 ( .A(n11763), .B(n11762), .Z(n11767) );
  NANDN U12370 ( .A(n11765), .B(n11764), .Z(n11766) );
  NAND U12371 ( .A(n11767), .B(n11766), .Z(n12288) );
  NANDN U12372 ( .A(n2978), .B(o[34]), .Z(n12284) );
  NANDN U12373 ( .A(n11769), .B(n11768), .Z(n11773) );
  NANDN U12374 ( .A(n11771), .B(n11770), .Z(n11772) );
  NAND U12375 ( .A(n11773), .B(n11772), .Z(n12282) );
  NANDN U12376 ( .A(n2980), .B(o[32]), .Z(n12278) );
  NANDN U12377 ( .A(n11775), .B(n11774), .Z(n11779) );
  NANDN U12378 ( .A(n11777), .B(n11776), .Z(n11778) );
  NAND U12379 ( .A(n11779), .B(n11778), .Z(n12276) );
  NANDN U12380 ( .A(n2982), .B(o[30]), .Z(n12272) );
  NANDN U12381 ( .A(n11781), .B(n11780), .Z(n11785) );
  NANDN U12382 ( .A(n11783), .B(n11782), .Z(n11784) );
  NAND U12383 ( .A(n11785), .B(n11784), .Z(n12270) );
  NANDN U12384 ( .A(n2984), .B(o[28]), .Z(n12266) );
  OR U12385 ( .A(n11786), .B(n16433), .Z(n11790) );
  NANDN U12386 ( .A(n11788), .B(n11787), .Z(n11789) );
  NAND U12387 ( .A(n11790), .B(n11789), .Z(n12264) );
  NANDN U12388 ( .A(n3020), .B(\stack[1][29] ), .Z(n12260) );
  NANDN U12389 ( .A(n11792), .B(n11791), .Z(n11796) );
  NANDN U12390 ( .A(n11794), .B(n11793), .Z(n11795) );
  NAND U12391 ( .A(n11796), .B(n11795), .Z(n12258) );
  NANDN U12392 ( .A(n3018), .B(\stack[1][31] ), .Z(n12118) );
  NANDN U12393 ( .A(n11798), .B(n11797), .Z(n11802) );
  NANDN U12394 ( .A(n11800), .B(n11799), .Z(n11801) );
  NAND U12395 ( .A(n11802), .B(n11801), .Z(n12116) );
  NANDN U12396 ( .A(n3016), .B(\stack[1][33] ), .Z(n12254) );
  NANDN U12397 ( .A(n11804), .B(n11803), .Z(n11808) );
  NANDN U12398 ( .A(n11806), .B(n11805), .Z(n11807) );
  NAND U12399 ( .A(n11808), .B(n11807), .Z(n12252) );
  AND U12400 ( .A(\stack[1][34] ), .B(o[21]), .Z(n12127) );
  OR U12401 ( .A(n11810), .B(n11809), .Z(n11814) );
  OR U12402 ( .A(n11812), .B(n11811), .Z(n11813) );
  NAND U12403 ( .A(n11814), .B(n11813), .Z(n12128) );
  XNOR U12404 ( .A(n12127), .B(n12128), .Z(n12130) );
  NANDN U12405 ( .A(n3013), .B(\stack[1][36] ), .Z(n12134) );
  OR U12406 ( .A(n11816), .B(n11815), .Z(n11820) );
  NANDN U12407 ( .A(n11818), .B(n11817), .Z(n11819) );
  AND U12408 ( .A(n11820), .B(n11819), .Z(n12133) );
  XNOR U12409 ( .A(n12134), .B(n12133), .Z(n12135) );
  OR U12410 ( .A(n11822), .B(n11821), .Z(n11826) );
  OR U12411 ( .A(n11824), .B(n11823), .Z(n11825) );
  NAND U12412 ( .A(n11826), .B(n11825), .Z(n12140) );
  ANDN U12413 ( .B(\stack[1][38] ), .A(n3011), .Z(n12148) );
  OR U12414 ( .A(n11828), .B(n11827), .Z(n11832) );
  NANDN U12415 ( .A(n11830), .B(n11829), .Z(n11831) );
  AND U12416 ( .A(n11832), .B(n11831), .Z(n12145) );
  OR U12417 ( .A(n11834), .B(n11833), .Z(n11838) );
  OR U12418 ( .A(n11836), .B(n11835), .Z(n11837) );
  AND U12419 ( .A(n11838), .B(n11837), .Z(n12151) );
  NANDN U12420 ( .A(n3010), .B(\stack[1][39] ), .Z(n12152) );
  XOR U12421 ( .A(n12151), .B(n12152), .Z(n12153) );
  OR U12422 ( .A(n11840), .B(n11839), .Z(n11844) );
  OR U12423 ( .A(n11842), .B(n11841), .Z(n11843) );
  AND U12424 ( .A(n11844), .B(n11843), .Z(n12235) );
  NANDN U12425 ( .A(n3006), .B(\stack[1][43] ), .Z(n12164) );
  AND U12426 ( .A(\stack[1][44] ), .B(o[11]), .Z(n12172) );
  OR U12427 ( .A(n11846), .B(n11845), .Z(n11850) );
  NANDN U12428 ( .A(n11848), .B(n11847), .Z(n11849) );
  AND U12429 ( .A(n11850), .B(n11849), .Z(n12169) );
  AND U12430 ( .A(\stack[1][45] ), .B(o[10]), .Z(n12178) );
  AND U12431 ( .A(\stack[1][46] ), .B(o[9]), .Z(n12229) );
  NANDN U12432 ( .A(n11852), .B(n11851), .Z(n11856) );
  NAND U12433 ( .A(n11854), .B(n11853), .Z(n11855) );
  AND U12434 ( .A(n11856), .B(n11855), .Z(n12218) );
  AND U12435 ( .A(\stack[1][50] ), .B(o[5]), .Z(n12212) );
  OR U12436 ( .A(n11858), .B(n11857), .Z(n11862) );
  NANDN U12437 ( .A(n11860), .B(n11859), .Z(n11861) );
  AND U12438 ( .A(n11862), .B(n11861), .Z(n12209) );
  AND U12439 ( .A(\stack[1][51] ), .B(o[4]), .Z(n12190) );
  AND U12440 ( .A(\stack[1][52] ), .B(o[3]), .Z(n12206) );
  NANDN U12441 ( .A(n11863), .B(n12193), .Z(n11864) );
  AND U12442 ( .A(n11865), .B(n11864), .Z(n11869) );
  OR U12443 ( .A(n11867), .B(n11866), .Z(n11868) );
  AND U12444 ( .A(n11869), .B(n11868), .Z(n12203) );
  AND U12445 ( .A(\stack[1][55] ), .B(o[1]), .Z(n12201) );
  ANDN U12446 ( .B(n12201), .A(n11870), .Z(n12521) );
  XNOR U12447 ( .A(n12521), .B(n12193), .Z(n11872) );
  NAND U12448 ( .A(o[0]), .B(\stack[1][55] ), .Z(n12200) );
  NANDN U12449 ( .A(n11871), .B(n12200), .Z(n12195) );
  NAND U12450 ( .A(n11872), .B(n12195), .Z(n12197) );
  ANDN U12451 ( .B(\stack[1][53] ), .A(n2996), .Z(n12196) );
  XNOR U12452 ( .A(n12197), .B(n12196), .Z(n12204) );
  XOR U12453 ( .A(n12203), .B(n12204), .Z(n12205) );
  XOR U12454 ( .A(n12206), .B(n12205), .Z(n12188) );
  OR U12455 ( .A(n11874), .B(n11873), .Z(n11878) );
  NANDN U12456 ( .A(n11876), .B(n11875), .Z(n11877) );
  AND U12457 ( .A(n11878), .B(n11877), .Z(n12187) );
  XOR U12458 ( .A(n12188), .B(n12187), .Z(n12189) );
  XOR U12459 ( .A(n12190), .B(n12189), .Z(n12210) );
  XNOR U12460 ( .A(n12209), .B(n12210), .Z(n12211) );
  OR U12461 ( .A(n11880), .B(n11879), .Z(n11884) );
  OR U12462 ( .A(n11882), .B(n11881), .Z(n11883) );
  NAND U12463 ( .A(n11884), .B(n11883), .Z(n12182) );
  ANDN U12464 ( .B(\stack[1][49] ), .A(n3000), .Z(n12181) );
  XNOR U12465 ( .A(n12182), .B(n12181), .Z(n12184) );
  XNOR U12466 ( .A(n12183), .B(n12184), .Z(n12216) );
  ANDN U12467 ( .B(o[7]), .A(n15623), .Z(n12215) );
  XOR U12468 ( .A(n12216), .B(n12215), .Z(n12217) );
  NANDN U12469 ( .A(n11886), .B(n11885), .Z(n11890) );
  OR U12470 ( .A(n11888), .B(n11887), .Z(n11889) );
  AND U12471 ( .A(n11890), .B(n11889), .Z(n12221) );
  XNOR U12472 ( .A(n12222), .B(n12221), .Z(n12224) );
  AND U12473 ( .A(\stack[1][47] ), .B(o[8]), .Z(n12223) );
  XNOR U12474 ( .A(n12224), .B(n12223), .Z(n12227) );
  OR U12475 ( .A(n11892), .B(n11891), .Z(n11896) );
  NANDN U12476 ( .A(n11894), .B(n11893), .Z(n11895) );
  NAND U12477 ( .A(n11896), .B(n11895), .Z(n12228) );
  XNOR U12478 ( .A(n12227), .B(n12228), .Z(n12230) );
  XNOR U12479 ( .A(n12229), .B(n12230), .Z(n12176) );
  OR U12480 ( .A(n11898), .B(n11897), .Z(n11902) );
  OR U12481 ( .A(n11900), .B(n11899), .Z(n11901) );
  AND U12482 ( .A(n11902), .B(n11901), .Z(n12175) );
  XOR U12483 ( .A(n12176), .B(n12175), .Z(n12177) );
  XOR U12484 ( .A(n12178), .B(n12177), .Z(n12170) );
  XNOR U12485 ( .A(n12169), .B(n12170), .Z(n12171) );
  XOR U12486 ( .A(n12164), .B(n12163), .Z(n12166) );
  NANDN U12487 ( .A(n11904), .B(n11903), .Z(n11908) );
  NANDN U12488 ( .A(n11906), .B(n11905), .Z(n11907) );
  NAND U12489 ( .A(n11908), .B(n11907), .Z(n12165) );
  XNOR U12490 ( .A(n12166), .B(n12165), .Z(n12234) );
  ANDN U12491 ( .B(o[13]), .A(n15857), .Z(n12233) );
  XOR U12492 ( .A(n12234), .B(n12233), .Z(n12236) );
  XNOR U12493 ( .A(n12235), .B(n12236), .Z(n12240) );
  NANDN U12494 ( .A(n11910), .B(n11909), .Z(n11914) );
  OR U12495 ( .A(n11912), .B(n11911), .Z(n11913) );
  AND U12496 ( .A(n11914), .B(n11913), .Z(n12239) );
  XNOR U12497 ( .A(n12240), .B(n12239), .Z(n12242) );
  ANDN U12498 ( .B(o[14]), .A(n15896), .Z(n12241) );
  XOR U12499 ( .A(n12242), .B(n12241), .Z(n12158) );
  OR U12500 ( .A(n11916), .B(n11915), .Z(n11920) );
  NANDN U12501 ( .A(n11918), .B(n11917), .Z(n11919) );
  AND U12502 ( .A(n11920), .B(n11919), .Z(n12157) );
  XNOR U12503 ( .A(n12158), .B(n12157), .Z(n12160) );
  ANDN U12504 ( .B(o[15]), .A(n15935), .Z(n12159) );
  XOR U12505 ( .A(n12160), .B(n12159), .Z(n12154) );
  XNOR U12506 ( .A(n12153), .B(n12154), .Z(n12146) );
  XNOR U12507 ( .A(n12145), .B(n12146), .Z(n12147) );
  XOR U12508 ( .A(n12140), .B(n12139), .Z(n12142) );
  NANDN U12509 ( .A(n3012), .B(\stack[1][37] ), .Z(n12141) );
  XNOR U12510 ( .A(n12142), .B(n12141), .Z(n12136) );
  NANDN U12511 ( .A(n11922), .B(n11921), .Z(n11926) );
  NANDN U12512 ( .A(n11924), .B(n11923), .Z(n11925) );
  AND U12513 ( .A(n11926), .B(n11925), .Z(n12246) );
  XNOR U12514 ( .A(n12245), .B(n12246), .Z(n12248) );
  AND U12515 ( .A(\stack[1][35] ), .B(o[20]), .Z(n12247) );
  XNOR U12516 ( .A(n12248), .B(n12247), .Z(n12129) );
  XOR U12517 ( .A(n12130), .B(n12129), .Z(n12251) );
  XNOR U12518 ( .A(n12252), .B(n12251), .Z(n12253) );
  XNOR U12519 ( .A(n12254), .B(n12253), .Z(n12123) );
  NANDN U12520 ( .A(n2989), .B(o[23]), .Z(n12121) );
  OR U12521 ( .A(n11928), .B(n11927), .Z(n11932) );
  OR U12522 ( .A(n11930), .B(n11929), .Z(n11931) );
  NAND U12523 ( .A(n11932), .B(n11931), .Z(n12122) );
  XOR U12524 ( .A(n12121), .B(n12122), .Z(n12124) );
  XNOR U12525 ( .A(n12123), .B(n12124), .Z(n12115) );
  XNOR U12526 ( .A(n12116), .B(n12115), .Z(n12117) );
  XNOR U12527 ( .A(n12118), .B(n12117), .Z(n12111) );
  NANDN U12528 ( .A(n2987), .B(o[25]), .Z(n12109) );
  OR U12529 ( .A(n11934), .B(n11933), .Z(n11938) );
  OR U12530 ( .A(n11936), .B(n11935), .Z(n11937) );
  NAND U12531 ( .A(n11938), .B(n11937), .Z(n12110) );
  XOR U12532 ( .A(n12109), .B(n12110), .Z(n12112) );
  XNOR U12533 ( .A(n12111), .B(n12112), .Z(n12257) );
  XNOR U12534 ( .A(n12258), .B(n12257), .Z(n12259) );
  XNOR U12535 ( .A(n12260), .B(n12259), .Z(n12105) );
  NANDN U12536 ( .A(n2985), .B(o[27]), .Z(n12103) );
  OR U12537 ( .A(n11940), .B(n11939), .Z(n11944) );
  OR U12538 ( .A(n11942), .B(n11941), .Z(n11943) );
  NAND U12539 ( .A(n11944), .B(n11943), .Z(n12104) );
  XOR U12540 ( .A(n12103), .B(n12104), .Z(n12106) );
  XNOR U12541 ( .A(n12105), .B(n12106), .Z(n12263) );
  XNOR U12542 ( .A(n12264), .B(n12263), .Z(n12265) );
  XNOR U12543 ( .A(n12266), .B(n12265), .Z(n12099) );
  NANDN U12544 ( .A(n2983), .B(o[29]), .Z(n12097) );
  OR U12545 ( .A(n11946), .B(n11945), .Z(n11950) );
  OR U12546 ( .A(n11948), .B(n11947), .Z(n11949) );
  NAND U12547 ( .A(n11950), .B(n11949), .Z(n12098) );
  XOR U12548 ( .A(n12097), .B(n12098), .Z(n12100) );
  XNOR U12549 ( .A(n12099), .B(n12100), .Z(n12269) );
  XNOR U12550 ( .A(n12270), .B(n12269), .Z(n12271) );
  XNOR U12551 ( .A(n12272), .B(n12271), .Z(n12093) );
  NANDN U12552 ( .A(n2981), .B(o[31]), .Z(n12091) );
  OR U12553 ( .A(n11952), .B(n11951), .Z(n11956) );
  OR U12554 ( .A(n11954), .B(n11953), .Z(n11955) );
  NAND U12555 ( .A(n11956), .B(n11955), .Z(n12092) );
  XOR U12556 ( .A(n12091), .B(n12092), .Z(n12094) );
  XNOR U12557 ( .A(n12093), .B(n12094), .Z(n12275) );
  XNOR U12558 ( .A(n12276), .B(n12275), .Z(n12277) );
  XNOR U12559 ( .A(n12278), .B(n12277), .Z(n12087) );
  NANDN U12560 ( .A(n2979), .B(o[33]), .Z(n12085) );
  OR U12561 ( .A(n11958), .B(n11957), .Z(n11962) );
  OR U12562 ( .A(n11960), .B(n11959), .Z(n11961) );
  NAND U12563 ( .A(n11962), .B(n11961), .Z(n12086) );
  XOR U12564 ( .A(n12085), .B(n12086), .Z(n12088) );
  XNOR U12565 ( .A(n12087), .B(n12088), .Z(n12281) );
  XNOR U12566 ( .A(n12282), .B(n12281), .Z(n12283) );
  XNOR U12567 ( .A(n12284), .B(n12283), .Z(n12081) );
  NANDN U12568 ( .A(n16712), .B(o[35]), .Z(n12079) );
  OR U12569 ( .A(n11964), .B(n11963), .Z(n11968) );
  OR U12570 ( .A(n11966), .B(n11965), .Z(n11967) );
  NAND U12571 ( .A(n11968), .B(n11967), .Z(n12080) );
  XOR U12572 ( .A(n12079), .B(n12080), .Z(n12082) );
  XNOR U12573 ( .A(n12081), .B(n12082), .Z(n12287) );
  XNOR U12574 ( .A(n12288), .B(n12287), .Z(n12289) );
  XNOR U12575 ( .A(n12290), .B(n12289), .Z(n12075) );
  NANDN U12576 ( .A(n16786), .B(o[37]), .Z(n12073) );
  OR U12577 ( .A(n11970), .B(n11969), .Z(n11974) );
  OR U12578 ( .A(n11972), .B(n11971), .Z(n11973) );
  NAND U12579 ( .A(n11974), .B(n11973), .Z(n12074) );
  XOR U12580 ( .A(n12073), .B(n12074), .Z(n12076) );
  XNOR U12581 ( .A(n12075), .B(n12076), .Z(n12293) );
  XNOR U12582 ( .A(n12294), .B(n12293), .Z(n12295) );
  XNOR U12583 ( .A(n12296), .B(n12295), .Z(n12069) );
  NANDN U12584 ( .A(n2977), .B(o[39]), .Z(n12067) );
  OR U12585 ( .A(n11976), .B(n11975), .Z(n11980) );
  OR U12586 ( .A(n11978), .B(n11977), .Z(n11979) );
  NAND U12587 ( .A(n11980), .B(n11979), .Z(n12068) );
  XOR U12588 ( .A(n12067), .B(n12068), .Z(n12070) );
  XNOR U12589 ( .A(n12069), .B(n12070), .Z(n12299) );
  XNOR U12590 ( .A(n12300), .B(n12299), .Z(n12301) );
  XNOR U12591 ( .A(n12302), .B(n12301), .Z(n12063) );
  NANDN U12592 ( .A(n2975), .B(o[41]), .Z(n12061) );
  OR U12593 ( .A(n11982), .B(n11981), .Z(n11986) );
  OR U12594 ( .A(n11984), .B(n11983), .Z(n11985) );
  NAND U12595 ( .A(n11986), .B(n11985), .Z(n12062) );
  XOR U12596 ( .A(n12061), .B(n12062), .Z(n12064) );
  XNOR U12597 ( .A(n12063), .B(n12064), .Z(n12305) );
  XNOR U12598 ( .A(n12306), .B(n12305), .Z(n12307) );
  XNOR U12599 ( .A(n12308), .B(n12307), .Z(n12057) );
  NANDN U12600 ( .A(n2973), .B(o[43]), .Z(n12055) );
  OR U12601 ( .A(n11988), .B(n11987), .Z(n11992) );
  OR U12602 ( .A(n11990), .B(n11989), .Z(n11991) );
  NAND U12603 ( .A(n11992), .B(n11991), .Z(n12056) );
  XOR U12604 ( .A(n12055), .B(n12056), .Z(n12058) );
  XNOR U12605 ( .A(n12057), .B(n12058), .Z(n12311) );
  XNOR U12606 ( .A(n12312), .B(n12311), .Z(n12313) );
  XNOR U12607 ( .A(n12314), .B(n12313), .Z(n12051) );
  NANDN U12608 ( .A(n17101), .B(o[45]), .Z(n12049) );
  OR U12609 ( .A(n11994), .B(n11993), .Z(n11998) );
  OR U12610 ( .A(n11996), .B(n11995), .Z(n11997) );
  NAND U12611 ( .A(n11998), .B(n11997), .Z(n12050) );
  XOR U12612 ( .A(n12049), .B(n12050), .Z(n12052) );
  XNOR U12613 ( .A(n12051), .B(n12052), .Z(n12317) );
  XNOR U12614 ( .A(n12318), .B(n12317), .Z(n12319) );
  XNOR U12615 ( .A(n12320), .B(n12319), .Z(n12045) );
  NANDN U12616 ( .A(n17179), .B(o[47]), .Z(n12043) );
  OR U12617 ( .A(n12000), .B(n11999), .Z(n12004) );
  OR U12618 ( .A(n12002), .B(n12001), .Z(n12003) );
  NAND U12619 ( .A(n12004), .B(n12003), .Z(n12044) );
  XOR U12620 ( .A(n12043), .B(n12044), .Z(n12046) );
  XNOR U12621 ( .A(n12045), .B(n12046), .Z(n12323) );
  XNOR U12622 ( .A(n12324), .B(n12323), .Z(n12325) );
  XNOR U12623 ( .A(n12326), .B(n12325), .Z(n12039) );
  NANDN U12624 ( .A(n17256), .B(o[49]), .Z(n12037) );
  OR U12625 ( .A(n12006), .B(n12005), .Z(n12010) );
  OR U12626 ( .A(n12008), .B(n12007), .Z(n12009) );
  NAND U12627 ( .A(n12010), .B(n12009), .Z(n12038) );
  XOR U12628 ( .A(n12037), .B(n12038), .Z(n12040) );
  XNOR U12629 ( .A(n12039), .B(n12040), .Z(n12329) );
  XNOR U12630 ( .A(n12330), .B(n12329), .Z(n12331) );
  XNOR U12631 ( .A(n12332), .B(n12331), .Z(n12033) );
  AND U12632 ( .A(o[51]), .B(\stack[1][4] ), .Z(n12031) );
  OR U12633 ( .A(n12012), .B(n12011), .Z(n12016) );
  OR U12634 ( .A(n12014), .B(n12013), .Z(n12015) );
  NAND U12635 ( .A(n12016), .B(n12015), .Z(n12032) );
  XNOR U12636 ( .A(n12031), .B(n12032), .Z(n12034) );
  XNOR U12637 ( .A(n12033), .B(n12034), .Z(n12335) );
  XNOR U12638 ( .A(n12336), .B(n12335), .Z(n12337) );
  XOR U12639 ( .A(n12338), .B(n12337), .Z(n12028) );
  AND U12640 ( .A(o[53]), .B(\stack[1][2] ), .Z(n12025) );
  OR U12641 ( .A(n12018), .B(n12017), .Z(n12022) );
  OR U12642 ( .A(n12020), .B(n12019), .Z(n12021) );
  NAND U12643 ( .A(n12022), .B(n12021), .Z(n12026) );
  XOR U12644 ( .A(n12025), .B(n12026), .Z(n12027) );
  XNOR U12645 ( .A(n12028), .B(n12027), .Z(n12341) );
  XNOR U12646 ( .A(n12342), .B(n12341), .Z(n12343) );
  XOR U12647 ( .A(n12344), .B(n12343), .Z(n15357) );
  OR U12648 ( .A(n15356), .B(n15357), .Z(n12023) );
  AND U12649 ( .A(n12024), .B(n12023), .Z(n12348) );
  NANDN U12650 ( .A(n2970), .B(o[54]), .Z(n12678) );
  OR U12651 ( .A(n12026), .B(n12025), .Z(n12030) );
  NANDN U12652 ( .A(n12028), .B(n12027), .Z(n12029) );
  NAND U12653 ( .A(n12030), .B(n12029), .Z(n12676) );
  NANDN U12654 ( .A(n2971), .B(o[52]), .Z(n12672) );
  OR U12655 ( .A(n12032), .B(n12031), .Z(n12036) );
  NANDN U12656 ( .A(n12034), .B(n12033), .Z(n12035) );
  NAND U12657 ( .A(n12036), .B(n12035), .Z(n12670) );
  NANDN U12658 ( .A(n17256), .B(o[50]), .Z(n12666) );
  NANDN U12659 ( .A(n12038), .B(n12037), .Z(n12042) );
  NANDN U12660 ( .A(n12040), .B(n12039), .Z(n12041) );
  NAND U12661 ( .A(n12042), .B(n12041), .Z(n12664) );
  NANDN U12662 ( .A(n17179), .B(o[48]), .Z(n12660) );
  NANDN U12663 ( .A(n12044), .B(n12043), .Z(n12048) );
  NANDN U12664 ( .A(n12046), .B(n12045), .Z(n12047) );
  NAND U12665 ( .A(n12048), .B(n12047), .Z(n12658) );
  NANDN U12666 ( .A(n17101), .B(o[46]), .Z(n12654) );
  NANDN U12667 ( .A(n12050), .B(n12049), .Z(n12054) );
  NANDN U12668 ( .A(n12052), .B(n12051), .Z(n12053) );
  NAND U12669 ( .A(n12054), .B(n12053), .Z(n12652) );
  NANDN U12670 ( .A(n2973), .B(o[44]), .Z(n12648) );
  NANDN U12671 ( .A(n12056), .B(n12055), .Z(n12060) );
  NANDN U12672 ( .A(n12058), .B(n12057), .Z(n12059) );
  NAND U12673 ( .A(n12060), .B(n12059), .Z(n12646) );
  NANDN U12674 ( .A(n2975), .B(o[42]), .Z(n12642) );
  NANDN U12675 ( .A(n12062), .B(n12061), .Z(n12066) );
  NANDN U12676 ( .A(n12064), .B(n12063), .Z(n12065) );
  NAND U12677 ( .A(n12066), .B(n12065), .Z(n12640) );
  NANDN U12678 ( .A(n2977), .B(o[40]), .Z(n12636) );
  NANDN U12679 ( .A(n12068), .B(n12067), .Z(n12072) );
  NANDN U12680 ( .A(n12070), .B(n12069), .Z(n12071) );
  NAND U12681 ( .A(n12072), .B(n12071), .Z(n12634) );
  NANDN U12682 ( .A(n16786), .B(o[38]), .Z(n12630) );
  NANDN U12683 ( .A(n12074), .B(n12073), .Z(n12078) );
  NANDN U12684 ( .A(n12076), .B(n12075), .Z(n12077) );
  NAND U12685 ( .A(n12078), .B(n12077), .Z(n12628) );
  NANDN U12686 ( .A(n16712), .B(o[36]), .Z(n12624) );
  NANDN U12687 ( .A(n12080), .B(n12079), .Z(n12084) );
  NANDN U12688 ( .A(n12082), .B(n12081), .Z(n12083) );
  NAND U12689 ( .A(n12084), .B(n12083), .Z(n12622) );
  NANDN U12690 ( .A(n2979), .B(o[34]), .Z(n12618) );
  NANDN U12691 ( .A(n12086), .B(n12085), .Z(n12090) );
  NANDN U12692 ( .A(n12088), .B(n12087), .Z(n12089) );
  NAND U12693 ( .A(n12090), .B(n12089), .Z(n12616) );
  NANDN U12694 ( .A(n2981), .B(o[32]), .Z(n12612) );
  NANDN U12695 ( .A(n12092), .B(n12091), .Z(n12096) );
  NANDN U12696 ( .A(n12094), .B(n12093), .Z(n12095) );
  NAND U12697 ( .A(n12096), .B(n12095), .Z(n12610) );
  NANDN U12698 ( .A(n2983), .B(o[30]), .Z(n12606) );
  NANDN U12699 ( .A(n12098), .B(n12097), .Z(n12102) );
  NANDN U12700 ( .A(n12100), .B(n12099), .Z(n12101) );
  NAND U12701 ( .A(n12102), .B(n12101), .Z(n12604) );
  NOR U12702 ( .A(n3021), .B(n2985), .Z(n12599) );
  NANDN U12703 ( .A(n12104), .B(n12103), .Z(n12108) );
  NANDN U12704 ( .A(n12106), .B(n12105), .Z(n12107) );
  NAND U12705 ( .A(n12108), .B(n12107), .Z(n12598) );
  AND U12706 ( .A(\stack[1][30] ), .B(o[26]), .Z(n12446) );
  NANDN U12707 ( .A(n12110), .B(n12109), .Z(n12114) );
  NANDN U12708 ( .A(n12112), .B(n12111), .Z(n12113) );
  AND U12709 ( .A(n12114), .B(n12113), .Z(n12443) );
  AND U12710 ( .A(\stack[1][31] ), .B(o[25]), .Z(n12591) );
  OR U12711 ( .A(n12116), .B(n12115), .Z(n12120) );
  OR U12712 ( .A(n12118), .B(n12117), .Z(n12119) );
  NAND U12713 ( .A(n12120), .B(n12119), .Z(n12592) );
  XNOR U12714 ( .A(n12591), .B(n12592), .Z(n12594) );
  NANDN U12715 ( .A(n12122), .B(n12121), .Z(n12126) );
  NANDN U12716 ( .A(n12124), .B(n12123), .Z(n12125) );
  AND U12717 ( .A(n12126), .B(n12125), .Z(n12449) );
  OR U12718 ( .A(n12128), .B(n12127), .Z(n12132) );
  OR U12719 ( .A(n12130), .B(n12129), .Z(n12131) );
  NAND U12720 ( .A(n12132), .B(n12131), .Z(n12586) );
  AND U12721 ( .A(\stack[1][36] ), .B(o[20]), .Z(n12581) );
  OR U12722 ( .A(n12134), .B(n12133), .Z(n12138) );
  OR U12723 ( .A(n12136), .B(n12135), .Z(n12137) );
  NAND U12724 ( .A(n12138), .B(n12137), .Z(n12580) );
  AND U12725 ( .A(\stack[1][37] ), .B(o[19]), .Z(n12467) );
  NANDN U12726 ( .A(n12140), .B(n12139), .Z(n12144) );
  OR U12727 ( .A(n12142), .B(n12141), .Z(n12143) );
  NAND U12728 ( .A(n12144), .B(n12143), .Z(n12468) );
  XNOR U12729 ( .A(n12467), .B(n12468), .Z(n12470) );
  ANDN U12730 ( .B(\stack[1][38] ), .A(n3012), .Z(n12475) );
  OR U12731 ( .A(n12146), .B(n12145), .Z(n12150) );
  OR U12732 ( .A(n12148), .B(n12147), .Z(n12149) );
  AND U12733 ( .A(n12150), .B(n12149), .Z(n12473) );
  OR U12734 ( .A(n12152), .B(n12151), .Z(n12156) );
  NANDN U12735 ( .A(n12154), .B(n12153), .Z(n12155) );
  AND U12736 ( .A(n12156), .B(n12155), .Z(n12576) );
  OR U12737 ( .A(n12158), .B(n12157), .Z(n12162) );
  NANDN U12738 ( .A(n12160), .B(n12159), .Z(n12161) );
  AND U12739 ( .A(n12162), .B(n12161), .Z(n12479) );
  NANDN U12740 ( .A(n3010), .B(\stack[1][40] ), .Z(n12480) );
  XOR U12741 ( .A(n12479), .B(n12480), .Z(n12482) );
  NANDN U12742 ( .A(n3009), .B(\stack[1][41] ), .Z(n12488) );
  NANDN U12743 ( .A(n12164), .B(n12163), .Z(n12168) );
  OR U12744 ( .A(n12166), .B(n12165), .Z(n12167) );
  AND U12745 ( .A(n12168), .B(n12167), .Z(n12564) );
  OR U12746 ( .A(n12170), .B(n12169), .Z(n12174) );
  OR U12747 ( .A(n12172), .B(n12171), .Z(n12173) );
  NAND U12748 ( .A(n12174), .B(n12173), .Z(n12494) );
  NANDN U12749 ( .A(n3006), .B(\stack[1][44] ), .Z(n12492) );
  NANDN U12750 ( .A(n15740), .B(o[11]), .Z(n12499) );
  OR U12751 ( .A(n12176), .B(n12175), .Z(n12180) );
  NANDN U12752 ( .A(n12178), .B(n12177), .Z(n12179) );
  AND U12753 ( .A(n12180), .B(n12179), .Z(n12498) );
  NANDN U12754 ( .A(n15701), .B(o[10]), .Z(n12505) );
  AND U12755 ( .A(\stack[1][47] ), .B(o[9]), .Z(n12557) );
  NANDN U12756 ( .A(n12182), .B(n12181), .Z(n12186) );
  NAND U12757 ( .A(n12184), .B(n12183), .Z(n12185) );
  AND U12758 ( .A(n12186), .B(n12185), .Z(n12546) );
  AND U12759 ( .A(\stack[1][51] ), .B(o[5]), .Z(n12540) );
  OR U12760 ( .A(n12188), .B(n12187), .Z(n12192) );
  NANDN U12761 ( .A(n12190), .B(n12189), .Z(n12191) );
  AND U12762 ( .A(n12192), .B(n12191), .Z(n12537) );
  AND U12763 ( .A(\stack[1][52] ), .B(o[4]), .Z(n12518) );
  ANDN U12764 ( .B(\stack[1][53] ), .A(n2997), .Z(n12534) );
  NANDN U12765 ( .A(n12193), .B(n12521), .Z(n12194) );
  AND U12766 ( .A(n12195), .B(n12194), .Z(n12199) );
  OR U12767 ( .A(n12197), .B(n12196), .Z(n12198) );
  AND U12768 ( .A(n12199), .B(n12198), .Z(n12531) );
  AND U12769 ( .A(\stack[1][56] ), .B(o[1]), .Z(n12529) );
  ANDN U12770 ( .B(n12529), .A(n12200), .Z(n12857) );
  XNOR U12771 ( .A(n12857), .B(n12521), .Z(n12202) );
  NAND U12772 ( .A(\stack[1][56] ), .B(o[0]), .Z(n12528) );
  NANDN U12773 ( .A(n12201), .B(n12528), .Z(n12523) );
  NAND U12774 ( .A(n12202), .B(n12523), .Z(n12525) );
  ANDN U12775 ( .B(\stack[1][54] ), .A(n2996), .Z(n12524) );
  XNOR U12776 ( .A(n12525), .B(n12524), .Z(n12532) );
  XOR U12777 ( .A(n12531), .B(n12532), .Z(n12533) );
  XOR U12778 ( .A(n12534), .B(n12533), .Z(n12516) );
  OR U12779 ( .A(n12204), .B(n12203), .Z(n12208) );
  NANDN U12780 ( .A(n12206), .B(n12205), .Z(n12207) );
  AND U12781 ( .A(n12208), .B(n12207), .Z(n12515) );
  XOR U12782 ( .A(n12516), .B(n12515), .Z(n12517) );
  XOR U12783 ( .A(n12518), .B(n12517), .Z(n12538) );
  XNOR U12784 ( .A(n12537), .B(n12538), .Z(n12539) );
  OR U12785 ( .A(n12210), .B(n12209), .Z(n12214) );
  OR U12786 ( .A(n12212), .B(n12211), .Z(n12213) );
  NAND U12787 ( .A(n12214), .B(n12213), .Z(n12510) );
  IV U12788 ( .A(\stack[1][50] ), .Z(n15546) );
  ANDN U12789 ( .B(o[6]), .A(n15546), .Z(n12509) );
  XNOR U12790 ( .A(n12510), .B(n12509), .Z(n12512) );
  XNOR U12791 ( .A(n12511), .B(n12512), .Z(n12544) );
  ANDN U12792 ( .B(\stack[1][49] ), .A(n3001), .Z(n12543) );
  XOR U12793 ( .A(n12544), .B(n12543), .Z(n12545) );
  NANDN U12794 ( .A(n12216), .B(n12215), .Z(n12220) );
  OR U12795 ( .A(n12218), .B(n12217), .Z(n12219) );
  AND U12796 ( .A(n12220), .B(n12219), .Z(n12549) );
  XNOR U12797 ( .A(n12550), .B(n12549), .Z(n12552) );
  AND U12798 ( .A(\stack[1][48] ), .B(o[8]), .Z(n12551) );
  XNOR U12799 ( .A(n12552), .B(n12551), .Z(n12555) );
  OR U12800 ( .A(n12222), .B(n12221), .Z(n12226) );
  NANDN U12801 ( .A(n12224), .B(n12223), .Z(n12225) );
  NAND U12802 ( .A(n12226), .B(n12225), .Z(n12556) );
  XNOR U12803 ( .A(n12555), .B(n12556), .Z(n12558) );
  XNOR U12804 ( .A(n12557), .B(n12558), .Z(n12504) );
  OR U12805 ( .A(n12228), .B(n12227), .Z(n12232) );
  OR U12806 ( .A(n12230), .B(n12229), .Z(n12231) );
  AND U12807 ( .A(n12232), .B(n12231), .Z(n12503) );
  XNOR U12808 ( .A(n12504), .B(n12503), .Z(n12506) );
  XNOR U12809 ( .A(n12505), .B(n12506), .Z(n12497) );
  XOR U12810 ( .A(n12498), .B(n12497), .Z(n12500) );
  XNOR U12811 ( .A(n12499), .B(n12500), .Z(n12491) );
  XNOR U12812 ( .A(n12492), .B(n12491), .Z(n12493) );
  XNOR U12813 ( .A(n12494), .B(n12493), .Z(n12562) );
  ANDN U12814 ( .B(o[13]), .A(n15818), .Z(n12561) );
  XOR U12815 ( .A(n12562), .B(n12561), .Z(n12563) );
  NANDN U12816 ( .A(n12234), .B(n12233), .Z(n12238) );
  OR U12817 ( .A(n12236), .B(n12235), .Z(n12237) );
  AND U12818 ( .A(n12238), .B(n12237), .Z(n12567) );
  XNOR U12819 ( .A(n12568), .B(n12567), .Z(n12570) );
  ANDN U12820 ( .B(o[14]), .A(n15857), .Z(n12569) );
  XOR U12821 ( .A(n12570), .B(n12569), .Z(n12486) );
  OR U12822 ( .A(n12240), .B(n12239), .Z(n12244) );
  NANDN U12823 ( .A(n12242), .B(n12241), .Z(n12243) );
  AND U12824 ( .A(n12244), .B(n12243), .Z(n12485) );
  XNOR U12825 ( .A(n12486), .B(n12485), .Z(n12487) );
  XOR U12826 ( .A(n12488), .B(n12487), .Z(n12481) );
  XNOR U12827 ( .A(n12482), .B(n12481), .Z(n12574) );
  NANDN U12828 ( .A(n3011), .B(\stack[1][39] ), .Z(n12573) );
  XOR U12829 ( .A(n12574), .B(n12573), .Z(n12575) );
  XNOR U12830 ( .A(n12576), .B(n12575), .Z(n12474) );
  XNOR U12831 ( .A(n12473), .B(n12474), .Z(n12476) );
  XNOR U12832 ( .A(n12475), .B(n12476), .Z(n12469) );
  XNOR U12833 ( .A(n12470), .B(n12469), .Z(n12579) );
  XNOR U12834 ( .A(n12580), .B(n12579), .Z(n12582) );
  XNOR U12835 ( .A(n12581), .B(n12582), .Z(n12464) );
  OR U12836 ( .A(n12246), .B(n12245), .Z(n12250) );
  OR U12837 ( .A(n12248), .B(n12247), .Z(n12249) );
  AND U12838 ( .A(n12250), .B(n12249), .Z(n12462) );
  NANDN U12839 ( .A(n2992), .B(o[21]), .Z(n12461) );
  XOR U12840 ( .A(n12462), .B(n12461), .Z(n12463) );
  XNOR U12841 ( .A(n12464), .B(n12463), .Z(n12585) );
  XOR U12842 ( .A(n12586), .B(n12585), .Z(n12588) );
  AND U12843 ( .A(\stack[1][34] ), .B(o[22]), .Z(n12587) );
  XNOR U12844 ( .A(n12588), .B(n12587), .Z(n12457) );
  AND U12845 ( .A(\stack[1][33] ), .B(o[23]), .Z(n12455) );
  OR U12846 ( .A(n12252), .B(n12251), .Z(n12256) );
  OR U12847 ( .A(n12254), .B(n12253), .Z(n12255) );
  NAND U12848 ( .A(n12256), .B(n12255), .Z(n12456) );
  XNOR U12849 ( .A(n12455), .B(n12456), .Z(n12458) );
  XNOR U12850 ( .A(n12457), .B(n12458), .Z(n12450) );
  XNOR U12851 ( .A(n12449), .B(n12450), .Z(n12451) );
  AND U12852 ( .A(\stack[1][32] ), .B(o[24]), .Z(n12452) );
  XNOR U12853 ( .A(n12594), .B(n12593), .Z(n12444) );
  XOR U12854 ( .A(n12443), .B(n12444), .Z(n12445) );
  XOR U12855 ( .A(n12446), .B(n12445), .Z(n12440) );
  AND U12856 ( .A(o[27]), .B(\stack[1][29] ), .Z(n12437) );
  OR U12857 ( .A(n12258), .B(n12257), .Z(n12262) );
  OR U12858 ( .A(n12260), .B(n12259), .Z(n12261) );
  NAND U12859 ( .A(n12262), .B(n12261), .Z(n12438) );
  XNOR U12860 ( .A(n12437), .B(n12438), .Z(n12439) );
  XOR U12861 ( .A(n12440), .B(n12439), .Z(n12597) );
  XNOR U12862 ( .A(n12598), .B(n12597), .Z(n12600) );
  XOR U12863 ( .A(n12599), .B(n12600), .Z(n12433) );
  NANDN U12864 ( .A(n2984), .B(o[29]), .Z(n12431) );
  OR U12865 ( .A(n12264), .B(n12263), .Z(n12268) );
  OR U12866 ( .A(n12266), .B(n12265), .Z(n12267) );
  NAND U12867 ( .A(n12268), .B(n12267), .Z(n12432) );
  XOR U12868 ( .A(n12431), .B(n12432), .Z(n12434) );
  XNOR U12869 ( .A(n12433), .B(n12434), .Z(n12603) );
  XNOR U12870 ( .A(n12604), .B(n12603), .Z(n12605) );
  XNOR U12871 ( .A(n12606), .B(n12605), .Z(n12427) );
  NANDN U12872 ( .A(n2982), .B(o[31]), .Z(n12425) );
  OR U12873 ( .A(n12270), .B(n12269), .Z(n12274) );
  OR U12874 ( .A(n12272), .B(n12271), .Z(n12273) );
  NAND U12875 ( .A(n12274), .B(n12273), .Z(n12426) );
  XOR U12876 ( .A(n12425), .B(n12426), .Z(n12428) );
  XNOR U12877 ( .A(n12427), .B(n12428), .Z(n12609) );
  XNOR U12878 ( .A(n12610), .B(n12609), .Z(n12611) );
  XNOR U12879 ( .A(n12612), .B(n12611), .Z(n12421) );
  NANDN U12880 ( .A(n2980), .B(o[33]), .Z(n12419) );
  OR U12881 ( .A(n12276), .B(n12275), .Z(n12280) );
  OR U12882 ( .A(n12278), .B(n12277), .Z(n12279) );
  NAND U12883 ( .A(n12280), .B(n12279), .Z(n12420) );
  XOR U12884 ( .A(n12419), .B(n12420), .Z(n12422) );
  XNOR U12885 ( .A(n12421), .B(n12422), .Z(n12615) );
  XNOR U12886 ( .A(n12616), .B(n12615), .Z(n12617) );
  XNOR U12887 ( .A(n12618), .B(n12617), .Z(n12415) );
  NANDN U12888 ( .A(n2978), .B(o[35]), .Z(n12413) );
  OR U12889 ( .A(n12282), .B(n12281), .Z(n12286) );
  OR U12890 ( .A(n12284), .B(n12283), .Z(n12285) );
  NAND U12891 ( .A(n12286), .B(n12285), .Z(n12414) );
  XOR U12892 ( .A(n12413), .B(n12414), .Z(n12416) );
  XNOR U12893 ( .A(n12415), .B(n12416), .Z(n12621) );
  XNOR U12894 ( .A(n12622), .B(n12621), .Z(n12623) );
  XNOR U12895 ( .A(n12624), .B(n12623), .Z(n12409) );
  NANDN U12896 ( .A(n16746), .B(o[37]), .Z(n12407) );
  OR U12897 ( .A(n12288), .B(n12287), .Z(n12292) );
  OR U12898 ( .A(n12290), .B(n12289), .Z(n12291) );
  NAND U12899 ( .A(n12292), .B(n12291), .Z(n12408) );
  XOR U12900 ( .A(n12407), .B(n12408), .Z(n12410) );
  XNOR U12901 ( .A(n12409), .B(n12410), .Z(n12627) );
  XNOR U12902 ( .A(n12628), .B(n12627), .Z(n12629) );
  XNOR U12903 ( .A(n12630), .B(n12629), .Z(n12403) );
  NANDN U12904 ( .A(n16826), .B(o[39]), .Z(n12401) );
  OR U12905 ( .A(n12294), .B(n12293), .Z(n12298) );
  OR U12906 ( .A(n12296), .B(n12295), .Z(n12297) );
  NAND U12907 ( .A(n12298), .B(n12297), .Z(n12402) );
  XOR U12908 ( .A(n12401), .B(n12402), .Z(n12404) );
  XNOR U12909 ( .A(n12403), .B(n12404), .Z(n12633) );
  XNOR U12910 ( .A(n12634), .B(n12633), .Z(n12635) );
  XNOR U12911 ( .A(n12636), .B(n12635), .Z(n12397) );
  NANDN U12912 ( .A(n2976), .B(o[41]), .Z(n12395) );
  OR U12913 ( .A(n12300), .B(n12299), .Z(n12304) );
  OR U12914 ( .A(n12302), .B(n12301), .Z(n12303) );
  NAND U12915 ( .A(n12304), .B(n12303), .Z(n12396) );
  XOR U12916 ( .A(n12395), .B(n12396), .Z(n12398) );
  XNOR U12917 ( .A(n12397), .B(n12398), .Z(n12639) );
  XNOR U12918 ( .A(n12640), .B(n12639), .Z(n12641) );
  XNOR U12919 ( .A(n12642), .B(n12641), .Z(n12391) );
  NANDN U12920 ( .A(n2974), .B(o[43]), .Z(n12389) );
  OR U12921 ( .A(n12306), .B(n12305), .Z(n12310) );
  OR U12922 ( .A(n12308), .B(n12307), .Z(n12309) );
  NAND U12923 ( .A(n12310), .B(n12309), .Z(n12390) );
  XOR U12924 ( .A(n12389), .B(n12390), .Z(n12392) );
  XNOR U12925 ( .A(n12391), .B(n12392), .Z(n12645) );
  XNOR U12926 ( .A(n12646), .B(n12645), .Z(n12647) );
  XNOR U12927 ( .A(n12648), .B(n12647), .Z(n12385) );
  NANDN U12928 ( .A(n2972), .B(o[45]), .Z(n12383) );
  OR U12929 ( .A(n12312), .B(n12311), .Z(n12316) );
  OR U12930 ( .A(n12314), .B(n12313), .Z(n12315) );
  NAND U12931 ( .A(n12316), .B(n12315), .Z(n12384) );
  XOR U12932 ( .A(n12383), .B(n12384), .Z(n12386) );
  XNOR U12933 ( .A(n12385), .B(n12386), .Z(n12651) );
  XNOR U12934 ( .A(n12652), .B(n12651), .Z(n12653) );
  XNOR U12935 ( .A(n12654), .B(n12653), .Z(n12379) );
  NANDN U12936 ( .A(n17145), .B(o[47]), .Z(n12377) );
  OR U12937 ( .A(n12318), .B(n12317), .Z(n12322) );
  OR U12938 ( .A(n12320), .B(n12319), .Z(n12321) );
  NAND U12939 ( .A(n12322), .B(n12321), .Z(n12378) );
  XOR U12940 ( .A(n12377), .B(n12378), .Z(n12380) );
  XNOR U12941 ( .A(n12379), .B(n12380), .Z(n12657) );
  XNOR U12942 ( .A(n12658), .B(n12657), .Z(n12659) );
  XNOR U12943 ( .A(n12660), .B(n12659), .Z(n12373) );
  NANDN U12944 ( .A(n17219), .B(o[49]), .Z(n12371) );
  OR U12945 ( .A(n12324), .B(n12323), .Z(n12328) );
  OR U12946 ( .A(n12326), .B(n12325), .Z(n12327) );
  NAND U12947 ( .A(n12328), .B(n12327), .Z(n12372) );
  XOR U12948 ( .A(n12371), .B(n12372), .Z(n12374) );
  XNOR U12949 ( .A(n12373), .B(n12374), .Z(n12663) );
  XNOR U12950 ( .A(n12664), .B(n12663), .Z(n12665) );
  XNOR U12951 ( .A(n12666), .B(n12665), .Z(n12367) );
  NANDN U12952 ( .A(n17296), .B(o[51]), .Z(n12365) );
  OR U12953 ( .A(n12330), .B(n12329), .Z(n12334) );
  OR U12954 ( .A(n12332), .B(n12331), .Z(n12333) );
  NAND U12955 ( .A(n12334), .B(n12333), .Z(n12366) );
  XOR U12956 ( .A(n12365), .B(n12366), .Z(n12368) );
  XNOR U12957 ( .A(n12367), .B(n12368), .Z(n12669) );
  XNOR U12958 ( .A(n12670), .B(n12669), .Z(n12671) );
  XNOR U12959 ( .A(n12672), .B(n12671), .Z(n12361) );
  NANDN U12960 ( .A(n17375), .B(o[53]), .Z(n12359) );
  OR U12961 ( .A(n12336), .B(n12335), .Z(n12340) );
  OR U12962 ( .A(n12338), .B(n12337), .Z(n12339) );
  NAND U12963 ( .A(n12340), .B(n12339), .Z(n12360) );
  XOR U12964 ( .A(n12359), .B(n12360), .Z(n12362) );
  XNOR U12965 ( .A(n12361), .B(n12362), .Z(n12675) );
  XNOR U12966 ( .A(n12676), .B(n12675), .Z(n12677) );
  AND U12967 ( .A(o[55]), .B(\stack[1][1] ), .Z(n12353) );
  OR U12968 ( .A(n12342), .B(n12341), .Z(n12346) );
  OR U12969 ( .A(n12344), .B(n12343), .Z(n12345) );
  NAND U12970 ( .A(n12346), .B(n12345), .Z(n12354) );
  XNOR U12971 ( .A(n12353), .B(n12354), .Z(n12356) );
  XOR U12972 ( .A(n12355), .B(n12356), .Z(n12347) );
  NANDN U12973 ( .A(n12348), .B(n12347), .Z(n12350) );
  XOR U12974 ( .A(n12348), .B(n12347), .Z(n15318) );
  AND U12975 ( .A(o[56]), .B(\stack[1][0] ), .Z(n15319) );
  OR U12976 ( .A(n15318), .B(n15319), .Z(n12349) );
  AND U12977 ( .A(n12350), .B(n12349), .Z(n12352) );
  OR U12978 ( .A(n12351), .B(n12352), .Z(n12682) );
  XNOR U12979 ( .A(n12352), .B(n12351), .Z(n15279) );
  NANDN U12980 ( .A(n2969), .B(o[56]), .Z(n13014) );
  OR U12981 ( .A(n12354), .B(n12353), .Z(n12358) );
  OR U12982 ( .A(n12356), .B(n12355), .Z(n12357) );
  NAND U12983 ( .A(n12358), .B(n12357), .Z(n13012) );
  NANDN U12984 ( .A(n17375), .B(o[54]), .Z(n13008) );
  NANDN U12985 ( .A(n12360), .B(n12359), .Z(n12364) );
  NANDN U12986 ( .A(n12362), .B(n12361), .Z(n12363) );
  NAND U12987 ( .A(n12364), .B(n12363), .Z(n13006) );
  NANDN U12988 ( .A(n17296), .B(o[52]), .Z(n13002) );
  NANDN U12989 ( .A(n12366), .B(n12365), .Z(n12370) );
  NANDN U12990 ( .A(n12368), .B(n12367), .Z(n12369) );
  NAND U12991 ( .A(n12370), .B(n12369), .Z(n13000) );
  NANDN U12992 ( .A(n17219), .B(o[50]), .Z(n12996) );
  NANDN U12993 ( .A(n12372), .B(n12371), .Z(n12376) );
  NANDN U12994 ( .A(n12374), .B(n12373), .Z(n12375) );
  NAND U12995 ( .A(n12376), .B(n12375), .Z(n12994) );
  NANDN U12996 ( .A(n17145), .B(o[48]), .Z(n12990) );
  NANDN U12997 ( .A(n12378), .B(n12377), .Z(n12382) );
  NANDN U12998 ( .A(n12380), .B(n12379), .Z(n12381) );
  NAND U12999 ( .A(n12382), .B(n12381), .Z(n12988) );
  NANDN U13000 ( .A(n2972), .B(o[46]), .Z(n12984) );
  NANDN U13001 ( .A(n12384), .B(n12383), .Z(n12388) );
  NANDN U13002 ( .A(n12386), .B(n12385), .Z(n12387) );
  NAND U13003 ( .A(n12388), .B(n12387), .Z(n12982) );
  NANDN U13004 ( .A(n2974), .B(o[44]), .Z(n12978) );
  NANDN U13005 ( .A(n12390), .B(n12389), .Z(n12394) );
  NANDN U13006 ( .A(n12392), .B(n12391), .Z(n12393) );
  NAND U13007 ( .A(n12394), .B(n12393), .Z(n12976) );
  NANDN U13008 ( .A(n2976), .B(o[42]), .Z(n12972) );
  NANDN U13009 ( .A(n12396), .B(n12395), .Z(n12400) );
  NANDN U13010 ( .A(n12398), .B(n12397), .Z(n12399) );
  NAND U13011 ( .A(n12400), .B(n12399), .Z(n12970) );
  NANDN U13012 ( .A(n16826), .B(o[40]), .Z(n12966) );
  NANDN U13013 ( .A(n12402), .B(n12401), .Z(n12406) );
  NANDN U13014 ( .A(n12404), .B(n12403), .Z(n12405) );
  NAND U13015 ( .A(n12406), .B(n12405), .Z(n12964) );
  NANDN U13016 ( .A(n16746), .B(o[38]), .Z(n12960) );
  NANDN U13017 ( .A(n12408), .B(n12407), .Z(n12412) );
  NANDN U13018 ( .A(n12410), .B(n12409), .Z(n12411) );
  NAND U13019 ( .A(n12412), .B(n12411), .Z(n12958) );
  NANDN U13020 ( .A(n2978), .B(o[36]), .Z(n12954) );
  NANDN U13021 ( .A(n12414), .B(n12413), .Z(n12418) );
  NANDN U13022 ( .A(n12416), .B(n12415), .Z(n12417) );
  NAND U13023 ( .A(n12418), .B(n12417), .Z(n12952) );
  NANDN U13024 ( .A(n2980), .B(o[34]), .Z(n12948) );
  NANDN U13025 ( .A(n12420), .B(n12419), .Z(n12424) );
  NANDN U13026 ( .A(n12422), .B(n12421), .Z(n12423) );
  NAND U13027 ( .A(n12424), .B(n12423), .Z(n12946) );
  NANDN U13028 ( .A(n2982), .B(o[32]), .Z(n12942) );
  NANDN U13029 ( .A(n12426), .B(n12425), .Z(n12430) );
  NANDN U13030 ( .A(n12428), .B(n12427), .Z(n12429) );
  NAND U13031 ( .A(n12430), .B(n12429), .Z(n12940) );
  NANDN U13032 ( .A(n2984), .B(o[30]), .Z(n12936) );
  NANDN U13033 ( .A(n12432), .B(n12431), .Z(n12436) );
  NANDN U13034 ( .A(n12434), .B(n12433), .Z(n12435) );
  NAND U13035 ( .A(n12436), .B(n12435), .Z(n12934) );
  AND U13036 ( .A(\stack[1][29] ), .B(o[28]), .Z(n12770) );
  OR U13037 ( .A(n12438), .B(n12437), .Z(n12442) );
  OR U13038 ( .A(n12440), .B(n12439), .Z(n12441) );
  AND U13039 ( .A(n12442), .B(n12441), .Z(n12767) );
  OR U13040 ( .A(n12444), .B(n12443), .Z(n12448) );
  NANDN U13041 ( .A(n12446), .B(n12445), .Z(n12447) );
  AND U13042 ( .A(n12448), .B(n12447), .Z(n12927) );
  AND U13043 ( .A(o[27]), .B(\stack[1][30] ), .Z(n12928) );
  XNOR U13044 ( .A(n12927), .B(n12928), .Z(n12930) );
  OR U13045 ( .A(n12450), .B(n12449), .Z(n12454) );
  OR U13046 ( .A(n12452), .B(n12451), .Z(n12453) );
  NAND U13047 ( .A(n12454), .B(n12453), .Z(n12780) );
  ANDN U13048 ( .B(o[25]), .A(n2989), .Z(n12779) );
  XOR U13049 ( .A(n12780), .B(n12779), .Z(n12781) );
  NANDN U13050 ( .A(n3018), .B(\stack[1][33] ), .Z(n12788) );
  OR U13051 ( .A(n12456), .B(n12455), .Z(n12460) );
  OR U13052 ( .A(n12458), .B(n12457), .Z(n12459) );
  NAND U13053 ( .A(n12460), .B(n12459), .Z(n12786) );
  NANDN U13054 ( .A(n3016), .B(\stack[1][35] ), .Z(n12924) );
  NANDN U13055 ( .A(n12462), .B(n12461), .Z(n12466) );
  OR U13056 ( .A(n12464), .B(n12463), .Z(n12465) );
  NAND U13057 ( .A(n12466), .B(n12465), .Z(n12922) );
  NANDN U13058 ( .A(n3014), .B(\stack[1][37] ), .Z(n12806) );
  OR U13059 ( .A(n12468), .B(n12467), .Z(n12472) );
  OR U13060 ( .A(n12470), .B(n12469), .Z(n12471) );
  NAND U13061 ( .A(n12472), .B(n12471), .Z(n12804) );
  NANDN U13062 ( .A(n3013), .B(\stack[1][38] ), .Z(n12811) );
  OR U13063 ( .A(n12474), .B(n12473), .Z(n12478) );
  OR U13064 ( .A(n12476), .B(n12475), .Z(n12477) );
  AND U13065 ( .A(n12478), .B(n12477), .Z(n12810) );
  OR U13066 ( .A(n12480), .B(n12479), .Z(n12484) );
  NAND U13067 ( .A(n12482), .B(n12481), .Z(n12483) );
  AND U13068 ( .A(n12484), .B(n12483), .Z(n12912) );
  OR U13069 ( .A(n12486), .B(n12485), .Z(n12490) );
  OR U13070 ( .A(n12488), .B(n12487), .Z(n12489) );
  AND U13071 ( .A(n12490), .B(n12489), .Z(n12815) );
  NANDN U13072 ( .A(n3010), .B(\stack[1][41] ), .Z(n12816) );
  XOR U13073 ( .A(n12815), .B(n12816), .Z(n12818) );
  NANDN U13074 ( .A(n3009), .B(\stack[1][42] ), .Z(n12824) );
  OR U13075 ( .A(n12492), .B(n12491), .Z(n12496) );
  OR U13076 ( .A(n12494), .B(n12493), .Z(n12495) );
  AND U13077 ( .A(n12496), .B(n12495), .Z(n12899) );
  NANDN U13078 ( .A(n12498), .B(n12497), .Z(n12502) );
  NANDN U13079 ( .A(n12500), .B(n12499), .Z(n12501) );
  NAND U13080 ( .A(n12502), .B(n12501), .Z(n12828) );
  AND U13081 ( .A(\stack[1][46] ), .B(o[11]), .Z(n12836) );
  OR U13082 ( .A(n12504), .B(n12503), .Z(n12508) );
  NANDN U13083 ( .A(n12506), .B(n12505), .Z(n12507) );
  AND U13084 ( .A(n12508), .B(n12507), .Z(n12833) );
  AND U13085 ( .A(\stack[1][47] ), .B(o[10]), .Z(n12842) );
  AND U13086 ( .A(\stack[1][48] ), .B(o[9]), .Z(n12893) );
  NANDN U13087 ( .A(n12510), .B(n12509), .Z(n12514) );
  NAND U13088 ( .A(n12512), .B(n12511), .Z(n12513) );
  AND U13089 ( .A(n12514), .B(n12513), .Z(n12882) );
  AND U13090 ( .A(\stack[1][52] ), .B(o[5]), .Z(n12876) );
  OR U13091 ( .A(n12516), .B(n12515), .Z(n12520) );
  NANDN U13092 ( .A(n12518), .B(n12517), .Z(n12519) );
  AND U13093 ( .A(n12520), .B(n12519), .Z(n12873) );
  ANDN U13094 ( .B(\stack[1][53] ), .A(n2998), .Z(n12854) );
  ANDN U13095 ( .B(\stack[1][54] ), .A(n2997), .Z(n12870) );
  NANDN U13096 ( .A(n12521), .B(n12857), .Z(n12522) );
  AND U13097 ( .A(n12523), .B(n12522), .Z(n12527) );
  OR U13098 ( .A(n12525), .B(n12524), .Z(n12526) );
  AND U13099 ( .A(n12527), .B(n12526), .Z(n12867) );
  AND U13100 ( .A(\stack[1][57] ), .B(o[1]), .Z(n12865) );
  ANDN U13101 ( .B(n12865), .A(n12528), .Z(n13203) );
  XNOR U13102 ( .A(n13203), .B(n12857), .Z(n12530) );
  NAND U13103 ( .A(o[0]), .B(\stack[1][57] ), .Z(n12864) );
  NANDN U13104 ( .A(n12529), .B(n12864), .Z(n12859) );
  NAND U13105 ( .A(n12530), .B(n12859), .Z(n12861) );
  ANDN U13106 ( .B(\stack[1][55] ), .A(n2996), .Z(n12860) );
  XNOR U13107 ( .A(n12861), .B(n12860), .Z(n12868) );
  XOR U13108 ( .A(n12867), .B(n12868), .Z(n12869) );
  XOR U13109 ( .A(n12870), .B(n12869), .Z(n12852) );
  OR U13110 ( .A(n12532), .B(n12531), .Z(n12536) );
  NANDN U13111 ( .A(n12534), .B(n12533), .Z(n12535) );
  AND U13112 ( .A(n12536), .B(n12535), .Z(n12851) );
  XOR U13113 ( .A(n12852), .B(n12851), .Z(n12853) );
  XOR U13114 ( .A(n12854), .B(n12853), .Z(n12874) );
  XNOR U13115 ( .A(n12873), .B(n12874), .Z(n12875) );
  OR U13116 ( .A(n12538), .B(n12537), .Z(n12542) );
  OR U13117 ( .A(n12540), .B(n12539), .Z(n12541) );
  NAND U13118 ( .A(n12542), .B(n12541), .Z(n12846) );
  IV U13119 ( .A(\stack[1][51] ), .Z(n15507) );
  ANDN U13120 ( .B(o[6]), .A(n15507), .Z(n12845) );
  XNOR U13121 ( .A(n12846), .B(n12845), .Z(n12848) );
  XNOR U13122 ( .A(n12847), .B(n12848), .Z(n12880) );
  ANDN U13123 ( .B(o[7]), .A(n15546), .Z(n12879) );
  XOR U13124 ( .A(n12880), .B(n12879), .Z(n12881) );
  NANDN U13125 ( .A(n12544), .B(n12543), .Z(n12548) );
  OR U13126 ( .A(n12546), .B(n12545), .Z(n12547) );
  AND U13127 ( .A(n12548), .B(n12547), .Z(n12885) );
  XNOR U13128 ( .A(n12886), .B(n12885), .Z(n12888) );
  ANDN U13129 ( .B(\stack[1][49] ), .A(n3002), .Z(n12887) );
  XNOR U13130 ( .A(n12888), .B(n12887), .Z(n12891) );
  OR U13131 ( .A(n12550), .B(n12549), .Z(n12554) );
  NANDN U13132 ( .A(n12552), .B(n12551), .Z(n12553) );
  NAND U13133 ( .A(n12554), .B(n12553), .Z(n12892) );
  XNOR U13134 ( .A(n12891), .B(n12892), .Z(n12894) );
  XNOR U13135 ( .A(n12893), .B(n12894), .Z(n12840) );
  OR U13136 ( .A(n12556), .B(n12555), .Z(n12560) );
  OR U13137 ( .A(n12558), .B(n12557), .Z(n12559) );
  AND U13138 ( .A(n12560), .B(n12559), .Z(n12839) );
  XOR U13139 ( .A(n12840), .B(n12839), .Z(n12841) );
  XOR U13140 ( .A(n12842), .B(n12841), .Z(n12834) );
  XNOR U13141 ( .A(n12833), .B(n12834), .Z(n12835) );
  XOR U13142 ( .A(n12828), .B(n12827), .Z(n12830) );
  ANDN U13143 ( .B(o[12]), .A(n15740), .Z(n12829) );
  XOR U13144 ( .A(n12830), .B(n12829), .Z(n12898) );
  ANDN U13145 ( .B(o[13]), .A(n15779), .Z(n12897) );
  XOR U13146 ( .A(n12898), .B(n12897), .Z(n12900) );
  XNOR U13147 ( .A(n12899), .B(n12900), .Z(n12904) );
  NANDN U13148 ( .A(n12562), .B(n12561), .Z(n12566) );
  OR U13149 ( .A(n12564), .B(n12563), .Z(n12565) );
  AND U13150 ( .A(n12566), .B(n12565), .Z(n12903) );
  XNOR U13151 ( .A(n12904), .B(n12903), .Z(n12906) );
  ANDN U13152 ( .B(o[14]), .A(n15818), .Z(n12905) );
  XOR U13153 ( .A(n12906), .B(n12905), .Z(n12822) );
  OR U13154 ( .A(n12568), .B(n12567), .Z(n12572) );
  NANDN U13155 ( .A(n12570), .B(n12569), .Z(n12571) );
  AND U13156 ( .A(n12572), .B(n12571), .Z(n12821) );
  XNOR U13157 ( .A(n12822), .B(n12821), .Z(n12823) );
  XOR U13158 ( .A(n12824), .B(n12823), .Z(n12817) );
  XNOR U13159 ( .A(n12818), .B(n12817), .Z(n12910) );
  ANDN U13160 ( .B(o[17]), .A(n15935), .Z(n12909) );
  XOR U13161 ( .A(n12910), .B(n12909), .Z(n12911) );
  OR U13162 ( .A(n12574), .B(n12573), .Z(n12578) );
  NANDN U13163 ( .A(n12576), .B(n12575), .Z(n12577) );
  AND U13164 ( .A(n12578), .B(n12577), .Z(n12915) );
  XNOR U13165 ( .A(n12916), .B(n12915), .Z(n12918) );
  ANDN U13166 ( .B(\stack[1][39] ), .A(n3012), .Z(n12917) );
  XOR U13167 ( .A(n12918), .B(n12917), .Z(n12809) );
  XOR U13168 ( .A(n12810), .B(n12809), .Z(n12812) );
  XNOR U13169 ( .A(n12811), .B(n12812), .Z(n12803) );
  XNOR U13170 ( .A(n12804), .B(n12803), .Z(n12805) );
  XNOR U13171 ( .A(n12806), .B(n12805), .Z(n12799) );
  OR U13172 ( .A(n12580), .B(n12579), .Z(n12584) );
  OR U13173 ( .A(n12582), .B(n12581), .Z(n12583) );
  AND U13174 ( .A(n12584), .B(n12583), .Z(n12798) );
  NANDN U13175 ( .A(n2993), .B(o[21]), .Z(n12797) );
  XOR U13176 ( .A(n12798), .B(n12797), .Z(n12800) );
  XNOR U13177 ( .A(n12799), .B(n12800), .Z(n12921) );
  XNOR U13178 ( .A(n12922), .B(n12921), .Z(n12923) );
  XNOR U13179 ( .A(n12924), .B(n12923), .Z(n12793) );
  AND U13180 ( .A(\stack[1][34] ), .B(o[23]), .Z(n12791) );
  NANDN U13181 ( .A(n12586), .B(n12585), .Z(n12590) );
  NANDN U13182 ( .A(n12588), .B(n12587), .Z(n12589) );
  NAND U13183 ( .A(n12590), .B(n12589), .Z(n12792) );
  XNOR U13184 ( .A(n12791), .B(n12792), .Z(n12794) );
  XNOR U13185 ( .A(n12793), .B(n12794), .Z(n12785) );
  XNOR U13186 ( .A(n12786), .B(n12785), .Z(n12787) );
  XNOR U13187 ( .A(n12788), .B(n12787), .Z(n12782) );
  OR U13188 ( .A(n12592), .B(n12591), .Z(n12596) );
  OR U13189 ( .A(n12594), .B(n12593), .Z(n12595) );
  AND U13190 ( .A(n12596), .B(n12595), .Z(n12774) );
  XNOR U13191 ( .A(n12773), .B(n12774), .Z(n12776) );
  AND U13192 ( .A(\stack[1][31] ), .B(o[26]), .Z(n12775) );
  XOR U13193 ( .A(n12776), .B(n12775), .Z(n12929) );
  XOR U13194 ( .A(n12930), .B(n12929), .Z(n12768) );
  XOR U13195 ( .A(n12767), .B(n12768), .Z(n12769) );
  XOR U13196 ( .A(n12770), .B(n12769), .Z(n12764) );
  AND U13197 ( .A(o[29]), .B(\stack[1][28] ), .Z(n12761) );
  OR U13198 ( .A(n12598), .B(n12597), .Z(n12602) );
  IV U13199 ( .A(n12599), .Z(n16399) );
  OR U13200 ( .A(n12600), .B(n16399), .Z(n12601) );
  NAND U13201 ( .A(n12602), .B(n12601), .Z(n12762) );
  XNOR U13202 ( .A(n12761), .B(n12762), .Z(n12763) );
  XOR U13203 ( .A(n12764), .B(n12763), .Z(n12933) );
  XNOR U13204 ( .A(n12934), .B(n12933), .Z(n12935) );
  XNOR U13205 ( .A(n12936), .B(n12935), .Z(n12757) );
  NANDN U13206 ( .A(n2983), .B(o[31]), .Z(n12755) );
  OR U13207 ( .A(n12604), .B(n12603), .Z(n12608) );
  OR U13208 ( .A(n12606), .B(n12605), .Z(n12607) );
  NAND U13209 ( .A(n12608), .B(n12607), .Z(n12756) );
  XOR U13210 ( .A(n12755), .B(n12756), .Z(n12758) );
  XNOR U13211 ( .A(n12757), .B(n12758), .Z(n12939) );
  XNOR U13212 ( .A(n12940), .B(n12939), .Z(n12941) );
  XNOR U13213 ( .A(n12942), .B(n12941), .Z(n12751) );
  NANDN U13214 ( .A(n2981), .B(o[33]), .Z(n12749) );
  OR U13215 ( .A(n12610), .B(n12609), .Z(n12614) );
  OR U13216 ( .A(n12612), .B(n12611), .Z(n12613) );
  NAND U13217 ( .A(n12614), .B(n12613), .Z(n12750) );
  XOR U13218 ( .A(n12749), .B(n12750), .Z(n12752) );
  XNOR U13219 ( .A(n12751), .B(n12752), .Z(n12945) );
  XNOR U13220 ( .A(n12946), .B(n12945), .Z(n12947) );
  XNOR U13221 ( .A(n12948), .B(n12947), .Z(n12745) );
  NANDN U13222 ( .A(n2979), .B(o[35]), .Z(n12743) );
  OR U13223 ( .A(n12616), .B(n12615), .Z(n12620) );
  OR U13224 ( .A(n12618), .B(n12617), .Z(n12619) );
  NAND U13225 ( .A(n12620), .B(n12619), .Z(n12744) );
  XOR U13226 ( .A(n12743), .B(n12744), .Z(n12746) );
  XNOR U13227 ( .A(n12745), .B(n12746), .Z(n12951) );
  XNOR U13228 ( .A(n12952), .B(n12951), .Z(n12953) );
  XNOR U13229 ( .A(n12954), .B(n12953), .Z(n12739) );
  NANDN U13230 ( .A(n16712), .B(o[37]), .Z(n12737) );
  OR U13231 ( .A(n12622), .B(n12621), .Z(n12626) );
  OR U13232 ( .A(n12624), .B(n12623), .Z(n12625) );
  NAND U13233 ( .A(n12626), .B(n12625), .Z(n12738) );
  XOR U13234 ( .A(n12737), .B(n12738), .Z(n12740) );
  XNOR U13235 ( .A(n12739), .B(n12740), .Z(n12957) );
  XNOR U13236 ( .A(n12958), .B(n12957), .Z(n12959) );
  XNOR U13237 ( .A(n12960), .B(n12959), .Z(n12733) );
  NANDN U13238 ( .A(n16786), .B(o[39]), .Z(n12731) );
  OR U13239 ( .A(n12628), .B(n12627), .Z(n12632) );
  OR U13240 ( .A(n12630), .B(n12629), .Z(n12631) );
  NAND U13241 ( .A(n12632), .B(n12631), .Z(n12732) );
  XOR U13242 ( .A(n12731), .B(n12732), .Z(n12734) );
  XNOR U13243 ( .A(n12733), .B(n12734), .Z(n12963) );
  XNOR U13244 ( .A(n12964), .B(n12963), .Z(n12965) );
  XNOR U13245 ( .A(n12966), .B(n12965), .Z(n12727) );
  NANDN U13246 ( .A(n2977), .B(o[41]), .Z(n12725) );
  OR U13247 ( .A(n12634), .B(n12633), .Z(n12638) );
  OR U13248 ( .A(n12636), .B(n12635), .Z(n12637) );
  NAND U13249 ( .A(n12638), .B(n12637), .Z(n12726) );
  XOR U13250 ( .A(n12725), .B(n12726), .Z(n12728) );
  XNOR U13251 ( .A(n12727), .B(n12728), .Z(n12969) );
  XNOR U13252 ( .A(n12970), .B(n12969), .Z(n12971) );
  XNOR U13253 ( .A(n12972), .B(n12971), .Z(n12721) );
  NANDN U13254 ( .A(n2975), .B(o[43]), .Z(n12719) );
  OR U13255 ( .A(n12640), .B(n12639), .Z(n12644) );
  OR U13256 ( .A(n12642), .B(n12641), .Z(n12643) );
  NAND U13257 ( .A(n12644), .B(n12643), .Z(n12720) );
  XOR U13258 ( .A(n12719), .B(n12720), .Z(n12722) );
  XNOR U13259 ( .A(n12721), .B(n12722), .Z(n12975) );
  XNOR U13260 ( .A(n12976), .B(n12975), .Z(n12977) );
  XNOR U13261 ( .A(n12978), .B(n12977), .Z(n12715) );
  NANDN U13262 ( .A(n2973), .B(o[45]), .Z(n12713) );
  OR U13263 ( .A(n12646), .B(n12645), .Z(n12650) );
  OR U13264 ( .A(n12648), .B(n12647), .Z(n12649) );
  NAND U13265 ( .A(n12650), .B(n12649), .Z(n12714) );
  XOR U13266 ( .A(n12713), .B(n12714), .Z(n12716) );
  XNOR U13267 ( .A(n12715), .B(n12716), .Z(n12981) );
  XNOR U13268 ( .A(n12982), .B(n12981), .Z(n12983) );
  XNOR U13269 ( .A(n12984), .B(n12983), .Z(n12709) );
  NANDN U13270 ( .A(n17101), .B(o[47]), .Z(n12707) );
  OR U13271 ( .A(n12652), .B(n12651), .Z(n12656) );
  OR U13272 ( .A(n12654), .B(n12653), .Z(n12655) );
  NAND U13273 ( .A(n12656), .B(n12655), .Z(n12708) );
  XOR U13274 ( .A(n12707), .B(n12708), .Z(n12710) );
  XNOR U13275 ( .A(n12709), .B(n12710), .Z(n12987) );
  XNOR U13276 ( .A(n12988), .B(n12987), .Z(n12989) );
  XNOR U13277 ( .A(n12990), .B(n12989), .Z(n12703) );
  NANDN U13278 ( .A(n17179), .B(o[49]), .Z(n12701) );
  OR U13279 ( .A(n12658), .B(n12657), .Z(n12662) );
  OR U13280 ( .A(n12660), .B(n12659), .Z(n12661) );
  NAND U13281 ( .A(n12662), .B(n12661), .Z(n12702) );
  XOR U13282 ( .A(n12701), .B(n12702), .Z(n12704) );
  XNOR U13283 ( .A(n12703), .B(n12704), .Z(n12993) );
  XNOR U13284 ( .A(n12994), .B(n12993), .Z(n12995) );
  XNOR U13285 ( .A(n12996), .B(n12995), .Z(n12697) );
  NANDN U13286 ( .A(n17256), .B(o[51]), .Z(n12695) );
  OR U13287 ( .A(n12664), .B(n12663), .Z(n12668) );
  OR U13288 ( .A(n12666), .B(n12665), .Z(n12667) );
  NAND U13289 ( .A(n12668), .B(n12667), .Z(n12696) );
  XOR U13290 ( .A(n12695), .B(n12696), .Z(n12698) );
  XNOR U13291 ( .A(n12697), .B(n12698), .Z(n12999) );
  XNOR U13292 ( .A(n13000), .B(n12999), .Z(n13001) );
  XNOR U13293 ( .A(n13002), .B(n13001), .Z(n12691) );
  AND U13294 ( .A(o[53]), .B(\stack[1][4] ), .Z(n12689) );
  OR U13295 ( .A(n12670), .B(n12669), .Z(n12674) );
  OR U13296 ( .A(n12672), .B(n12671), .Z(n12673) );
  NAND U13297 ( .A(n12674), .B(n12673), .Z(n12690) );
  XNOR U13298 ( .A(n12689), .B(n12690), .Z(n12692) );
  XNOR U13299 ( .A(n12691), .B(n12692), .Z(n13005) );
  XNOR U13300 ( .A(n13006), .B(n13005), .Z(n13007) );
  XOR U13301 ( .A(n13008), .B(n13007), .Z(n12686) );
  AND U13302 ( .A(o[55]), .B(\stack[1][2] ), .Z(n12683) );
  OR U13303 ( .A(n12676), .B(n12675), .Z(n12680) );
  OR U13304 ( .A(n12678), .B(n12677), .Z(n12679) );
  NAND U13305 ( .A(n12680), .B(n12679), .Z(n12684) );
  XOR U13306 ( .A(n12683), .B(n12684), .Z(n12685) );
  XNOR U13307 ( .A(n12686), .B(n12685), .Z(n13011) );
  XNOR U13308 ( .A(n13012), .B(n13011), .Z(n13013) );
  XOR U13309 ( .A(n13014), .B(n13013), .Z(n15280) );
  OR U13310 ( .A(n15279), .B(n15280), .Z(n12681) );
  AND U13311 ( .A(n12682), .B(n12681), .Z(n13018) );
  NANDN U13312 ( .A(n2970), .B(o[56]), .Z(n13360) );
  OR U13313 ( .A(n12684), .B(n12683), .Z(n12688) );
  NANDN U13314 ( .A(n12686), .B(n12685), .Z(n12687) );
  NAND U13315 ( .A(n12688), .B(n12687), .Z(n13358) );
  NANDN U13316 ( .A(n2971), .B(o[54]), .Z(n13354) );
  OR U13317 ( .A(n12690), .B(n12689), .Z(n12694) );
  NANDN U13318 ( .A(n12692), .B(n12691), .Z(n12693) );
  NAND U13319 ( .A(n12694), .B(n12693), .Z(n13352) );
  NANDN U13320 ( .A(n17256), .B(o[52]), .Z(n13348) );
  NANDN U13321 ( .A(n12696), .B(n12695), .Z(n12700) );
  NANDN U13322 ( .A(n12698), .B(n12697), .Z(n12699) );
  NAND U13323 ( .A(n12700), .B(n12699), .Z(n13346) );
  NANDN U13324 ( .A(n17179), .B(o[50]), .Z(n13342) );
  NANDN U13325 ( .A(n12702), .B(n12701), .Z(n12706) );
  NANDN U13326 ( .A(n12704), .B(n12703), .Z(n12705) );
  NAND U13327 ( .A(n12706), .B(n12705), .Z(n13340) );
  NANDN U13328 ( .A(n17101), .B(o[48]), .Z(n13336) );
  NANDN U13329 ( .A(n12708), .B(n12707), .Z(n12712) );
  NANDN U13330 ( .A(n12710), .B(n12709), .Z(n12711) );
  NAND U13331 ( .A(n12712), .B(n12711), .Z(n13334) );
  NANDN U13332 ( .A(n2973), .B(o[46]), .Z(n13330) );
  NANDN U13333 ( .A(n12714), .B(n12713), .Z(n12718) );
  NANDN U13334 ( .A(n12716), .B(n12715), .Z(n12717) );
  NAND U13335 ( .A(n12718), .B(n12717), .Z(n13328) );
  NANDN U13336 ( .A(n2975), .B(o[44]), .Z(n13324) );
  NANDN U13337 ( .A(n12720), .B(n12719), .Z(n12724) );
  NANDN U13338 ( .A(n12722), .B(n12721), .Z(n12723) );
  NAND U13339 ( .A(n12724), .B(n12723), .Z(n13322) );
  NANDN U13340 ( .A(n2977), .B(o[42]), .Z(n13318) );
  NANDN U13341 ( .A(n12726), .B(n12725), .Z(n12730) );
  NANDN U13342 ( .A(n12728), .B(n12727), .Z(n12729) );
  NAND U13343 ( .A(n12730), .B(n12729), .Z(n13316) );
  NANDN U13344 ( .A(n16786), .B(o[40]), .Z(n13312) );
  NANDN U13345 ( .A(n12732), .B(n12731), .Z(n12736) );
  NANDN U13346 ( .A(n12734), .B(n12733), .Z(n12735) );
  NAND U13347 ( .A(n12736), .B(n12735), .Z(n13310) );
  NANDN U13348 ( .A(n16712), .B(o[38]), .Z(n13306) );
  NANDN U13349 ( .A(n12738), .B(n12737), .Z(n12742) );
  NANDN U13350 ( .A(n12740), .B(n12739), .Z(n12741) );
  NAND U13351 ( .A(n12742), .B(n12741), .Z(n13304) );
  NANDN U13352 ( .A(n2979), .B(o[36]), .Z(n13300) );
  NANDN U13353 ( .A(n12744), .B(n12743), .Z(n12748) );
  NANDN U13354 ( .A(n12746), .B(n12745), .Z(n12747) );
  NAND U13355 ( .A(n12748), .B(n12747), .Z(n13298) );
  NANDN U13356 ( .A(n2981), .B(o[34]), .Z(n13294) );
  NANDN U13357 ( .A(n12750), .B(n12749), .Z(n12754) );
  NANDN U13358 ( .A(n12752), .B(n12751), .Z(n12753) );
  NAND U13359 ( .A(n12754), .B(n12753), .Z(n13292) );
  NANDN U13360 ( .A(n2983), .B(o[32]), .Z(n13288) );
  NANDN U13361 ( .A(n12756), .B(n12755), .Z(n12760) );
  NANDN U13362 ( .A(n12758), .B(n12757), .Z(n12759) );
  NAND U13363 ( .A(n12760), .B(n12759), .Z(n13286) );
  AND U13364 ( .A(o[30]), .B(\stack[1][28] ), .Z(n13110) );
  OR U13365 ( .A(n12762), .B(n12761), .Z(n12766) );
  OR U13366 ( .A(n12764), .B(n12763), .Z(n12765) );
  AND U13367 ( .A(n12766), .B(n12765), .Z(n13107) );
  AND U13368 ( .A(o[29]), .B(\stack[1][29] ), .Z(n13279) );
  OR U13369 ( .A(n12768), .B(n12767), .Z(n12772) );
  NANDN U13370 ( .A(n12770), .B(n12769), .Z(n12771) );
  AND U13371 ( .A(n12772), .B(n12771), .Z(n13280) );
  XNOR U13372 ( .A(n13279), .B(n13280), .Z(n13282) );
  OR U13373 ( .A(n12774), .B(n12773), .Z(n12778) );
  OR U13374 ( .A(n12776), .B(n12775), .Z(n12777) );
  NAND U13375 ( .A(n12778), .B(n12777), .Z(n13120) );
  ANDN U13376 ( .B(o[27]), .A(n2988), .Z(n13119) );
  XNOR U13377 ( .A(n13120), .B(n13119), .Z(n13121) );
  NANDN U13378 ( .A(n3020), .B(\stack[1][32] ), .Z(n13276) );
  NANDN U13379 ( .A(n12780), .B(n12779), .Z(n12784) );
  OR U13380 ( .A(n12782), .B(n12781), .Z(n12783) );
  AND U13381 ( .A(n12784), .B(n12783), .Z(n13273) );
  AND U13382 ( .A(\stack[1][33] ), .B(o[25]), .Z(n13125) );
  OR U13383 ( .A(n12786), .B(n12785), .Z(n12790) );
  OR U13384 ( .A(n12788), .B(n12787), .Z(n12789) );
  NAND U13385 ( .A(n12790), .B(n12789), .Z(n13126) );
  XNOR U13386 ( .A(n13125), .B(n13126), .Z(n13128) );
  OR U13387 ( .A(n12792), .B(n12791), .Z(n12796) );
  NANDN U13388 ( .A(n12794), .B(n12793), .Z(n12795) );
  AND U13389 ( .A(n12796), .B(n12795), .Z(n13131) );
  NANDN U13390 ( .A(n12798), .B(n12797), .Z(n12802) );
  NANDN U13391 ( .A(n12800), .B(n12799), .Z(n12801) );
  NAND U13392 ( .A(n12802), .B(n12801), .Z(n13268) );
  AND U13393 ( .A(\stack[1][37] ), .B(o[21]), .Z(n13143) );
  OR U13394 ( .A(n12804), .B(n12803), .Z(n12808) );
  OR U13395 ( .A(n12806), .B(n12805), .Z(n12807) );
  NAND U13396 ( .A(n12808), .B(n12807), .Z(n13144) );
  XNOR U13397 ( .A(n13143), .B(n13144), .Z(n13146) );
  NANDN U13398 ( .A(n3014), .B(\stack[1][38] ), .Z(n13151) );
  NANDN U13399 ( .A(n12810), .B(n12809), .Z(n12814) );
  NANDN U13400 ( .A(n12812), .B(n12811), .Z(n12813) );
  AND U13401 ( .A(n12814), .B(n12813), .Z(n13149) );
  NANDN U13402 ( .A(n3013), .B(\stack[1][39] ), .Z(n13262) );
  OR U13403 ( .A(n12816), .B(n12815), .Z(n12820) );
  NAND U13404 ( .A(n12818), .B(n12817), .Z(n12819) );
  AND U13405 ( .A(n12820), .B(n12819), .Z(n13258) );
  OR U13406 ( .A(n12822), .B(n12821), .Z(n12826) );
  OR U13407 ( .A(n12824), .B(n12823), .Z(n12825) );
  AND U13408 ( .A(n12826), .B(n12825), .Z(n13161) );
  NANDN U13409 ( .A(n3010), .B(\stack[1][42] ), .Z(n13162) );
  XOR U13410 ( .A(n13161), .B(n13162), .Z(n13164) );
  NANDN U13411 ( .A(n3009), .B(\stack[1][43] ), .Z(n13170) );
  NANDN U13412 ( .A(n12828), .B(n12827), .Z(n12832) );
  NANDN U13413 ( .A(n12830), .B(n12829), .Z(n12831) );
  AND U13414 ( .A(n12832), .B(n12831), .Z(n13245) );
  OR U13415 ( .A(n12834), .B(n12833), .Z(n12838) );
  OR U13416 ( .A(n12836), .B(n12835), .Z(n12837) );
  NAND U13417 ( .A(n12838), .B(n12837), .Z(n13174) );
  AND U13418 ( .A(\stack[1][47] ), .B(o[11]), .Z(n13182) );
  OR U13419 ( .A(n12840), .B(n12839), .Z(n12844) );
  NANDN U13420 ( .A(n12842), .B(n12841), .Z(n12843) );
  AND U13421 ( .A(n12844), .B(n12843), .Z(n13179) );
  AND U13422 ( .A(\stack[1][48] ), .B(o[10]), .Z(n13188) );
  ANDN U13423 ( .B(\stack[1][49] ), .A(n3003), .Z(n13239) );
  NANDN U13424 ( .A(n12846), .B(n12845), .Z(n12850) );
  NAND U13425 ( .A(n12848), .B(n12847), .Z(n12849) );
  AND U13426 ( .A(n12850), .B(n12849), .Z(n13228) );
  ANDN U13427 ( .B(\stack[1][53] ), .A(n2999), .Z(n13222) );
  OR U13428 ( .A(n12852), .B(n12851), .Z(n12856) );
  NANDN U13429 ( .A(n12854), .B(n12853), .Z(n12855) );
  AND U13430 ( .A(n12856), .B(n12855), .Z(n13219) );
  ANDN U13431 ( .B(\stack[1][54] ), .A(n2998), .Z(n13200) );
  ANDN U13432 ( .B(\stack[1][55] ), .A(n2997), .Z(n13216) );
  NANDN U13433 ( .A(n12857), .B(n13203), .Z(n12858) );
  AND U13434 ( .A(n12859), .B(n12858), .Z(n12863) );
  OR U13435 ( .A(n12861), .B(n12860), .Z(n12862) );
  AND U13436 ( .A(n12863), .B(n12862), .Z(n13213) );
  AND U13437 ( .A(\stack[1][58] ), .B(o[1]), .Z(n13211) );
  ANDN U13438 ( .B(n13211), .A(n12864), .Z(n13533) );
  XNOR U13439 ( .A(n13533), .B(n13203), .Z(n12866) );
  NAND U13440 ( .A(\stack[1][58] ), .B(o[0]), .Z(n13210) );
  NANDN U13441 ( .A(n12865), .B(n13210), .Z(n13205) );
  NAND U13442 ( .A(n12866), .B(n13205), .Z(n13207) );
  AND U13443 ( .A(\stack[1][56] ), .B(o[2]), .Z(n13206) );
  XNOR U13444 ( .A(n13207), .B(n13206), .Z(n13214) );
  XOR U13445 ( .A(n13213), .B(n13214), .Z(n13215) );
  XOR U13446 ( .A(n13216), .B(n13215), .Z(n13198) );
  OR U13447 ( .A(n12868), .B(n12867), .Z(n12872) );
  NANDN U13448 ( .A(n12870), .B(n12869), .Z(n12871) );
  AND U13449 ( .A(n12872), .B(n12871), .Z(n13197) );
  XOR U13450 ( .A(n13198), .B(n13197), .Z(n13199) );
  XOR U13451 ( .A(n13200), .B(n13199), .Z(n13220) );
  XNOR U13452 ( .A(n13219), .B(n13220), .Z(n13221) );
  OR U13453 ( .A(n12874), .B(n12873), .Z(n12878) );
  OR U13454 ( .A(n12876), .B(n12875), .Z(n12877) );
  NAND U13455 ( .A(n12878), .B(n12877), .Z(n13192) );
  IV U13456 ( .A(\stack[1][52] ), .Z(n15468) );
  ANDN U13457 ( .B(o[6]), .A(n15468), .Z(n13191) );
  XNOR U13458 ( .A(n13192), .B(n13191), .Z(n13194) );
  XNOR U13459 ( .A(n13193), .B(n13194), .Z(n13226) );
  ANDN U13460 ( .B(o[7]), .A(n15507), .Z(n13225) );
  XOR U13461 ( .A(n13226), .B(n13225), .Z(n13227) );
  NANDN U13462 ( .A(n12880), .B(n12879), .Z(n12884) );
  OR U13463 ( .A(n12882), .B(n12881), .Z(n12883) );
  AND U13464 ( .A(n12884), .B(n12883), .Z(n13231) );
  XNOR U13465 ( .A(n13232), .B(n13231), .Z(n13234) );
  AND U13466 ( .A(\stack[1][50] ), .B(o[8]), .Z(n13233) );
  XNOR U13467 ( .A(n13234), .B(n13233), .Z(n13237) );
  OR U13468 ( .A(n12886), .B(n12885), .Z(n12890) );
  NANDN U13469 ( .A(n12888), .B(n12887), .Z(n12889) );
  NAND U13470 ( .A(n12890), .B(n12889), .Z(n13238) );
  XNOR U13471 ( .A(n13237), .B(n13238), .Z(n13240) );
  XNOR U13472 ( .A(n13239), .B(n13240), .Z(n13186) );
  OR U13473 ( .A(n12892), .B(n12891), .Z(n12896) );
  OR U13474 ( .A(n12894), .B(n12893), .Z(n12895) );
  AND U13475 ( .A(n12896), .B(n12895), .Z(n13185) );
  XOR U13476 ( .A(n13186), .B(n13185), .Z(n13187) );
  XOR U13477 ( .A(n13188), .B(n13187), .Z(n13180) );
  XNOR U13478 ( .A(n13179), .B(n13180), .Z(n13181) );
  XOR U13479 ( .A(n13174), .B(n13173), .Z(n13176) );
  ANDN U13480 ( .B(o[12]), .A(n15701), .Z(n13175) );
  XOR U13481 ( .A(n13176), .B(n13175), .Z(n13244) );
  ANDN U13482 ( .B(o[13]), .A(n15740), .Z(n13243) );
  XOR U13483 ( .A(n13244), .B(n13243), .Z(n13246) );
  XNOR U13484 ( .A(n13245), .B(n13246), .Z(n13250) );
  NANDN U13485 ( .A(n12898), .B(n12897), .Z(n12902) );
  OR U13486 ( .A(n12900), .B(n12899), .Z(n12901) );
  AND U13487 ( .A(n12902), .B(n12901), .Z(n13249) );
  XNOR U13488 ( .A(n13250), .B(n13249), .Z(n13252) );
  ANDN U13489 ( .B(o[14]), .A(n15779), .Z(n13251) );
  XOR U13490 ( .A(n13252), .B(n13251), .Z(n13168) );
  OR U13491 ( .A(n12904), .B(n12903), .Z(n12908) );
  NANDN U13492 ( .A(n12906), .B(n12905), .Z(n12907) );
  AND U13493 ( .A(n12908), .B(n12907), .Z(n13167) );
  XNOR U13494 ( .A(n13168), .B(n13167), .Z(n13169) );
  XOR U13495 ( .A(n13170), .B(n13169), .Z(n13163) );
  XNOR U13496 ( .A(n13164), .B(n13163), .Z(n13256) );
  ANDN U13497 ( .B(o[17]), .A(n15896), .Z(n13255) );
  XOR U13498 ( .A(n13256), .B(n13255), .Z(n13257) );
  NANDN U13499 ( .A(n12910), .B(n12909), .Z(n12914) );
  OR U13500 ( .A(n12912), .B(n12911), .Z(n12913) );
  AND U13501 ( .A(n12914), .B(n12913), .Z(n13155) );
  XNOR U13502 ( .A(n13156), .B(n13155), .Z(n13158) );
  NANDN U13503 ( .A(n3012), .B(\stack[1][40] ), .Z(n13157) );
  XOR U13504 ( .A(n13158), .B(n13157), .Z(n13261) );
  XOR U13505 ( .A(n13262), .B(n13261), .Z(n13264) );
  OR U13506 ( .A(n12916), .B(n12915), .Z(n12920) );
  NANDN U13507 ( .A(n12918), .B(n12917), .Z(n12919) );
  AND U13508 ( .A(n12920), .B(n12919), .Z(n13263) );
  XOR U13509 ( .A(n13264), .B(n13263), .Z(n13150) );
  XNOR U13510 ( .A(n13149), .B(n13150), .Z(n13152) );
  XNOR U13511 ( .A(n13151), .B(n13152), .Z(n13145) );
  XNOR U13512 ( .A(n13146), .B(n13145), .Z(n13267) );
  XNOR U13513 ( .A(n13268), .B(n13267), .Z(n13270) );
  AND U13514 ( .A(\stack[1][36] ), .B(o[22]), .Z(n13269) );
  XNOR U13515 ( .A(n13270), .B(n13269), .Z(n13139) );
  AND U13516 ( .A(\stack[1][35] ), .B(o[23]), .Z(n13137) );
  OR U13517 ( .A(n12922), .B(n12921), .Z(n12926) );
  OR U13518 ( .A(n12924), .B(n12923), .Z(n12925) );
  NAND U13519 ( .A(n12926), .B(n12925), .Z(n13138) );
  XNOR U13520 ( .A(n13137), .B(n13138), .Z(n13140) );
  XNOR U13521 ( .A(n13139), .B(n13140), .Z(n13132) );
  XOR U13522 ( .A(n13131), .B(n13132), .Z(n13133) );
  AND U13523 ( .A(\stack[1][34] ), .B(o[24]), .Z(n13134) );
  XOR U13524 ( .A(n13133), .B(n13134), .Z(n13127) );
  XOR U13525 ( .A(n13128), .B(n13127), .Z(n13274) );
  XNOR U13526 ( .A(n13273), .B(n13274), .Z(n13275) );
  XOR U13527 ( .A(n13121), .B(n13122), .Z(n13113) );
  OR U13528 ( .A(n12928), .B(n12927), .Z(n12932) );
  NANDN U13529 ( .A(n12930), .B(n12929), .Z(n12931) );
  AND U13530 ( .A(n12932), .B(n12931), .Z(n13114) );
  XOR U13531 ( .A(n13113), .B(n13114), .Z(n13116) );
  AND U13532 ( .A(\stack[1][30] ), .B(o[28]), .Z(n13115) );
  XOR U13533 ( .A(n13116), .B(n13115), .Z(n13281) );
  XOR U13534 ( .A(n13282), .B(n13281), .Z(n13108) );
  XOR U13535 ( .A(n13107), .B(n13108), .Z(n13109) );
  XOR U13536 ( .A(n13110), .B(n13109), .Z(n13104) );
  AND U13537 ( .A(o[31]), .B(\stack[1][27] ), .Z(n13101) );
  OR U13538 ( .A(n12934), .B(n12933), .Z(n12938) );
  OR U13539 ( .A(n12936), .B(n12935), .Z(n12937) );
  NAND U13540 ( .A(n12938), .B(n12937), .Z(n13102) );
  XNOR U13541 ( .A(n13101), .B(n13102), .Z(n13103) );
  XOR U13542 ( .A(n13104), .B(n13103), .Z(n13285) );
  XNOR U13543 ( .A(n13286), .B(n13285), .Z(n13287) );
  XNOR U13544 ( .A(n13288), .B(n13287), .Z(n13097) );
  NANDN U13545 ( .A(n2982), .B(o[33]), .Z(n13095) );
  OR U13546 ( .A(n12940), .B(n12939), .Z(n12944) );
  OR U13547 ( .A(n12942), .B(n12941), .Z(n12943) );
  NAND U13548 ( .A(n12944), .B(n12943), .Z(n13096) );
  XOR U13549 ( .A(n13095), .B(n13096), .Z(n13098) );
  XNOR U13550 ( .A(n13097), .B(n13098), .Z(n13291) );
  XNOR U13551 ( .A(n13292), .B(n13291), .Z(n13293) );
  XNOR U13552 ( .A(n13294), .B(n13293), .Z(n13091) );
  NANDN U13553 ( .A(n2980), .B(o[35]), .Z(n13089) );
  OR U13554 ( .A(n12946), .B(n12945), .Z(n12950) );
  OR U13555 ( .A(n12948), .B(n12947), .Z(n12949) );
  NAND U13556 ( .A(n12950), .B(n12949), .Z(n13090) );
  XOR U13557 ( .A(n13089), .B(n13090), .Z(n13092) );
  XNOR U13558 ( .A(n13091), .B(n13092), .Z(n13297) );
  XNOR U13559 ( .A(n13298), .B(n13297), .Z(n13299) );
  XNOR U13560 ( .A(n13300), .B(n13299), .Z(n13085) );
  NANDN U13561 ( .A(n2978), .B(o[37]), .Z(n13083) );
  OR U13562 ( .A(n12952), .B(n12951), .Z(n12956) );
  OR U13563 ( .A(n12954), .B(n12953), .Z(n12955) );
  NAND U13564 ( .A(n12956), .B(n12955), .Z(n13084) );
  XOR U13565 ( .A(n13083), .B(n13084), .Z(n13086) );
  XNOR U13566 ( .A(n13085), .B(n13086), .Z(n13303) );
  XNOR U13567 ( .A(n13304), .B(n13303), .Z(n13305) );
  XNOR U13568 ( .A(n13306), .B(n13305), .Z(n13079) );
  NANDN U13569 ( .A(n16746), .B(o[39]), .Z(n13077) );
  OR U13570 ( .A(n12958), .B(n12957), .Z(n12962) );
  OR U13571 ( .A(n12960), .B(n12959), .Z(n12961) );
  NAND U13572 ( .A(n12962), .B(n12961), .Z(n13078) );
  XOR U13573 ( .A(n13077), .B(n13078), .Z(n13080) );
  XNOR U13574 ( .A(n13079), .B(n13080), .Z(n13309) );
  XNOR U13575 ( .A(n13310), .B(n13309), .Z(n13311) );
  XNOR U13576 ( .A(n13312), .B(n13311), .Z(n13073) );
  NANDN U13577 ( .A(n16826), .B(o[41]), .Z(n13071) );
  OR U13578 ( .A(n12964), .B(n12963), .Z(n12968) );
  OR U13579 ( .A(n12966), .B(n12965), .Z(n12967) );
  NAND U13580 ( .A(n12968), .B(n12967), .Z(n13072) );
  XOR U13581 ( .A(n13071), .B(n13072), .Z(n13074) );
  XNOR U13582 ( .A(n13073), .B(n13074), .Z(n13315) );
  XNOR U13583 ( .A(n13316), .B(n13315), .Z(n13317) );
  XNOR U13584 ( .A(n13318), .B(n13317), .Z(n13067) );
  NANDN U13585 ( .A(n2976), .B(o[43]), .Z(n13065) );
  OR U13586 ( .A(n12970), .B(n12969), .Z(n12974) );
  OR U13587 ( .A(n12972), .B(n12971), .Z(n12973) );
  NAND U13588 ( .A(n12974), .B(n12973), .Z(n13066) );
  XOR U13589 ( .A(n13065), .B(n13066), .Z(n13068) );
  XNOR U13590 ( .A(n13067), .B(n13068), .Z(n13321) );
  XNOR U13591 ( .A(n13322), .B(n13321), .Z(n13323) );
  XNOR U13592 ( .A(n13324), .B(n13323), .Z(n13061) );
  NANDN U13593 ( .A(n2974), .B(o[45]), .Z(n13059) );
  OR U13594 ( .A(n12976), .B(n12975), .Z(n12980) );
  OR U13595 ( .A(n12978), .B(n12977), .Z(n12979) );
  NAND U13596 ( .A(n12980), .B(n12979), .Z(n13060) );
  XOR U13597 ( .A(n13059), .B(n13060), .Z(n13062) );
  XNOR U13598 ( .A(n13061), .B(n13062), .Z(n13327) );
  XNOR U13599 ( .A(n13328), .B(n13327), .Z(n13329) );
  XNOR U13600 ( .A(n13330), .B(n13329), .Z(n13055) );
  NANDN U13601 ( .A(n2972), .B(o[47]), .Z(n13053) );
  OR U13602 ( .A(n12982), .B(n12981), .Z(n12986) );
  OR U13603 ( .A(n12984), .B(n12983), .Z(n12985) );
  NAND U13604 ( .A(n12986), .B(n12985), .Z(n13054) );
  XOR U13605 ( .A(n13053), .B(n13054), .Z(n13056) );
  XNOR U13606 ( .A(n13055), .B(n13056), .Z(n13333) );
  XNOR U13607 ( .A(n13334), .B(n13333), .Z(n13335) );
  XNOR U13608 ( .A(n13336), .B(n13335), .Z(n13049) );
  NANDN U13609 ( .A(n17145), .B(o[49]), .Z(n13047) );
  OR U13610 ( .A(n12988), .B(n12987), .Z(n12992) );
  OR U13611 ( .A(n12990), .B(n12989), .Z(n12991) );
  NAND U13612 ( .A(n12992), .B(n12991), .Z(n13048) );
  XOR U13613 ( .A(n13047), .B(n13048), .Z(n13050) );
  XNOR U13614 ( .A(n13049), .B(n13050), .Z(n13339) );
  XNOR U13615 ( .A(n13340), .B(n13339), .Z(n13341) );
  XNOR U13616 ( .A(n13342), .B(n13341), .Z(n13043) );
  NANDN U13617 ( .A(n17219), .B(o[51]), .Z(n13041) );
  OR U13618 ( .A(n12994), .B(n12993), .Z(n12998) );
  OR U13619 ( .A(n12996), .B(n12995), .Z(n12997) );
  NAND U13620 ( .A(n12998), .B(n12997), .Z(n13042) );
  XOR U13621 ( .A(n13041), .B(n13042), .Z(n13044) );
  XNOR U13622 ( .A(n13043), .B(n13044), .Z(n13345) );
  XNOR U13623 ( .A(n13346), .B(n13345), .Z(n13347) );
  XNOR U13624 ( .A(n13348), .B(n13347), .Z(n13037) );
  NANDN U13625 ( .A(n17296), .B(o[53]), .Z(n13035) );
  OR U13626 ( .A(n13000), .B(n12999), .Z(n13004) );
  OR U13627 ( .A(n13002), .B(n13001), .Z(n13003) );
  NAND U13628 ( .A(n13004), .B(n13003), .Z(n13036) );
  XOR U13629 ( .A(n13035), .B(n13036), .Z(n13038) );
  XNOR U13630 ( .A(n13037), .B(n13038), .Z(n13351) );
  XNOR U13631 ( .A(n13352), .B(n13351), .Z(n13353) );
  XNOR U13632 ( .A(n13354), .B(n13353), .Z(n13031) );
  NANDN U13633 ( .A(n17375), .B(o[55]), .Z(n13029) );
  OR U13634 ( .A(n13006), .B(n13005), .Z(n13010) );
  OR U13635 ( .A(n13008), .B(n13007), .Z(n13009) );
  NAND U13636 ( .A(n13010), .B(n13009), .Z(n13030) );
  XOR U13637 ( .A(n13029), .B(n13030), .Z(n13032) );
  XNOR U13638 ( .A(n13031), .B(n13032), .Z(n13357) );
  XNOR U13639 ( .A(n13358), .B(n13357), .Z(n13359) );
  AND U13640 ( .A(o[57]), .B(\stack[1][1] ), .Z(n13023) );
  OR U13641 ( .A(n13012), .B(n13011), .Z(n13016) );
  OR U13642 ( .A(n13014), .B(n13013), .Z(n13015) );
  NAND U13643 ( .A(n13016), .B(n13015), .Z(n13024) );
  XNOR U13644 ( .A(n13023), .B(n13024), .Z(n13026) );
  XOR U13645 ( .A(n13025), .B(n13026), .Z(n13017) );
  NANDN U13646 ( .A(n13018), .B(n13017), .Z(n13020) );
  XOR U13647 ( .A(n13018), .B(n13017), .Z(n15241) );
  AND U13648 ( .A(o[58]), .B(\stack[1][0] ), .Z(n15242) );
  OR U13649 ( .A(n15241), .B(n15242), .Z(n13019) );
  AND U13650 ( .A(n13020), .B(n13019), .Z(n13022) );
  OR U13651 ( .A(n13021), .B(n13022), .Z(n13364) );
  XNOR U13652 ( .A(n13022), .B(n13021), .Z(n15202) );
  NANDN U13653 ( .A(n2969), .B(o[58]), .Z(n13708) );
  OR U13654 ( .A(n13024), .B(n13023), .Z(n13028) );
  OR U13655 ( .A(n13026), .B(n13025), .Z(n13027) );
  NAND U13656 ( .A(n13028), .B(n13027), .Z(n13706) );
  NANDN U13657 ( .A(n17375), .B(o[56]), .Z(n13702) );
  NANDN U13658 ( .A(n13030), .B(n13029), .Z(n13034) );
  NANDN U13659 ( .A(n13032), .B(n13031), .Z(n13033) );
  NAND U13660 ( .A(n13034), .B(n13033), .Z(n13700) );
  NANDN U13661 ( .A(n17296), .B(o[54]), .Z(n13696) );
  NANDN U13662 ( .A(n13036), .B(n13035), .Z(n13040) );
  NANDN U13663 ( .A(n13038), .B(n13037), .Z(n13039) );
  NAND U13664 ( .A(n13040), .B(n13039), .Z(n13694) );
  NANDN U13665 ( .A(n17219), .B(o[52]), .Z(n13690) );
  NANDN U13666 ( .A(n13042), .B(n13041), .Z(n13046) );
  NANDN U13667 ( .A(n13044), .B(n13043), .Z(n13045) );
  NAND U13668 ( .A(n13046), .B(n13045), .Z(n13688) );
  NANDN U13669 ( .A(n17145), .B(o[50]), .Z(n13684) );
  NANDN U13670 ( .A(n13048), .B(n13047), .Z(n13052) );
  NANDN U13671 ( .A(n13050), .B(n13049), .Z(n13051) );
  NAND U13672 ( .A(n13052), .B(n13051), .Z(n13682) );
  NANDN U13673 ( .A(n2972), .B(o[48]), .Z(n13678) );
  NANDN U13674 ( .A(n13054), .B(n13053), .Z(n13058) );
  NANDN U13675 ( .A(n13056), .B(n13055), .Z(n13057) );
  NAND U13676 ( .A(n13058), .B(n13057), .Z(n13676) );
  NANDN U13677 ( .A(n2974), .B(o[46]), .Z(n13672) );
  NANDN U13678 ( .A(n13060), .B(n13059), .Z(n13064) );
  NANDN U13679 ( .A(n13062), .B(n13061), .Z(n13063) );
  NAND U13680 ( .A(n13064), .B(n13063), .Z(n13670) );
  NANDN U13681 ( .A(n2976), .B(o[44]), .Z(n13666) );
  NANDN U13682 ( .A(n13066), .B(n13065), .Z(n13070) );
  NANDN U13683 ( .A(n13068), .B(n13067), .Z(n13069) );
  NAND U13684 ( .A(n13070), .B(n13069), .Z(n13664) );
  NANDN U13685 ( .A(n16826), .B(o[42]), .Z(n13660) );
  NANDN U13686 ( .A(n13072), .B(n13071), .Z(n13076) );
  NANDN U13687 ( .A(n13074), .B(n13073), .Z(n13075) );
  NAND U13688 ( .A(n13076), .B(n13075), .Z(n13658) );
  NANDN U13689 ( .A(n16746), .B(o[40]), .Z(n13654) );
  NANDN U13690 ( .A(n13078), .B(n13077), .Z(n13082) );
  NANDN U13691 ( .A(n13080), .B(n13079), .Z(n13081) );
  NAND U13692 ( .A(n13082), .B(n13081), .Z(n13652) );
  NANDN U13693 ( .A(n2978), .B(o[38]), .Z(n13648) );
  NANDN U13694 ( .A(n13084), .B(n13083), .Z(n13088) );
  NANDN U13695 ( .A(n13086), .B(n13085), .Z(n13087) );
  NAND U13696 ( .A(n13088), .B(n13087), .Z(n13646) );
  NANDN U13697 ( .A(n2980), .B(o[36]), .Z(n13642) );
  NANDN U13698 ( .A(n13090), .B(n13089), .Z(n13094) );
  NANDN U13699 ( .A(n13092), .B(n13091), .Z(n13093) );
  NAND U13700 ( .A(n13094), .B(n13093), .Z(n13640) );
  NANDN U13701 ( .A(n2982), .B(o[34]), .Z(n13636) );
  NANDN U13702 ( .A(n13096), .B(n13095), .Z(n13100) );
  NANDN U13703 ( .A(n13098), .B(n13097), .Z(n13099) );
  NAND U13704 ( .A(n13100), .B(n13099), .Z(n13634) );
  AND U13705 ( .A(o[32]), .B(\stack[1][27] ), .Z(n13630) );
  OR U13706 ( .A(n13102), .B(n13101), .Z(n13106) );
  OR U13707 ( .A(n13104), .B(n13103), .Z(n13105) );
  AND U13708 ( .A(n13106), .B(n13105), .Z(n13627) );
  OR U13709 ( .A(n13108), .B(n13107), .Z(n13112) );
  NANDN U13710 ( .A(n13110), .B(n13109), .Z(n13111) );
  AND U13711 ( .A(n13112), .B(n13111), .Z(n13443) );
  AND U13712 ( .A(o[31]), .B(\stack[1][28] ), .Z(n13444) );
  XNOR U13713 ( .A(n13443), .B(n13444), .Z(n13446) );
  NANDN U13714 ( .A(n13114), .B(n13113), .Z(n13118) );
  OR U13715 ( .A(n13116), .B(n13115), .Z(n13117) );
  NAND U13716 ( .A(n13118), .B(n13117), .Z(n13450) );
  ANDN U13717 ( .B(o[29]), .A(n2987), .Z(n13449) );
  XNOR U13718 ( .A(n13450), .B(n13449), .Z(n13451) );
  NANDN U13719 ( .A(n3021), .B(\stack[1][31] ), .Z(n13618) );
  NANDN U13720 ( .A(n13120), .B(n13119), .Z(n13124) );
  NANDN U13721 ( .A(n13122), .B(n13121), .Z(n13123) );
  AND U13722 ( .A(n13124), .B(n13123), .Z(n13615) );
  NANDN U13723 ( .A(n3020), .B(\stack[1][33] ), .Z(n13612) );
  OR U13724 ( .A(n13126), .B(n13125), .Z(n13130) );
  OR U13725 ( .A(n13128), .B(n13127), .Z(n13129) );
  NAND U13726 ( .A(n13130), .B(n13129), .Z(n13610) );
  OR U13727 ( .A(n13132), .B(n13131), .Z(n13136) );
  NANDN U13728 ( .A(n13134), .B(n13133), .Z(n13135) );
  AND U13729 ( .A(n13136), .B(n13135), .Z(n13461) );
  AND U13730 ( .A(\stack[1][34] ), .B(o[25]), .Z(n13462) );
  XNOR U13731 ( .A(n13461), .B(n13462), .Z(n13464) );
  OR U13732 ( .A(n13138), .B(n13137), .Z(n13142) );
  OR U13733 ( .A(n13140), .B(n13139), .Z(n13141) );
  AND U13734 ( .A(n13142), .B(n13141), .Z(n13603) );
  OR U13735 ( .A(n13144), .B(n13143), .Z(n13148) );
  NANDN U13736 ( .A(n13146), .B(n13145), .Z(n13147) );
  NAND U13737 ( .A(n13148), .B(n13147), .Z(n13474) );
  ANDN U13738 ( .B(\stack[1][38] ), .A(n3015), .Z(n13482) );
  OR U13739 ( .A(n13150), .B(n13149), .Z(n13154) );
  NANDN U13740 ( .A(n13152), .B(n13151), .Z(n13153) );
  AND U13741 ( .A(n13154), .B(n13153), .Z(n13479) );
  NANDN U13742 ( .A(n3013), .B(\stack[1][40] ), .Z(n13600) );
  OR U13743 ( .A(n13156), .B(n13155), .Z(n13160) );
  OR U13744 ( .A(n13158), .B(n13157), .Z(n13159) );
  AND U13745 ( .A(n13160), .B(n13159), .Z(n13598) );
  OR U13746 ( .A(n13162), .B(n13161), .Z(n13166) );
  NAND U13747 ( .A(n13164), .B(n13163), .Z(n13165) );
  AND U13748 ( .A(n13166), .B(n13165), .Z(n13588) );
  OR U13749 ( .A(n13168), .B(n13167), .Z(n13172) );
  OR U13750 ( .A(n13170), .B(n13169), .Z(n13171) );
  AND U13751 ( .A(n13172), .B(n13171), .Z(n13491) );
  NANDN U13752 ( .A(n3010), .B(\stack[1][43] ), .Z(n13492) );
  XOR U13753 ( .A(n13491), .B(n13492), .Z(n13494) );
  NANDN U13754 ( .A(n3009), .B(\stack[1][44] ), .Z(n13500) );
  NANDN U13755 ( .A(n13174), .B(n13173), .Z(n13178) );
  NANDN U13756 ( .A(n13176), .B(n13175), .Z(n13177) );
  AND U13757 ( .A(n13178), .B(n13177), .Z(n13576) );
  NANDN U13758 ( .A(n3006), .B(\stack[1][47] ), .Z(n13506) );
  OR U13759 ( .A(n13180), .B(n13179), .Z(n13184) );
  OR U13760 ( .A(n13182), .B(n13181), .Z(n13183) );
  NAND U13761 ( .A(n13184), .B(n13183), .Z(n13504) );
  NANDN U13762 ( .A(n15623), .B(o[11]), .Z(n13511) );
  OR U13763 ( .A(n13186), .B(n13185), .Z(n13190) );
  NANDN U13764 ( .A(n13188), .B(n13187), .Z(n13189) );
  AND U13765 ( .A(n13190), .B(n13189), .Z(n13510) );
  NANDN U13766 ( .A(n3004), .B(\stack[1][49] ), .Z(n13517) );
  AND U13767 ( .A(\stack[1][50] ), .B(o[9]), .Z(n13569) );
  NANDN U13768 ( .A(n13192), .B(n13191), .Z(n13196) );
  NAND U13769 ( .A(n13194), .B(n13193), .Z(n13195) );
  AND U13770 ( .A(n13196), .B(n13195), .Z(n13558) );
  ANDN U13771 ( .B(\stack[1][54] ), .A(n2999), .Z(n13552) );
  OR U13772 ( .A(n13198), .B(n13197), .Z(n13202) );
  NANDN U13773 ( .A(n13200), .B(n13199), .Z(n13201) );
  AND U13774 ( .A(n13202), .B(n13201), .Z(n13549) );
  ANDN U13775 ( .B(\stack[1][55] ), .A(n2998), .Z(n13530) );
  AND U13776 ( .A(\stack[1][56] ), .B(o[3]), .Z(n13546) );
  NANDN U13777 ( .A(n13203), .B(n13533), .Z(n13204) );
  AND U13778 ( .A(n13205), .B(n13204), .Z(n13209) );
  OR U13779 ( .A(n13207), .B(n13206), .Z(n13208) );
  AND U13780 ( .A(n13209), .B(n13208), .Z(n13543) );
  AND U13781 ( .A(\stack[1][59] ), .B(o[1]), .Z(n13541) );
  ANDN U13782 ( .B(n13541), .A(n13210), .Z(n13885) );
  XNOR U13783 ( .A(n13885), .B(n13533), .Z(n13212) );
  NAND U13784 ( .A(\stack[1][59] ), .B(o[0]), .Z(n13540) );
  NANDN U13785 ( .A(n13211), .B(n13540), .Z(n13535) );
  NAND U13786 ( .A(n13212), .B(n13535), .Z(n13537) );
  ANDN U13787 ( .B(\stack[1][57] ), .A(n2996), .Z(n13536) );
  XNOR U13788 ( .A(n13537), .B(n13536), .Z(n13544) );
  XOR U13789 ( .A(n13543), .B(n13544), .Z(n13545) );
  XOR U13790 ( .A(n13546), .B(n13545), .Z(n13528) );
  OR U13791 ( .A(n13214), .B(n13213), .Z(n13218) );
  NANDN U13792 ( .A(n13216), .B(n13215), .Z(n13217) );
  AND U13793 ( .A(n13218), .B(n13217), .Z(n13527) );
  XOR U13794 ( .A(n13528), .B(n13527), .Z(n13529) );
  XOR U13795 ( .A(n13530), .B(n13529), .Z(n13550) );
  XNOR U13796 ( .A(n13549), .B(n13550), .Z(n13551) );
  OR U13797 ( .A(n13220), .B(n13219), .Z(n13224) );
  OR U13798 ( .A(n13222), .B(n13221), .Z(n13223) );
  NAND U13799 ( .A(n13224), .B(n13223), .Z(n13522) );
  ANDN U13800 ( .B(\stack[1][53] ), .A(n3000), .Z(n13521) );
  XNOR U13801 ( .A(n13522), .B(n13521), .Z(n13524) );
  XNOR U13802 ( .A(n13523), .B(n13524), .Z(n13556) );
  ANDN U13803 ( .B(o[7]), .A(n15468), .Z(n13555) );
  XOR U13804 ( .A(n13556), .B(n13555), .Z(n13557) );
  NANDN U13805 ( .A(n13226), .B(n13225), .Z(n13230) );
  OR U13806 ( .A(n13228), .B(n13227), .Z(n13229) );
  AND U13807 ( .A(n13230), .B(n13229), .Z(n13561) );
  XNOR U13808 ( .A(n13562), .B(n13561), .Z(n13564) );
  AND U13809 ( .A(\stack[1][51] ), .B(o[8]), .Z(n13563) );
  XNOR U13810 ( .A(n13564), .B(n13563), .Z(n13567) );
  OR U13811 ( .A(n13232), .B(n13231), .Z(n13236) );
  NANDN U13812 ( .A(n13234), .B(n13233), .Z(n13235) );
  NAND U13813 ( .A(n13236), .B(n13235), .Z(n13568) );
  XNOR U13814 ( .A(n13567), .B(n13568), .Z(n13570) );
  XNOR U13815 ( .A(n13569), .B(n13570), .Z(n13516) );
  OR U13816 ( .A(n13238), .B(n13237), .Z(n13242) );
  OR U13817 ( .A(n13240), .B(n13239), .Z(n13241) );
  AND U13818 ( .A(n13242), .B(n13241), .Z(n13515) );
  XNOR U13819 ( .A(n13516), .B(n13515), .Z(n13518) );
  XNOR U13820 ( .A(n13517), .B(n13518), .Z(n13509) );
  XOR U13821 ( .A(n13510), .B(n13509), .Z(n13512) );
  XNOR U13822 ( .A(n13511), .B(n13512), .Z(n13503) );
  XNOR U13823 ( .A(n13504), .B(n13503), .Z(n13505) );
  XNOR U13824 ( .A(n13506), .B(n13505), .Z(n13574) );
  ANDN U13825 ( .B(o[13]), .A(n15701), .Z(n13573) );
  XOR U13826 ( .A(n13574), .B(n13573), .Z(n13575) );
  NANDN U13827 ( .A(n13244), .B(n13243), .Z(n13248) );
  OR U13828 ( .A(n13246), .B(n13245), .Z(n13247) );
  AND U13829 ( .A(n13248), .B(n13247), .Z(n13579) );
  XNOR U13830 ( .A(n13580), .B(n13579), .Z(n13582) );
  ANDN U13831 ( .B(o[14]), .A(n15740), .Z(n13581) );
  XOR U13832 ( .A(n13582), .B(n13581), .Z(n13498) );
  OR U13833 ( .A(n13250), .B(n13249), .Z(n13254) );
  NANDN U13834 ( .A(n13252), .B(n13251), .Z(n13253) );
  AND U13835 ( .A(n13254), .B(n13253), .Z(n13497) );
  XNOR U13836 ( .A(n13498), .B(n13497), .Z(n13499) );
  XOR U13837 ( .A(n13500), .B(n13499), .Z(n13493) );
  XNOR U13838 ( .A(n13494), .B(n13493), .Z(n13586) );
  ANDN U13839 ( .B(o[17]), .A(n15857), .Z(n13585) );
  XOR U13840 ( .A(n13586), .B(n13585), .Z(n13587) );
  NANDN U13841 ( .A(n13256), .B(n13255), .Z(n13260) );
  OR U13842 ( .A(n13258), .B(n13257), .Z(n13259) );
  AND U13843 ( .A(n13260), .B(n13259), .Z(n13591) );
  XNOR U13844 ( .A(n13592), .B(n13591), .Z(n13594) );
  NANDN U13845 ( .A(n3012), .B(\stack[1][41] ), .Z(n13593) );
  XOR U13846 ( .A(n13594), .B(n13593), .Z(n13597) );
  XOR U13847 ( .A(n13598), .B(n13597), .Z(n13599) );
  XNOR U13848 ( .A(n13600), .B(n13599), .Z(n13485) );
  NANDN U13849 ( .A(n13262), .B(n13261), .Z(n13266) );
  OR U13850 ( .A(n13264), .B(n13263), .Z(n13265) );
  NAND U13851 ( .A(n13266), .B(n13265), .Z(n13486) );
  XOR U13852 ( .A(n13485), .B(n13486), .Z(n13488) );
  AND U13853 ( .A(\stack[1][39] ), .B(o[20]), .Z(n13487) );
  XNOR U13854 ( .A(n13488), .B(n13487), .Z(n13480) );
  XNOR U13855 ( .A(n13479), .B(n13480), .Z(n13481) );
  XOR U13856 ( .A(n13474), .B(n13473), .Z(n13476) );
  AND U13857 ( .A(\stack[1][37] ), .B(o[22]), .Z(n13475) );
  XNOR U13858 ( .A(n13476), .B(n13475), .Z(n13469) );
  AND U13859 ( .A(\stack[1][36] ), .B(o[23]), .Z(n13467) );
  OR U13860 ( .A(n13268), .B(n13267), .Z(n13272) );
  NANDN U13861 ( .A(n13270), .B(n13269), .Z(n13271) );
  NAND U13862 ( .A(n13272), .B(n13271), .Z(n13468) );
  XNOR U13863 ( .A(n13467), .B(n13468), .Z(n13470) );
  XNOR U13864 ( .A(n13469), .B(n13470), .Z(n13604) );
  XOR U13865 ( .A(n13603), .B(n13604), .Z(n13605) );
  AND U13866 ( .A(\stack[1][35] ), .B(o[24]), .Z(n13606) );
  XOR U13867 ( .A(n13605), .B(n13606), .Z(n13463) );
  XOR U13868 ( .A(n13464), .B(n13463), .Z(n13609) );
  XNOR U13869 ( .A(n13610), .B(n13609), .Z(n13611) );
  XNOR U13870 ( .A(n13612), .B(n13611), .Z(n13457) );
  NANDN U13871 ( .A(n2989), .B(o[27]), .Z(n13455) );
  OR U13872 ( .A(n13274), .B(n13273), .Z(n13278) );
  OR U13873 ( .A(n13276), .B(n13275), .Z(n13277) );
  NAND U13874 ( .A(n13278), .B(n13277), .Z(n13456) );
  XOR U13875 ( .A(n13455), .B(n13456), .Z(n13458) );
  XNOR U13876 ( .A(n13457), .B(n13458), .Z(n13616) );
  XNOR U13877 ( .A(n13615), .B(n13616), .Z(n13617) );
  XOR U13878 ( .A(n13451), .B(n13452), .Z(n13621) );
  OR U13879 ( .A(n13280), .B(n13279), .Z(n13284) );
  NANDN U13880 ( .A(n13282), .B(n13281), .Z(n13283) );
  AND U13881 ( .A(n13284), .B(n13283), .Z(n13622) );
  XOR U13882 ( .A(n13621), .B(n13622), .Z(n13624) );
  AND U13883 ( .A(o[30]), .B(\stack[1][29] ), .Z(n13623) );
  XOR U13884 ( .A(n13624), .B(n13623), .Z(n13445) );
  XOR U13885 ( .A(n13446), .B(n13445), .Z(n13628) );
  XOR U13886 ( .A(n13627), .B(n13628), .Z(n13629) );
  XOR U13887 ( .A(n13630), .B(n13629), .Z(n13440) );
  AND U13888 ( .A(o[33]), .B(\stack[1][26] ), .Z(n13437) );
  OR U13889 ( .A(n13286), .B(n13285), .Z(n13290) );
  OR U13890 ( .A(n13288), .B(n13287), .Z(n13289) );
  NAND U13891 ( .A(n13290), .B(n13289), .Z(n13438) );
  XNOR U13892 ( .A(n13437), .B(n13438), .Z(n13439) );
  XOR U13893 ( .A(n13440), .B(n13439), .Z(n13633) );
  XNOR U13894 ( .A(n13634), .B(n13633), .Z(n13635) );
  XNOR U13895 ( .A(n13636), .B(n13635), .Z(n13433) );
  NANDN U13896 ( .A(n2981), .B(o[35]), .Z(n13431) );
  OR U13897 ( .A(n13292), .B(n13291), .Z(n13296) );
  OR U13898 ( .A(n13294), .B(n13293), .Z(n13295) );
  NAND U13899 ( .A(n13296), .B(n13295), .Z(n13432) );
  XOR U13900 ( .A(n13431), .B(n13432), .Z(n13434) );
  XNOR U13901 ( .A(n13433), .B(n13434), .Z(n13639) );
  XNOR U13902 ( .A(n13640), .B(n13639), .Z(n13641) );
  XNOR U13903 ( .A(n13642), .B(n13641), .Z(n13427) );
  NANDN U13904 ( .A(n2979), .B(o[37]), .Z(n13425) );
  OR U13905 ( .A(n13298), .B(n13297), .Z(n13302) );
  OR U13906 ( .A(n13300), .B(n13299), .Z(n13301) );
  NAND U13907 ( .A(n13302), .B(n13301), .Z(n13426) );
  XOR U13908 ( .A(n13425), .B(n13426), .Z(n13428) );
  XNOR U13909 ( .A(n13427), .B(n13428), .Z(n13645) );
  XNOR U13910 ( .A(n13646), .B(n13645), .Z(n13647) );
  XNOR U13911 ( .A(n13648), .B(n13647), .Z(n13421) );
  NANDN U13912 ( .A(n16712), .B(o[39]), .Z(n13419) );
  OR U13913 ( .A(n13304), .B(n13303), .Z(n13308) );
  OR U13914 ( .A(n13306), .B(n13305), .Z(n13307) );
  NAND U13915 ( .A(n13308), .B(n13307), .Z(n13420) );
  XOR U13916 ( .A(n13419), .B(n13420), .Z(n13422) );
  XNOR U13917 ( .A(n13421), .B(n13422), .Z(n13651) );
  XNOR U13918 ( .A(n13652), .B(n13651), .Z(n13653) );
  XNOR U13919 ( .A(n13654), .B(n13653), .Z(n13415) );
  NANDN U13920 ( .A(n16786), .B(o[41]), .Z(n13413) );
  OR U13921 ( .A(n13310), .B(n13309), .Z(n13314) );
  OR U13922 ( .A(n13312), .B(n13311), .Z(n13313) );
  NAND U13923 ( .A(n13314), .B(n13313), .Z(n13414) );
  XOR U13924 ( .A(n13413), .B(n13414), .Z(n13416) );
  XNOR U13925 ( .A(n13415), .B(n13416), .Z(n13657) );
  XNOR U13926 ( .A(n13658), .B(n13657), .Z(n13659) );
  XNOR U13927 ( .A(n13660), .B(n13659), .Z(n13409) );
  NANDN U13928 ( .A(n2977), .B(o[43]), .Z(n13407) );
  OR U13929 ( .A(n13316), .B(n13315), .Z(n13320) );
  OR U13930 ( .A(n13318), .B(n13317), .Z(n13319) );
  NAND U13931 ( .A(n13320), .B(n13319), .Z(n13408) );
  XOR U13932 ( .A(n13407), .B(n13408), .Z(n13410) );
  XNOR U13933 ( .A(n13409), .B(n13410), .Z(n13663) );
  XNOR U13934 ( .A(n13664), .B(n13663), .Z(n13665) );
  XNOR U13935 ( .A(n13666), .B(n13665), .Z(n13403) );
  NANDN U13936 ( .A(n2975), .B(o[45]), .Z(n13401) );
  OR U13937 ( .A(n13322), .B(n13321), .Z(n13326) );
  OR U13938 ( .A(n13324), .B(n13323), .Z(n13325) );
  NAND U13939 ( .A(n13326), .B(n13325), .Z(n13402) );
  XOR U13940 ( .A(n13401), .B(n13402), .Z(n13404) );
  XNOR U13941 ( .A(n13403), .B(n13404), .Z(n13669) );
  XNOR U13942 ( .A(n13670), .B(n13669), .Z(n13671) );
  XNOR U13943 ( .A(n13672), .B(n13671), .Z(n13397) );
  NANDN U13944 ( .A(n2973), .B(o[47]), .Z(n13395) );
  OR U13945 ( .A(n13328), .B(n13327), .Z(n13332) );
  OR U13946 ( .A(n13330), .B(n13329), .Z(n13331) );
  NAND U13947 ( .A(n13332), .B(n13331), .Z(n13396) );
  XOR U13948 ( .A(n13395), .B(n13396), .Z(n13398) );
  XNOR U13949 ( .A(n13397), .B(n13398), .Z(n13675) );
  XNOR U13950 ( .A(n13676), .B(n13675), .Z(n13677) );
  XNOR U13951 ( .A(n13678), .B(n13677), .Z(n13391) );
  NANDN U13952 ( .A(n17101), .B(o[49]), .Z(n13389) );
  OR U13953 ( .A(n13334), .B(n13333), .Z(n13338) );
  OR U13954 ( .A(n13336), .B(n13335), .Z(n13337) );
  NAND U13955 ( .A(n13338), .B(n13337), .Z(n13390) );
  XOR U13956 ( .A(n13389), .B(n13390), .Z(n13392) );
  XNOR U13957 ( .A(n13391), .B(n13392), .Z(n13681) );
  XNOR U13958 ( .A(n13682), .B(n13681), .Z(n13683) );
  XNOR U13959 ( .A(n13684), .B(n13683), .Z(n13385) );
  NANDN U13960 ( .A(n17179), .B(o[51]), .Z(n13383) );
  OR U13961 ( .A(n13340), .B(n13339), .Z(n13344) );
  OR U13962 ( .A(n13342), .B(n13341), .Z(n13343) );
  NAND U13963 ( .A(n13344), .B(n13343), .Z(n13384) );
  XOR U13964 ( .A(n13383), .B(n13384), .Z(n13386) );
  XNOR U13965 ( .A(n13385), .B(n13386), .Z(n13687) );
  XNOR U13966 ( .A(n13688), .B(n13687), .Z(n13689) );
  XNOR U13967 ( .A(n13690), .B(n13689), .Z(n13379) );
  NANDN U13968 ( .A(n17256), .B(o[53]), .Z(n13377) );
  OR U13969 ( .A(n13346), .B(n13345), .Z(n13350) );
  OR U13970 ( .A(n13348), .B(n13347), .Z(n13349) );
  NAND U13971 ( .A(n13350), .B(n13349), .Z(n13378) );
  XOR U13972 ( .A(n13377), .B(n13378), .Z(n13380) );
  XNOR U13973 ( .A(n13379), .B(n13380), .Z(n13693) );
  XNOR U13974 ( .A(n13694), .B(n13693), .Z(n13695) );
  XNOR U13975 ( .A(n13696), .B(n13695), .Z(n13373) );
  AND U13976 ( .A(o[55]), .B(\stack[1][4] ), .Z(n13371) );
  OR U13977 ( .A(n13352), .B(n13351), .Z(n13356) );
  OR U13978 ( .A(n13354), .B(n13353), .Z(n13355) );
  NAND U13979 ( .A(n13356), .B(n13355), .Z(n13372) );
  XNOR U13980 ( .A(n13371), .B(n13372), .Z(n13374) );
  XNOR U13981 ( .A(n13373), .B(n13374), .Z(n13699) );
  XNOR U13982 ( .A(n13700), .B(n13699), .Z(n13701) );
  XOR U13983 ( .A(n13702), .B(n13701), .Z(n13368) );
  AND U13984 ( .A(o[57]), .B(\stack[1][2] ), .Z(n13365) );
  OR U13985 ( .A(n13358), .B(n13357), .Z(n13362) );
  OR U13986 ( .A(n13360), .B(n13359), .Z(n13361) );
  NAND U13987 ( .A(n13362), .B(n13361), .Z(n13366) );
  XOR U13988 ( .A(n13365), .B(n13366), .Z(n13367) );
  XNOR U13989 ( .A(n13368), .B(n13367), .Z(n13705) );
  XNOR U13990 ( .A(n13706), .B(n13705), .Z(n13707) );
  XOR U13991 ( .A(n13708), .B(n13707), .Z(n15203) );
  OR U13992 ( .A(n15202), .B(n15203), .Z(n13363) );
  AND U13993 ( .A(n13364), .B(n13363), .Z(n13712) );
  NANDN U13994 ( .A(n2970), .B(o[58]), .Z(n14066) );
  OR U13995 ( .A(n13366), .B(n13365), .Z(n13370) );
  NANDN U13996 ( .A(n13368), .B(n13367), .Z(n13369) );
  NAND U13997 ( .A(n13370), .B(n13369), .Z(n14064) );
  NANDN U13998 ( .A(n2971), .B(o[56]), .Z(n14060) );
  OR U13999 ( .A(n13372), .B(n13371), .Z(n13376) );
  NANDN U14000 ( .A(n13374), .B(n13373), .Z(n13375) );
  NAND U14001 ( .A(n13376), .B(n13375), .Z(n14058) );
  NANDN U14002 ( .A(n17256), .B(o[54]), .Z(n14054) );
  NANDN U14003 ( .A(n13378), .B(n13377), .Z(n13382) );
  NANDN U14004 ( .A(n13380), .B(n13379), .Z(n13381) );
  NAND U14005 ( .A(n13382), .B(n13381), .Z(n14052) );
  NANDN U14006 ( .A(n17179), .B(o[52]), .Z(n14048) );
  NANDN U14007 ( .A(n13384), .B(n13383), .Z(n13388) );
  NANDN U14008 ( .A(n13386), .B(n13385), .Z(n13387) );
  NAND U14009 ( .A(n13388), .B(n13387), .Z(n14046) );
  NANDN U14010 ( .A(n17101), .B(o[50]), .Z(n14042) );
  NANDN U14011 ( .A(n13390), .B(n13389), .Z(n13394) );
  NANDN U14012 ( .A(n13392), .B(n13391), .Z(n13393) );
  NAND U14013 ( .A(n13394), .B(n13393), .Z(n14040) );
  NANDN U14014 ( .A(n2973), .B(o[48]), .Z(n14036) );
  NANDN U14015 ( .A(n13396), .B(n13395), .Z(n13400) );
  NANDN U14016 ( .A(n13398), .B(n13397), .Z(n13399) );
  NAND U14017 ( .A(n13400), .B(n13399), .Z(n14034) );
  NANDN U14018 ( .A(n2975), .B(o[46]), .Z(n14030) );
  NANDN U14019 ( .A(n13402), .B(n13401), .Z(n13406) );
  NANDN U14020 ( .A(n13404), .B(n13403), .Z(n13405) );
  NAND U14021 ( .A(n13406), .B(n13405), .Z(n14028) );
  NANDN U14022 ( .A(n2977), .B(o[44]), .Z(n14024) );
  NANDN U14023 ( .A(n13408), .B(n13407), .Z(n13412) );
  NANDN U14024 ( .A(n13410), .B(n13409), .Z(n13411) );
  NAND U14025 ( .A(n13412), .B(n13411), .Z(n14022) );
  NANDN U14026 ( .A(n16786), .B(o[42]), .Z(n14018) );
  NANDN U14027 ( .A(n13414), .B(n13413), .Z(n13418) );
  NANDN U14028 ( .A(n13416), .B(n13415), .Z(n13417) );
  NAND U14029 ( .A(n13418), .B(n13417), .Z(n14016) );
  NANDN U14030 ( .A(n16712), .B(o[40]), .Z(n14012) );
  NANDN U14031 ( .A(n13420), .B(n13419), .Z(n13424) );
  NANDN U14032 ( .A(n13422), .B(n13421), .Z(n13423) );
  NAND U14033 ( .A(n13424), .B(n13423), .Z(n14010) );
  NANDN U14034 ( .A(n2979), .B(o[38]), .Z(n14006) );
  NANDN U14035 ( .A(n13426), .B(n13425), .Z(n13430) );
  NANDN U14036 ( .A(n13428), .B(n13427), .Z(n13429) );
  NAND U14037 ( .A(n13430), .B(n13429), .Z(n14004) );
  NANDN U14038 ( .A(n2981), .B(o[36]), .Z(n14000) );
  NANDN U14039 ( .A(n13432), .B(n13431), .Z(n13436) );
  NANDN U14040 ( .A(n13434), .B(n13433), .Z(n13435) );
  NAND U14041 ( .A(n13436), .B(n13435), .Z(n13998) );
  NANDN U14042 ( .A(n2983), .B(o[34]), .Z(n13994) );
  OR U14043 ( .A(n13438), .B(n13437), .Z(n13442) );
  OR U14044 ( .A(n13440), .B(n13439), .Z(n13441) );
  NAND U14045 ( .A(n13442), .B(n13441), .Z(n13992) );
  NANDN U14046 ( .A(n2985), .B(o[32]), .Z(n13988) );
  OR U14047 ( .A(n13444), .B(n13443), .Z(n13448) );
  NANDN U14048 ( .A(n13446), .B(n13445), .Z(n13447) );
  NAND U14049 ( .A(n13448), .B(n13447), .Z(n13986) );
  ANDN U14050 ( .B(o[30]), .A(n2987), .Z(n13981) );
  NANDN U14051 ( .A(n13450), .B(n13449), .Z(n13454) );
  NANDN U14052 ( .A(n13452), .B(n13451), .Z(n13453) );
  AND U14053 ( .A(n13454), .B(n13453), .Z(n13979) );
  NANDN U14054 ( .A(n3021), .B(\stack[1][32] ), .Z(n13976) );
  NANDN U14055 ( .A(n13456), .B(n13455), .Z(n13460) );
  NANDN U14056 ( .A(n13458), .B(n13457), .Z(n13459) );
  NAND U14057 ( .A(n13460), .B(n13459), .Z(n13974) );
  NANDN U14058 ( .A(n3020), .B(\stack[1][34] ), .Z(n13822) );
  OR U14059 ( .A(n13462), .B(n13461), .Z(n13466) );
  OR U14060 ( .A(n13464), .B(n13463), .Z(n13465) );
  NAND U14061 ( .A(n13466), .B(n13465), .Z(n13820) );
  AND U14062 ( .A(\stack[1][36] ), .B(o[24]), .Z(n13828) );
  OR U14063 ( .A(n13468), .B(n13467), .Z(n13472) );
  OR U14064 ( .A(n13470), .B(n13469), .Z(n13471) );
  AND U14065 ( .A(n13472), .B(n13471), .Z(n13825) );
  AND U14066 ( .A(\stack[1][37] ), .B(o[23]), .Z(n13831) );
  NANDN U14067 ( .A(n13474), .B(n13473), .Z(n13478) );
  NANDN U14068 ( .A(n13476), .B(n13475), .Z(n13477) );
  NAND U14069 ( .A(n13478), .B(n13477), .Z(n13832) );
  XNOR U14070 ( .A(n13831), .B(n13832), .Z(n13834) );
  NANDN U14071 ( .A(n3016), .B(\stack[1][38] ), .Z(n13839) );
  OR U14072 ( .A(n13480), .B(n13479), .Z(n13484) );
  OR U14073 ( .A(n13482), .B(n13481), .Z(n13483) );
  AND U14074 ( .A(n13484), .B(n13483), .Z(n13838) );
  NANDN U14075 ( .A(n3015), .B(\stack[1][39] ), .Z(n13963) );
  NANDN U14076 ( .A(n13486), .B(n13485), .Z(n13490) );
  OR U14077 ( .A(n13488), .B(n13487), .Z(n13489) );
  AND U14078 ( .A(n13490), .B(n13489), .Z(n13962) );
  NANDN U14079 ( .A(n3013), .B(\stack[1][41] ), .Z(n13950) );
  OR U14080 ( .A(n13492), .B(n13491), .Z(n13496) );
  NAND U14081 ( .A(n13494), .B(n13493), .Z(n13495) );
  AND U14082 ( .A(n13496), .B(n13495), .Z(n13940) );
  OR U14083 ( .A(n13498), .B(n13497), .Z(n13502) );
  OR U14084 ( .A(n13500), .B(n13499), .Z(n13501) );
  AND U14085 ( .A(n13502), .B(n13501), .Z(n13843) );
  NANDN U14086 ( .A(n3010), .B(\stack[1][44] ), .Z(n13844) );
  XOR U14087 ( .A(n13843), .B(n13844), .Z(n13846) );
  NANDN U14088 ( .A(n3009), .B(\stack[1][45] ), .Z(n13852) );
  OR U14089 ( .A(n13504), .B(n13503), .Z(n13508) );
  OR U14090 ( .A(n13506), .B(n13505), .Z(n13507) );
  AND U14091 ( .A(n13508), .B(n13507), .Z(n13928) );
  NANDN U14092 ( .A(n13510), .B(n13509), .Z(n13514) );
  NANDN U14093 ( .A(n13512), .B(n13511), .Z(n13513) );
  NAND U14094 ( .A(n13514), .B(n13513), .Z(n13858) );
  NANDN U14095 ( .A(n3006), .B(\stack[1][48] ), .Z(n13856) );
  NANDN U14096 ( .A(n3005), .B(\stack[1][49] ), .Z(n13863) );
  OR U14097 ( .A(n13516), .B(n13515), .Z(n13520) );
  NANDN U14098 ( .A(n13518), .B(n13517), .Z(n13519) );
  AND U14099 ( .A(n13520), .B(n13519), .Z(n13862) );
  NANDN U14100 ( .A(n15546), .B(o[10]), .Z(n13869) );
  AND U14101 ( .A(\stack[1][51] ), .B(o[9]), .Z(n13921) );
  NANDN U14102 ( .A(n13522), .B(n13521), .Z(n13526) );
  NAND U14103 ( .A(n13524), .B(n13523), .Z(n13525) );
  AND U14104 ( .A(n13526), .B(n13525), .Z(n13910) );
  ANDN U14105 ( .B(\stack[1][55] ), .A(n2999), .Z(n13904) );
  OR U14106 ( .A(n13528), .B(n13527), .Z(n13532) );
  NANDN U14107 ( .A(n13530), .B(n13529), .Z(n13531) );
  AND U14108 ( .A(n13532), .B(n13531), .Z(n13901) );
  AND U14109 ( .A(\stack[1][56] ), .B(o[4]), .Z(n13882) );
  ANDN U14110 ( .B(\stack[1][57] ), .A(n2997), .Z(n13898) );
  NANDN U14111 ( .A(n13533), .B(n13885), .Z(n13534) );
  AND U14112 ( .A(n13535), .B(n13534), .Z(n13539) );
  OR U14113 ( .A(n13537), .B(n13536), .Z(n13538) );
  AND U14114 ( .A(n13539), .B(n13538), .Z(n13895) );
  AND U14115 ( .A(\stack[1][60] ), .B(o[1]), .Z(n13893) );
  ANDN U14116 ( .B(n13893), .A(n13540), .Z(n14233) );
  XNOR U14117 ( .A(n14233), .B(n13885), .Z(n13542) );
  NAND U14118 ( .A(\stack[1][60] ), .B(o[0]), .Z(n13892) );
  NANDN U14119 ( .A(n13541), .B(n13892), .Z(n13887) );
  NAND U14120 ( .A(n13542), .B(n13887), .Z(n13889) );
  AND U14121 ( .A(\stack[1][58] ), .B(o[2]), .Z(n13888) );
  XNOR U14122 ( .A(n13889), .B(n13888), .Z(n13896) );
  XOR U14123 ( .A(n13895), .B(n13896), .Z(n13897) );
  XOR U14124 ( .A(n13898), .B(n13897), .Z(n13880) );
  OR U14125 ( .A(n13544), .B(n13543), .Z(n13548) );
  NANDN U14126 ( .A(n13546), .B(n13545), .Z(n13547) );
  AND U14127 ( .A(n13548), .B(n13547), .Z(n13879) );
  XOR U14128 ( .A(n13880), .B(n13879), .Z(n13881) );
  XOR U14129 ( .A(n13882), .B(n13881), .Z(n13902) );
  XNOR U14130 ( .A(n13901), .B(n13902), .Z(n13903) );
  OR U14131 ( .A(n13550), .B(n13549), .Z(n13554) );
  OR U14132 ( .A(n13552), .B(n13551), .Z(n13553) );
  NAND U14133 ( .A(n13554), .B(n13553), .Z(n13874) );
  ANDN U14134 ( .B(\stack[1][54] ), .A(n3000), .Z(n13873) );
  XNOR U14135 ( .A(n13874), .B(n13873), .Z(n13876) );
  XNOR U14136 ( .A(n13875), .B(n13876), .Z(n13908) );
  ANDN U14137 ( .B(\stack[1][53] ), .A(n3001), .Z(n13907) );
  XOR U14138 ( .A(n13908), .B(n13907), .Z(n13909) );
  NANDN U14139 ( .A(n13556), .B(n13555), .Z(n13560) );
  OR U14140 ( .A(n13558), .B(n13557), .Z(n13559) );
  AND U14141 ( .A(n13560), .B(n13559), .Z(n13913) );
  XNOR U14142 ( .A(n13914), .B(n13913), .Z(n13916) );
  AND U14143 ( .A(\stack[1][52] ), .B(o[8]), .Z(n13915) );
  XNOR U14144 ( .A(n13916), .B(n13915), .Z(n13919) );
  OR U14145 ( .A(n13562), .B(n13561), .Z(n13566) );
  NANDN U14146 ( .A(n13564), .B(n13563), .Z(n13565) );
  NAND U14147 ( .A(n13566), .B(n13565), .Z(n13920) );
  XNOR U14148 ( .A(n13919), .B(n13920), .Z(n13922) );
  XNOR U14149 ( .A(n13921), .B(n13922), .Z(n13868) );
  OR U14150 ( .A(n13568), .B(n13567), .Z(n13572) );
  OR U14151 ( .A(n13570), .B(n13569), .Z(n13571) );
  AND U14152 ( .A(n13572), .B(n13571), .Z(n13867) );
  XNOR U14153 ( .A(n13868), .B(n13867), .Z(n13870) );
  XNOR U14154 ( .A(n13869), .B(n13870), .Z(n13861) );
  XOR U14155 ( .A(n13862), .B(n13861), .Z(n13864) );
  XNOR U14156 ( .A(n13863), .B(n13864), .Z(n13855) );
  XNOR U14157 ( .A(n13856), .B(n13855), .Z(n13857) );
  XNOR U14158 ( .A(n13858), .B(n13857), .Z(n13926) );
  ANDN U14159 ( .B(o[13]), .A(n15662), .Z(n13925) );
  XOR U14160 ( .A(n13926), .B(n13925), .Z(n13927) );
  NANDN U14161 ( .A(n13574), .B(n13573), .Z(n13578) );
  OR U14162 ( .A(n13576), .B(n13575), .Z(n13577) );
  AND U14163 ( .A(n13578), .B(n13577), .Z(n13931) );
  XNOR U14164 ( .A(n13932), .B(n13931), .Z(n13934) );
  ANDN U14165 ( .B(o[14]), .A(n15701), .Z(n13933) );
  XOR U14166 ( .A(n13934), .B(n13933), .Z(n13850) );
  OR U14167 ( .A(n13580), .B(n13579), .Z(n13584) );
  NANDN U14168 ( .A(n13582), .B(n13581), .Z(n13583) );
  AND U14169 ( .A(n13584), .B(n13583), .Z(n13849) );
  XNOR U14170 ( .A(n13850), .B(n13849), .Z(n13851) );
  XOR U14171 ( .A(n13852), .B(n13851), .Z(n13845) );
  XNOR U14172 ( .A(n13846), .B(n13845), .Z(n13938) );
  ANDN U14173 ( .B(o[17]), .A(n15818), .Z(n13937) );
  XOR U14174 ( .A(n13938), .B(n13937), .Z(n13939) );
  NANDN U14175 ( .A(n13586), .B(n13585), .Z(n13590) );
  OR U14176 ( .A(n13588), .B(n13587), .Z(n13589) );
  AND U14177 ( .A(n13590), .B(n13589), .Z(n13943) );
  XNOR U14178 ( .A(n13944), .B(n13943), .Z(n13946) );
  NANDN U14179 ( .A(n3012), .B(\stack[1][42] ), .Z(n13945) );
  XOR U14180 ( .A(n13946), .B(n13945), .Z(n13949) );
  XOR U14181 ( .A(n13950), .B(n13949), .Z(n13952) );
  OR U14182 ( .A(n13592), .B(n13591), .Z(n13596) );
  OR U14183 ( .A(n13594), .B(n13593), .Z(n13595) );
  AND U14184 ( .A(n13596), .B(n13595), .Z(n13951) );
  XNOR U14185 ( .A(n13952), .B(n13951), .Z(n13955) );
  NANDN U14186 ( .A(n13598), .B(n13597), .Z(n13602) );
  OR U14187 ( .A(n13600), .B(n13599), .Z(n13601) );
  AND U14188 ( .A(n13602), .B(n13601), .Z(n13956) );
  ANDN U14189 ( .B(o[20]), .A(n15935), .Z(n13957) );
  XOR U14190 ( .A(n13958), .B(n13957), .Z(n13961) );
  XOR U14191 ( .A(n13962), .B(n13961), .Z(n13964) );
  XNOR U14192 ( .A(n13963), .B(n13964), .Z(n13837) );
  XOR U14193 ( .A(n13838), .B(n13837), .Z(n13840) );
  XNOR U14194 ( .A(n13839), .B(n13840), .Z(n13833) );
  XOR U14195 ( .A(n13834), .B(n13833), .Z(n13826) );
  XOR U14196 ( .A(n13825), .B(n13826), .Z(n13827) );
  XOR U14197 ( .A(n13828), .B(n13827), .Z(n13970) );
  OR U14198 ( .A(n13604), .B(n13603), .Z(n13608) );
  NANDN U14199 ( .A(n13606), .B(n13605), .Z(n13607) );
  AND U14200 ( .A(n13608), .B(n13607), .Z(n13967) );
  AND U14201 ( .A(\stack[1][35] ), .B(o[25]), .Z(n13968) );
  XNOR U14202 ( .A(n13967), .B(n13968), .Z(n13969) );
  XOR U14203 ( .A(n13970), .B(n13969), .Z(n13819) );
  XNOR U14204 ( .A(n13820), .B(n13819), .Z(n13821) );
  XNOR U14205 ( .A(n13822), .B(n13821), .Z(n13815) );
  NANDN U14206 ( .A(n2990), .B(o[27]), .Z(n13813) );
  OR U14207 ( .A(n13610), .B(n13609), .Z(n13614) );
  OR U14208 ( .A(n13612), .B(n13611), .Z(n13613) );
  NAND U14209 ( .A(n13614), .B(n13613), .Z(n13814) );
  XOR U14210 ( .A(n13813), .B(n13814), .Z(n13816) );
  XNOR U14211 ( .A(n13815), .B(n13816), .Z(n13973) );
  XNOR U14212 ( .A(n13974), .B(n13973), .Z(n13975) );
  XOR U14213 ( .A(n13976), .B(n13975), .Z(n13809) );
  AND U14214 ( .A(o[29]), .B(\stack[1][31] ), .Z(n13807) );
  OR U14215 ( .A(n13616), .B(n13615), .Z(n13620) );
  OR U14216 ( .A(n13618), .B(n13617), .Z(n13619) );
  NAND U14217 ( .A(n13620), .B(n13619), .Z(n13808) );
  XNOR U14218 ( .A(n13807), .B(n13808), .Z(n13810) );
  XNOR U14219 ( .A(n13979), .B(n13980), .Z(n13982) );
  XOR U14220 ( .A(n13981), .B(n13982), .Z(n13803) );
  NANDN U14221 ( .A(n13622), .B(n13621), .Z(n13626) );
  OR U14222 ( .A(n13624), .B(n13623), .Z(n13625) );
  AND U14223 ( .A(n13626), .B(n13625), .Z(n13802) );
  NANDN U14224 ( .A(n2986), .B(o[31]), .Z(n13801) );
  XOR U14225 ( .A(n13802), .B(n13801), .Z(n13804) );
  XNOR U14226 ( .A(n13803), .B(n13804), .Z(n13985) );
  XNOR U14227 ( .A(n13986), .B(n13985), .Z(n13987) );
  XNOR U14228 ( .A(n13988), .B(n13987), .Z(n13797) );
  OR U14229 ( .A(n13628), .B(n13627), .Z(n13632) );
  NANDN U14230 ( .A(n13630), .B(n13629), .Z(n13631) );
  AND U14231 ( .A(n13632), .B(n13631), .Z(n13796) );
  NANDN U14232 ( .A(n2984), .B(o[33]), .Z(n13795) );
  XOR U14233 ( .A(n13796), .B(n13795), .Z(n13798) );
  XNOR U14234 ( .A(n13797), .B(n13798), .Z(n13991) );
  XNOR U14235 ( .A(n13992), .B(n13991), .Z(n13993) );
  XNOR U14236 ( .A(n13994), .B(n13993), .Z(n13791) );
  NANDN U14237 ( .A(n2982), .B(o[35]), .Z(n13789) );
  OR U14238 ( .A(n13634), .B(n13633), .Z(n13638) );
  OR U14239 ( .A(n13636), .B(n13635), .Z(n13637) );
  NAND U14240 ( .A(n13638), .B(n13637), .Z(n13790) );
  XOR U14241 ( .A(n13789), .B(n13790), .Z(n13792) );
  XNOR U14242 ( .A(n13791), .B(n13792), .Z(n13997) );
  XNOR U14243 ( .A(n13998), .B(n13997), .Z(n13999) );
  XNOR U14244 ( .A(n14000), .B(n13999), .Z(n13785) );
  NANDN U14245 ( .A(n2980), .B(o[37]), .Z(n13783) );
  OR U14246 ( .A(n13640), .B(n13639), .Z(n13644) );
  OR U14247 ( .A(n13642), .B(n13641), .Z(n13643) );
  NAND U14248 ( .A(n13644), .B(n13643), .Z(n13784) );
  XOR U14249 ( .A(n13783), .B(n13784), .Z(n13786) );
  XNOR U14250 ( .A(n13785), .B(n13786), .Z(n14003) );
  XNOR U14251 ( .A(n14004), .B(n14003), .Z(n14005) );
  XNOR U14252 ( .A(n14006), .B(n14005), .Z(n13779) );
  NANDN U14253 ( .A(n2978), .B(o[39]), .Z(n13777) );
  OR U14254 ( .A(n13646), .B(n13645), .Z(n13650) );
  OR U14255 ( .A(n13648), .B(n13647), .Z(n13649) );
  NAND U14256 ( .A(n13650), .B(n13649), .Z(n13778) );
  XOR U14257 ( .A(n13777), .B(n13778), .Z(n13780) );
  XNOR U14258 ( .A(n13779), .B(n13780), .Z(n14009) );
  XNOR U14259 ( .A(n14010), .B(n14009), .Z(n14011) );
  XNOR U14260 ( .A(n14012), .B(n14011), .Z(n13773) );
  NANDN U14261 ( .A(n16746), .B(o[41]), .Z(n13771) );
  OR U14262 ( .A(n13652), .B(n13651), .Z(n13656) );
  OR U14263 ( .A(n13654), .B(n13653), .Z(n13655) );
  NAND U14264 ( .A(n13656), .B(n13655), .Z(n13772) );
  XOR U14265 ( .A(n13771), .B(n13772), .Z(n13774) );
  XNOR U14266 ( .A(n13773), .B(n13774), .Z(n14015) );
  XNOR U14267 ( .A(n14016), .B(n14015), .Z(n14017) );
  XNOR U14268 ( .A(n14018), .B(n14017), .Z(n13767) );
  NANDN U14269 ( .A(n16826), .B(o[43]), .Z(n13765) );
  OR U14270 ( .A(n13658), .B(n13657), .Z(n13662) );
  OR U14271 ( .A(n13660), .B(n13659), .Z(n13661) );
  NAND U14272 ( .A(n13662), .B(n13661), .Z(n13766) );
  XOR U14273 ( .A(n13765), .B(n13766), .Z(n13768) );
  XNOR U14274 ( .A(n13767), .B(n13768), .Z(n14021) );
  XNOR U14275 ( .A(n14022), .B(n14021), .Z(n14023) );
  XNOR U14276 ( .A(n14024), .B(n14023), .Z(n13761) );
  NANDN U14277 ( .A(n2976), .B(o[45]), .Z(n13759) );
  OR U14278 ( .A(n13664), .B(n13663), .Z(n13668) );
  OR U14279 ( .A(n13666), .B(n13665), .Z(n13667) );
  NAND U14280 ( .A(n13668), .B(n13667), .Z(n13760) );
  XOR U14281 ( .A(n13759), .B(n13760), .Z(n13762) );
  XNOR U14282 ( .A(n13761), .B(n13762), .Z(n14027) );
  XNOR U14283 ( .A(n14028), .B(n14027), .Z(n14029) );
  XNOR U14284 ( .A(n14030), .B(n14029), .Z(n13755) );
  NANDN U14285 ( .A(n2974), .B(o[47]), .Z(n13753) );
  OR U14286 ( .A(n13670), .B(n13669), .Z(n13674) );
  OR U14287 ( .A(n13672), .B(n13671), .Z(n13673) );
  NAND U14288 ( .A(n13674), .B(n13673), .Z(n13754) );
  XOR U14289 ( .A(n13753), .B(n13754), .Z(n13756) );
  XNOR U14290 ( .A(n13755), .B(n13756), .Z(n14033) );
  XNOR U14291 ( .A(n14034), .B(n14033), .Z(n14035) );
  XNOR U14292 ( .A(n14036), .B(n14035), .Z(n13749) );
  NANDN U14293 ( .A(n2972), .B(o[49]), .Z(n13747) );
  OR U14294 ( .A(n13676), .B(n13675), .Z(n13680) );
  OR U14295 ( .A(n13678), .B(n13677), .Z(n13679) );
  NAND U14296 ( .A(n13680), .B(n13679), .Z(n13748) );
  XOR U14297 ( .A(n13747), .B(n13748), .Z(n13750) );
  XNOR U14298 ( .A(n13749), .B(n13750), .Z(n14039) );
  XNOR U14299 ( .A(n14040), .B(n14039), .Z(n14041) );
  XNOR U14300 ( .A(n14042), .B(n14041), .Z(n13743) );
  NANDN U14301 ( .A(n17145), .B(o[51]), .Z(n13741) );
  OR U14302 ( .A(n13682), .B(n13681), .Z(n13686) );
  OR U14303 ( .A(n13684), .B(n13683), .Z(n13685) );
  NAND U14304 ( .A(n13686), .B(n13685), .Z(n13742) );
  XOR U14305 ( .A(n13741), .B(n13742), .Z(n13744) );
  XNOR U14306 ( .A(n13743), .B(n13744), .Z(n14045) );
  XNOR U14307 ( .A(n14046), .B(n14045), .Z(n14047) );
  XNOR U14308 ( .A(n14048), .B(n14047), .Z(n13737) );
  NANDN U14309 ( .A(n17219), .B(o[53]), .Z(n13735) );
  OR U14310 ( .A(n13688), .B(n13687), .Z(n13692) );
  OR U14311 ( .A(n13690), .B(n13689), .Z(n13691) );
  NAND U14312 ( .A(n13692), .B(n13691), .Z(n13736) );
  XOR U14313 ( .A(n13735), .B(n13736), .Z(n13738) );
  XNOR U14314 ( .A(n13737), .B(n13738), .Z(n14051) );
  XNOR U14315 ( .A(n14052), .B(n14051), .Z(n14053) );
  XNOR U14316 ( .A(n14054), .B(n14053), .Z(n13731) );
  NANDN U14317 ( .A(n17296), .B(o[55]), .Z(n13729) );
  OR U14318 ( .A(n13694), .B(n13693), .Z(n13698) );
  OR U14319 ( .A(n13696), .B(n13695), .Z(n13697) );
  NAND U14320 ( .A(n13698), .B(n13697), .Z(n13730) );
  XOR U14321 ( .A(n13729), .B(n13730), .Z(n13732) );
  XNOR U14322 ( .A(n13731), .B(n13732), .Z(n14057) );
  XNOR U14323 ( .A(n14058), .B(n14057), .Z(n14059) );
  XNOR U14324 ( .A(n14060), .B(n14059), .Z(n13725) );
  NANDN U14325 ( .A(n17375), .B(o[57]), .Z(n13723) );
  OR U14326 ( .A(n13700), .B(n13699), .Z(n13704) );
  OR U14327 ( .A(n13702), .B(n13701), .Z(n13703) );
  NAND U14328 ( .A(n13704), .B(n13703), .Z(n13724) );
  XOR U14329 ( .A(n13723), .B(n13724), .Z(n13726) );
  XNOR U14330 ( .A(n13725), .B(n13726), .Z(n14063) );
  XNOR U14331 ( .A(n14064), .B(n14063), .Z(n14065) );
  AND U14332 ( .A(o[59]), .B(\stack[1][1] ), .Z(n13717) );
  OR U14333 ( .A(n13706), .B(n13705), .Z(n13710) );
  OR U14334 ( .A(n13708), .B(n13707), .Z(n13709) );
  NAND U14335 ( .A(n13710), .B(n13709), .Z(n13718) );
  XNOR U14336 ( .A(n13717), .B(n13718), .Z(n13720) );
  XOR U14337 ( .A(n13719), .B(n13720), .Z(n13711) );
  NANDN U14338 ( .A(n13712), .B(n13711), .Z(n13714) );
  XOR U14339 ( .A(n13712), .B(n13711), .Z(n15163) );
  AND U14340 ( .A(o[60]), .B(\stack[1][0] ), .Z(n15164) );
  OR U14341 ( .A(n15163), .B(n15164), .Z(n13713) );
  AND U14342 ( .A(n13714), .B(n13713), .Z(n13716) );
  OR U14343 ( .A(n13715), .B(n13716), .Z(n14070) );
  XNOR U14344 ( .A(n13716), .B(n13715), .Z(n15124) );
  NANDN U14345 ( .A(n2969), .B(o[60]), .Z(n14427) );
  OR U14346 ( .A(n13718), .B(n13717), .Z(n13722) );
  OR U14347 ( .A(n13720), .B(n13719), .Z(n13721) );
  NAND U14348 ( .A(n13722), .B(n13721), .Z(n14425) );
  NANDN U14349 ( .A(n17375), .B(o[58]), .Z(n14421) );
  NANDN U14350 ( .A(n13724), .B(n13723), .Z(n13728) );
  NANDN U14351 ( .A(n13726), .B(n13725), .Z(n13727) );
  NAND U14352 ( .A(n13728), .B(n13727), .Z(n14419) );
  NANDN U14353 ( .A(n17296), .B(o[56]), .Z(n14415) );
  NANDN U14354 ( .A(n13730), .B(n13729), .Z(n13734) );
  NANDN U14355 ( .A(n13732), .B(n13731), .Z(n13733) );
  NAND U14356 ( .A(n13734), .B(n13733), .Z(n14413) );
  NANDN U14357 ( .A(n17219), .B(o[54]), .Z(n14409) );
  NANDN U14358 ( .A(n13736), .B(n13735), .Z(n13740) );
  NANDN U14359 ( .A(n13738), .B(n13737), .Z(n13739) );
  NAND U14360 ( .A(n13740), .B(n13739), .Z(n14407) );
  NANDN U14361 ( .A(n17145), .B(o[52]), .Z(n14403) );
  NANDN U14362 ( .A(n13742), .B(n13741), .Z(n13746) );
  NANDN U14363 ( .A(n13744), .B(n13743), .Z(n13745) );
  NAND U14364 ( .A(n13746), .B(n13745), .Z(n14401) );
  NANDN U14365 ( .A(n2972), .B(o[50]), .Z(n14397) );
  NANDN U14366 ( .A(n13748), .B(n13747), .Z(n13752) );
  NANDN U14367 ( .A(n13750), .B(n13749), .Z(n13751) );
  NAND U14368 ( .A(n13752), .B(n13751), .Z(n14395) );
  NANDN U14369 ( .A(n2974), .B(o[48]), .Z(n14391) );
  NANDN U14370 ( .A(n13754), .B(n13753), .Z(n13758) );
  NANDN U14371 ( .A(n13756), .B(n13755), .Z(n13757) );
  NAND U14372 ( .A(n13758), .B(n13757), .Z(n14389) );
  NANDN U14373 ( .A(n2976), .B(o[46]), .Z(n14385) );
  NANDN U14374 ( .A(n13760), .B(n13759), .Z(n13764) );
  NANDN U14375 ( .A(n13762), .B(n13761), .Z(n13763) );
  NAND U14376 ( .A(n13764), .B(n13763), .Z(n14383) );
  NANDN U14377 ( .A(n16826), .B(o[44]), .Z(n14379) );
  NANDN U14378 ( .A(n13766), .B(n13765), .Z(n13770) );
  NANDN U14379 ( .A(n13768), .B(n13767), .Z(n13769) );
  NAND U14380 ( .A(n13770), .B(n13769), .Z(n14377) );
  NANDN U14381 ( .A(n16746), .B(o[42]), .Z(n14373) );
  NANDN U14382 ( .A(n13772), .B(n13771), .Z(n13776) );
  NANDN U14383 ( .A(n13774), .B(n13773), .Z(n13775) );
  NAND U14384 ( .A(n13776), .B(n13775), .Z(n14371) );
  NANDN U14385 ( .A(n2978), .B(o[40]), .Z(n14367) );
  NANDN U14386 ( .A(n13778), .B(n13777), .Z(n13782) );
  NANDN U14387 ( .A(n13780), .B(n13779), .Z(n13781) );
  NAND U14388 ( .A(n13782), .B(n13781), .Z(n14365) );
  NANDN U14389 ( .A(n2980), .B(o[38]), .Z(n14361) );
  NANDN U14390 ( .A(n13784), .B(n13783), .Z(n13788) );
  NANDN U14391 ( .A(n13786), .B(n13785), .Z(n13787) );
  NAND U14392 ( .A(n13788), .B(n13787), .Z(n14359) );
  NANDN U14393 ( .A(n2982), .B(o[36]), .Z(n14355) );
  NANDN U14394 ( .A(n13790), .B(n13789), .Z(n13794) );
  NANDN U14395 ( .A(n13792), .B(n13791), .Z(n13793) );
  NAND U14396 ( .A(n13794), .B(n13793), .Z(n14353) );
  NANDN U14397 ( .A(n2984), .B(o[34]), .Z(n14349) );
  NANDN U14398 ( .A(n13796), .B(n13795), .Z(n13800) );
  NANDN U14399 ( .A(n13798), .B(n13797), .Z(n13799) );
  NAND U14400 ( .A(n13800), .B(n13799), .Z(n14347) );
  NANDN U14401 ( .A(n2986), .B(o[32]), .Z(n14343) );
  NANDN U14402 ( .A(n13802), .B(n13801), .Z(n13806) );
  NANDN U14403 ( .A(n13804), .B(n13803), .Z(n13805) );
  NAND U14404 ( .A(n13806), .B(n13805), .Z(n14341) );
  NANDN U14405 ( .A(n2988), .B(o[30]), .Z(n14337) );
  OR U14406 ( .A(n13808), .B(n13807), .Z(n13812) );
  OR U14407 ( .A(n13810), .B(n13809), .Z(n13811) );
  NAND U14408 ( .A(n13812), .B(n13811), .Z(n14335) );
  AND U14409 ( .A(\stack[1][33] ), .B(o[28]), .Z(n14331) );
  NANDN U14410 ( .A(n13814), .B(n13813), .Z(n13818) );
  NANDN U14411 ( .A(n13816), .B(n13815), .Z(n13817) );
  AND U14412 ( .A(n13818), .B(n13817), .Z(n14328) );
  AND U14413 ( .A(o[27]), .B(\stack[1][34] ), .Z(n14167) );
  OR U14414 ( .A(n13820), .B(n13819), .Z(n13824) );
  OR U14415 ( .A(n13822), .B(n13821), .Z(n13823) );
  NAND U14416 ( .A(n13824), .B(n13823), .Z(n14168) );
  XNOR U14417 ( .A(n14167), .B(n14168), .Z(n14170) );
  OR U14418 ( .A(n13826), .B(n13825), .Z(n13830) );
  NANDN U14419 ( .A(n13828), .B(n13827), .Z(n13829) );
  NAND U14420 ( .A(n13830), .B(n13829), .Z(n14174) );
  ANDN U14421 ( .B(o[25]), .A(n2993), .Z(n14173) );
  XOR U14422 ( .A(n14174), .B(n14173), .Z(n14175) );
  OR U14423 ( .A(n13832), .B(n13831), .Z(n13836) );
  NANDN U14424 ( .A(n13834), .B(n13833), .Z(n13835) );
  NAND U14425 ( .A(n13836), .B(n13835), .Z(n14180) );
  ANDN U14426 ( .B(\stack[1][38] ), .A(n3017), .Z(n14188) );
  NANDN U14427 ( .A(n13838), .B(n13837), .Z(n13842) );
  NANDN U14428 ( .A(n13840), .B(n13839), .Z(n13841) );
  AND U14429 ( .A(n13842), .B(n13841), .Z(n14185) );
  AND U14430 ( .A(\stack[1][39] ), .B(o[22]), .Z(n14319) );
  AND U14431 ( .A(\stack[1][40] ), .B(o[21]), .Z(n14312) );
  OR U14432 ( .A(n13844), .B(n13843), .Z(n13848) );
  NAND U14433 ( .A(n13846), .B(n13845), .Z(n13847) );
  AND U14434 ( .A(n13848), .B(n13847), .Z(n14289) );
  OR U14435 ( .A(n13850), .B(n13849), .Z(n13854) );
  OR U14436 ( .A(n13852), .B(n13851), .Z(n13853) );
  AND U14437 ( .A(n13854), .B(n13853), .Z(n14191) );
  NANDN U14438 ( .A(n3010), .B(\stack[1][45] ), .Z(n14192) );
  XOR U14439 ( .A(n14191), .B(n14192), .Z(n14194) );
  NANDN U14440 ( .A(n3009), .B(\stack[1][46] ), .Z(n14200) );
  OR U14441 ( .A(n13856), .B(n13855), .Z(n13860) );
  OR U14442 ( .A(n13858), .B(n13857), .Z(n13859) );
  AND U14443 ( .A(n13860), .B(n13859), .Z(n14276) );
  NANDN U14444 ( .A(n13862), .B(n13861), .Z(n13866) );
  NANDN U14445 ( .A(n13864), .B(n13863), .Z(n13865) );
  NAND U14446 ( .A(n13866), .B(n13865), .Z(n14204) );
  AND U14447 ( .A(\stack[1][50] ), .B(o[11]), .Z(n14212) );
  OR U14448 ( .A(n13868), .B(n13867), .Z(n13872) );
  NANDN U14449 ( .A(n13870), .B(n13869), .Z(n13871) );
  AND U14450 ( .A(n13872), .B(n13871), .Z(n14209) );
  AND U14451 ( .A(\stack[1][51] ), .B(o[10]), .Z(n14218) );
  AND U14452 ( .A(\stack[1][52] ), .B(o[9]), .Z(n14270) );
  NANDN U14453 ( .A(n13874), .B(n13873), .Z(n13878) );
  NAND U14454 ( .A(n13876), .B(n13875), .Z(n13877) );
  AND U14455 ( .A(n13878), .B(n13877), .Z(n14259) );
  AND U14456 ( .A(\stack[1][56] ), .B(o[5]), .Z(n14253) );
  OR U14457 ( .A(n13880), .B(n13879), .Z(n13884) );
  NANDN U14458 ( .A(n13882), .B(n13881), .Z(n13883) );
  AND U14459 ( .A(n13884), .B(n13883), .Z(n14250) );
  ANDN U14460 ( .B(\stack[1][57] ), .A(n2998), .Z(n14230) );
  AND U14461 ( .A(\stack[1][58] ), .B(o[3]), .Z(n14247) );
  NANDN U14462 ( .A(n13885), .B(n14233), .Z(n13886) );
  AND U14463 ( .A(n13887), .B(n13886), .Z(n13891) );
  OR U14464 ( .A(n13889), .B(n13888), .Z(n13890) );
  AND U14465 ( .A(n13891), .B(n13890), .Z(n14244) );
  NANDN U14466 ( .A(n2995), .B(\stack[1][61] ), .Z(n14242) );
  NOR U14467 ( .A(n13892), .B(n14242), .Z(n14679) );
  XNOR U14468 ( .A(n14679), .B(n14233), .Z(n13894) );
  NAND U14469 ( .A(o[0]), .B(\stack[1][61] ), .Z(n14240) );
  NANDN U14470 ( .A(n13893), .B(n14240), .Z(n14235) );
  NAND U14471 ( .A(n13894), .B(n14235), .Z(n14237) );
  AND U14472 ( .A(\stack[1][59] ), .B(o[2]), .Z(n14236) );
  XNOR U14473 ( .A(n14237), .B(n14236), .Z(n14245) );
  XOR U14474 ( .A(n14244), .B(n14245), .Z(n14246) );
  XOR U14475 ( .A(n14247), .B(n14246), .Z(n14228) );
  OR U14476 ( .A(n13896), .B(n13895), .Z(n13900) );
  NANDN U14477 ( .A(n13898), .B(n13897), .Z(n13899) );
  AND U14478 ( .A(n13900), .B(n13899), .Z(n14227) );
  XOR U14479 ( .A(n14228), .B(n14227), .Z(n14229) );
  XOR U14480 ( .A(n14230), .B(n14229), .Z(n14251) );
  XNOR U14481 ( .A(n14250), .B(n14251), .Z(n14252) );
  OR U14482 ( .A(n13902), .B(n13901), .Z(n13906) );
  OR U14483 ( .A(n13904), .B(n13903), .Z(n13905) );
  NAND U14484 ( .A(n13906), .B(n13905), .Z(n14222) );
  ANDN U14485 ( .B(\stack[1][55] ), .A(n3000), .Z(n14221) );
  XNOR U14486 ( .A(n14222), .B(n14221), .Z(n14224) );
  XNOR U14487 ( .A(n14223), .B(n14224), .Z(n14257) );
  ANDN U14488 ( .B(\stack[1][54] ), .A(n3001), .Z(n14256) );
  XOR U14489 ( .A(n14257), .B(n14256), .Z(n14258) );
  NANDN U14490 ( .A(n13908), .B(n13907), .Z(n13912) );
  OR U14491 ( .A(n13910), .B(n13909), .Z(n13911) );
  AND U14492 ( .A(n13912), .B(n13911), .Z(n14262) );
  XNOR U14493 ( .A(n14263), .B(n14262), .Z(n14265) );
  ANDN U14494 ( .B(\stack[1][53] ), .A(n3002), .Z(n14264) );
  XNOR U14495 ( .A(n14265), .B(n14264), .Z(n14268) );
  OR U14496 ( .A(n13914), .B(n13913), .Z(n13918) );
  NANDN U14497 ( .A(n13916), .B(n13915), .Z(n13917) );
  NAND U14498 ( .A(n13918), .B(n13917), .Z(n14269) );
  XNOR U14499 ( .A(n14268), .B(n14269), .Z(n14271) );
  XNOR U14500 ( .A(n14270), .B(n14271), .Z(n14216) );
  OR U14501 ( .A(n13920), .B(n13919), .Z(n13924) );
  OR U14502 ( .A(n13922), .B(n13921), .Z(n13923) );
  AND U14503 ( .A(n13924), .B(n13923), .Z(n14215) );
  XOR U14504 ( .A(n14216), .B(n14215), .Z(n14217) );
  XOR U14505 ( .A(n14218), .B(n14217), .Z(n14210) );
  XNOR U14506 ( .A(n14209), .B(n14210), .Z(n14211) );
  XOR U14507 ( .A(n14204), .B(n14203), .Z(n14206) );
  ANDN U14508 ( .B(\stack[1][49] ), .A(n3006), .Z(n14205) );
  XOR U14509 ( .A(n14206), .B(n14205), .Z(n14275) );
  ANDN U14510 ( .B(o[13]), .A(n15623), .Z(n14274) );
  XOR U14511 ( .A(n14275), .B(n14274), .Z(n14277) );
  XNOR U14512 ( .A(n14276), .B(n14277), .Z(n14281) );
  NANDN U14513 ( .A(n13926), .B(n13925), .Z(n13930) );
  OR U14514 ( .A(n13928), .B(n13927), .Z(n13929) );
  AND U14515 ( .A(n13930), .B(n13929), .Z(n14280) );
  XNOR U14516 ( .A(n14281), .B(n14280), .Z(n14283) );
  ANDN U14517 ( .B(o[14]), .A(n15662), .Z(n14282) );
  XOR U14518 ( .A(n14283), .B(n14282), .Z(n14198) );
  OR U14519 ( .A(n13932), .B(n13931), .Z(n13936) );
  NANDN U14520 ( .A(n13934), .B(n13933), .Z(n13935) );
  AND U14521 ( .A(n13936), .B(n13935), .Z(n14197) );
  XNOR U14522 ( .A(n14198), .B(n14197), .Z(n14199) );
  XOR U14523 ( .A(n14200), .B(n14199), .Z(n14193) );
  XNOR U14524 ( .A(n14194), .B(n14193), .Z(n14287) );
  ANDN U14525 ( .B(o[17]), .A(n15779), .Z(n14286) );
  XOR U14526 ( .A(n14287), .B(n14286), .Z(n14288) );
  NANDN U14527 ( .A(n13938), .B(n13937), .Z(n13942) );
  OR U14528 ( .A(n13940), .B(n13939), .Z(n13941) );
  AND U14529 ( .A(n13942), .B(n13941), .Z(n14292) );
  XNOR U14530 ( .A(n14293), .B(n14292), .Z(n14295) );
  ANDN U14531 ( .B(o[18]), .A(n15818), .Z(n14294) );
  XOR U14532 ( .A(n14295), .B(n14294), .Z(n14299) );
  OR U14533 ( .A(n13944), .B(n13943), .Z(n13948) );
  OR U14534 ( .A(n13946), .B(n13945), .Z(n13947) );
  AND U14535 ( .A(n13948), .B(n13947), .Z(n14298) );
  XNOR U14536 ( .A(n14299), .B(n14298), .Z(n14301) );
  ANDN U14537 ( .B(o[19]), .A(n15857), .Z(n14300) );
  XOR U14538 ( .A(n14301), .B(n14300), .Z(n14305) );
  NANDN U14539 ( .A(n13950), .B(n13949), .Z(n13954) );
  OR U14540 ( .A(n13952), .B(n13951), .Z(n13953) );
  AND U14541 ( .A(n13954), .B(n13953), .Z(n14304) );
  XNOR U14542 ( .A(n14305), .B(n14304), .Z(n14307) );
  AND U14543 ( .A(\stack[1][41] ), .B(o[20]), .Z(n14306) );
  XNOR U14544 ( .A(n14307), .B(n14306), .Z(n14310) );
  OR U14545 ( .A(n13956), .B(n13955), .Z(n13960) );
  NANDN U14546 ( .A(n13958), .B(n13957), .Z(n13959) );
  NAND U14547 ( .A(n13960), .B(n13959), .Z(n14311) );
  XNOR U14548 ( .A(n14310), .B(n14311), .Z(n14313) );
  XNOR U14549 ( .A(n14312), .B(n14313), .Z(n14317) );
  NANDN U14550 ( .A(n13962), .B(n13961), .Z(n13966) );
  NANDN U14551 ( .A(n13964), .B(n13963), .Z(n13965) );
  AND U14552 ( .A(n13966), .B(n13965), .Z(n14316) );
  XOR U14553 ( .A(n14317), .B(n14316), .Z(n14318) );
  XOR U14554 ( .A(n14319), .B(n14318), .Z(n14186) );
  XNOR U14555 ( .A(n14185), .B(n14186), .Z(n14187) );
  XOR U14556 ( .A(n14180), .B(n14179), .Z(n14182) );
  NANDN U14557 ( .A(n3018), .B(\stack[1][37] ), .Z(n14181) );
  XNOR U14558 ( .A(n14182), .B(n14181), .Z(n14176) );
  OR U14559 ( .A(n13968), .B(n13967), .Z(n13972) );
  OR U14560 ( .A(n13970), .B(n13969), .Z(n13971) );
  AND U14561 ( .A(n13972), .B(n13971), .Z(n14323) );
  XNOR U14562 ( .A(n14322), .B(n14323), .Z(n14325) );
  AND U14563 ( .A(\stack[1][35] ), .B(o[26]), .Z(n14324) );
  XOR U14564 ( .A(n14325), .B(n14324), .Z(n14169) );
  XOR U14565 ( .A(n14170), .B(n14169), .Z(n14329) );
  XOR U14566 ( .A(n14328), .B(n14329), .Z(n14330) );
  XOR U14567 ( .A(n14331), .B(n14330), .Z(n14164) );
  AND U14568 ( .A(o[29]), .B(\stack[1][32] ), .Z(n14161) );
  OR U14569 ( .A(n13974), .B(n13973), .Z(n13978) );
  OR U14570 ( .A(n13976), .B(n13975), .Z(n13977) );
  NAND U14571 ( .A(n13978), .B(n13977), .Z(n14162) );
  XNOR U14572 ( .A(n14161), .B(n14162), .Z(n14163) );
  XOR U14573 ( .A(n14164), .B(n14163), .Z(n14334) );
  XNOR U14574 ( .A(n14335), .B(n14334), .Z(n14336) );
  XNOR U14575 ( .A(n14337), .B(n14336), .Z(n14157) );
  NANDN U14576 ( .A(n2987), .B(o[31]), .Z(n14155) );
  OR U14577 ( .A(n13980), .B(n13979), .Z(n13984) );
  IV U14578 ( .A(n13981), .Z(n16317) );
  OR U14579 ( .A(n13982), .B(n16317), .Z(n13983) );
  NAND U14580 ( .A(n13984), .B(n13983), .Z(n14156) );
  XOR U14581 ( .A(n14155), .B(n14156), .Z(n14158) );
  XNOR U14582 ( .A(n14157), .B(n14158), .Z(n14340) );
  XNOR U14583 ( .A(n14341), .B(n14340), .Z(n14342) );
  XNOR U14584 ( .A(n14343), .B(n14342), .Z(n14151) );
  NANDN U14585 ( .A(n2985), .B(o[33]), .Z(n14149) );
  OR U14586 ( .A(n13986), .B(n13985), .Z(n13990) );
  OR U14587 ( .A(n13988), .B(n13987), .Z(n13989) );
  NAND U14588 ( .A(n13990), .B(n13989), .Z(n14150) );
  XOR U14589 ( .A(n14149), .B(n14150), .Z(n14152) );
  XNOR U14590 ( .A(n14151), .B(n14152), .Z(n14346) );
  XNOR U14591 ( .A(n14347), .B(n14346), .Z(n14348) );
  XNOR U14592 ( .A(n14349), .B(n14348), .Z(n14145) );
  NANDN U14593 ( .A(n2983), .B(o[35]), .Z(n14143) );
  OR U14594 ( .A(n13992), .B(n13991), .Z(n13996) );
  OR U14595 ( .A(n13994), .B(n13993), .Z(n13995) );
  NAND U14596 ( .A(n13996), .B(n13995), .Z(n14144) );
  XOR U14597 ( .A(n14143), .B(n14144), .Z(n14146) );
  XNOR U14598 ( .A(n14145), .B(n14146), .Z(n14352) );
  XNOR U14599 ( .A(n14353), .B(n14352), .Z(n14354) );
  XNOR U14600 ( .A(n14355), .B(n14354), .Z(n14139) );
  NANDN U14601 ( .A(n2981), .B(o[37]), .Z(n14137) );
  OR U14602 ( .A(n13998), .B(n13997), .Z(n14002) );
  OR U14603 ( .A(n14000), .B(n13999), .Z(n14001) );
  NAND U14604 ( .A(n14002), .B(n14001), .Z(n14138) );
  XOR U14605 ( .A(n14137), .B(n14138), .Z(n14140) );
  XNOR U14606 ( .A(n14139), .B(n14140), .Z(n14358) );
  XNOR U14607 ( .A(n14359), .B(n14358), .Z(n14360) );
  XNOR U14608 ( .A(n14361), .B(n14360), .Z(n14133) );
  NANDN U14609 ( .A(n2979), .B(o[39]), .Z(n14131) );
  OR U14610 ( .A(n14004), .B(n14003), .Z(n14008) );
  OR U14611 ( .A(n14006), .B(n14005), .Z(n14007) );
  NAND U14612 ( .A(n14008), .B(n14007), .Z(n14132) );
  XOR U14613 ( .A(n14131), .B(n14132), .Z(n14134) );
  XNOR U14614 ( .A(n14133), .B(n14134), .Z(n14364) );
  XNOR U14615 ( .A(n14365), .B(n14364), .Z(n14366) );
  XNOR U14616 ( .A(n14367), .B(n14366), .Z(n14127) );
  NANDN U14617 ( .A(n16712), .B(o[41]), .Z(n14125) );
  OR U14618 ( .A(n14010), .B(n14009), .Z(n14014) );
  OR U14619 ( .A(n14012), .B(n14011), .Z(n14013) );
  NAND U14620 ( .A(n14014), .B(n14013), .Z(n14126) );
  XOR U14621 ( .A(n14125), .B(n14126), .Z(n14128) );
  XNOR U14622 ( .A(n14127), .B(n14128), .Z(n14370) );
  XNOR U14623 ( .A(n14371), .B(n14370), .Z(n14372) );
  XNOR U14624 ( .A(n14373), .B(n14372), .Z(n14121) );
  NANDN U14625 ( .A(n16786), .B(o[43]), .Z(n14119) );
  OR U14626 ( .A(n14016), .B(n14015), .Z(n14020) );
  OR U14627 ( .A(n14018), .B(n14017), .Z(n14019) );
  NAND U14628 ( .A(n14020), .B(n14019), .Z(n14120) );
  XOR U14629 ( .A(n14119), .B(n14120), .Z(n14122) );
  XNOR U14630 ( .A(n14121), .B(n14122), .Z(n14376) );
  XNOR U14631 ( .A(n14377), .B(n14376), .Z(n14378) );
  XNOR U14632 ( .A(n14379), .B(n14378), .Z(n14115) );
  NANDN U14633 ( .A(n2977), .B(o[45]), .Z(n14113) );
  OR U14634 ( .A(n14022), .B(n14021), .Z(n14026) );
  OR U14635 ( .A(n14024), .B(n14023), .Z(n14025) );
  NAND U14636 ( .A(n14026), .B(n14025), .Z(n14114) );
  XOR U14637 ( .A(n14113), .B(n14114), .Z(n14116) );
  XNOR U14638 ( .A(n14115), .B(n14116), .Z(n14382) );
  XNOR U14639 ( .A(n14383), .B(n14382), .Z(n14384) );
  XNOR U14640 ( .A(n14385), .B(n14384), .Z(n14109) );
  NANDN U14641 ( .A(n2975), .B(o[47]), .Z(n14107) );
  OR U14642 ( .A(n14028), .B(n14027), .Z(n14032) );
  OR U14643 ( .A(n14030), .B(n14029), .Z(n14031) );
  NAND U14644 ( .A(n14032), .B(n14031), .Z(n14108) );
  XOR U14645 ( .A(n14107), .B(n14108), .Z(n14110) );
  XNOR U14646 ( .A(n14109), .B(n14110), .Z(n14388) );
  XNOR U14647 ( .A(n14389), .B(n14388), .Z(n14390) );
  XNOR U14648 ( .A(n14391), .B(n14390), .Z(n14103) );
  NANDN U14649 ( .A(n2973), .B(o[49]), .Z(n14101) );
  OR U14650 ( .A(n14034), .B(n14033), .Z(n14038) );
  OR U14651 ( .A(n14036), .B(n14035), .Z(n14037) );
  NAND U14652 ( .A(n14038), .B(n14037), .Z(n14102) );
  XOR U14653 ( .A(n14101), .B(n14102), .Z(n14104) );
  XNOR U14654 ( .A(n14103), .B(n14104), .Z(n14394) );
  XNOR U14655 ( .A(n14395), .B(n14394), .Z(n14396) );
  XNOR U14656 ( .A(n14397), .B(n14396), .Z(n14097) );
  NANDN U14657 ( .A(n17101), .B(o[51]), .Z(n14095) );
  OR U14658 ( .A(n14040), .B(n14039), .Z(n14044) );
  OR U14659 ( .A(n14042), .B(n14041), .Z(n14043) );
  NAND U14660 ( .A(n14044), .B(n14043), .Z(n14096) );
  XOR U14661 ( .A(n14095), .B(n14096), .Z(n14098) );
  XNOR U14662 ( .A(n14097), .B(n14098), .Z(n14400) );
  XNOR U14663 ( .A(n14401), .B(n14400), .Z(n14402) );
  XNOR U14664 ( .A(n14403), .B(n14402), .Z(n14091) );
  NANDN U14665 ( .A(n17179), .B(o[53]), .Z(n14089) );
  OR U14666 ( .A(n14046), .B(n14045), .Z(n14050) );
  OR U14667 ( .A(n14048), .B(n14047), .Z(n14049) );
  NAND U14668 ( .A(n14050), .B(n14049), .Z(n14090) );
  XOR U14669 ( .A(n14089), .B(n14090), .Z(n14092) );
  XNOR U14670 ( .A(n14091), .B(n14092), .Z(n14406) );
  XNOR U14671 ( .A(n14407), .B(n14406), .Z(n14408) );
  XNOR U14672 ( .A(n14409), .B(n14408), .Z(n14085) );
  NANDN U14673 ( .A(n17256), .B(o[55]), .Z(n14083) );
  OR U14674 ( .A(n14052), .B(n14051), .Z(n14056) );
  OR U14675 ( .A(n14054), .B(n14053), .Z(n14055) );
  NAND U14676 ( .A(n14056), .B(n14055), .Z(n14084) );
  XOR U14677 ( .A(n14083), .B(n14084), .Z(n14086) );
  XNOR U14678 ( .A(n14085), .B(n14086), .Z(n14412) );
  XNOR U14679 ( .A(n14413), .B(n14412), .Z(n14414) );
  XNOR U14680 ( .A(n14415), .B(n14414), .Z(n14079) );
  AND U14681 ( .A(o[57]), .B(\stack[1][4] ), .Z(n14077) );
  OR U14682 ( .A(n14058), .B(n14057), .Z(n14062) );
  OR U14683 ( .A(n14060), .B(n14059), .Z(n14061) );
  NAND U14684 ( .A(n14062), .B(n14061), .Z(n14078) );
  XNOR U14685 ( .A(n14077), .B(n14078), .Z(n14080) );
  XNOR U14686 ( .A(n14079), .B(n14080), .Z(n14418) );
  XNOR U14687 ( .A(n14419), .B(n14418), .Z(n14420) );
  XOR U14688 ( .A(n14421), .B(n14420), .Z(n14074) );
  AND U14689 ( .A(o[59]), .B(\stack[1][2] ), .Z(n14071) );
  OR U14690 ( .A(n14064), .B(n14063), .Z(n14068) );
  OR U14691 ( .A(n14066), .B(n14065), .Z(n14067) );
  NAND U14692 ( .A(n14068), .B(n14067), .Z(n14072) );
  XOR U14693 ( .A(n14071), .B(n14072), .Z(n14073) );
  XNOR U14694 ( .A(n14074), .B(n14073), .Z(n14424) );
  XNOR U14695 ( .A(n14425), .B(n14424), .Z(n14426) );
  XOR U14696 ( .A(n14427), .B(n14426), .Z(n15125) );
  OR U14697 ( .A(n15124), .B(n15125), .Z(n14069) );
  AND U14698 ( .A(n14070), .B(n14069), .Z(n14430) );
  NANDN U14699 ( .A(n2970), .B(o[60]), .Z(n15035) );
  OR U14700 ( .A(n14072), .B(n14071), .Z(n14076) );
  NANDN U14701 ( .A(n14074), .B(n14073), .Z(n14075) );
  NAND U14702 ( .A(n14076), .B(n14075), .Z(n15034) );
  NANDN U14703 ( .A(n2971), .B(o[58]), .Z(n14435) );
  OR U14704 ( .A(n14078), .B(n14077), .Z(n14082) );
  NANDN U14705 ( .A(n14080), .B(n14079), .Z(n14081) );
  NAND U14706 ( .A(n14082), .B(n14081), .Z(n14437) );
  NANDN U14707 ( .A(n17256), .B(o[56]), .Z(n14992) );
  NANDN U14708 ( .A(n14084), .B(n14083), .Z(n14088) );
  NANDN U14709 ( .A(n14086), .B(n14085), .Z(n14087) );
  NAND U14710 ( .A(n14088), .B(n14087), .Z(n14994) );
  NANDN U14711 ( .A(n17179), .B(o[54]), .Z(n14441) );
  NANDN U14712 ( .A(n14090), .B(n14089), .Z(n14094) );
  NANDN U14713 ( .A(n14092), .B(n14091), .Z(n14093) );
  NAND U14714 ( .A(n14094), .B(n14093), .Z(n14443) );
  NANDN U14715 ( .A(n17101), .B(o[52]), .Z(n14447) );
  NANDN U14716 ( .A(n14096), .B(n14095), .Z(n14100) );
  NANDN U14717 ( .A(n14098), .B(n14097), .Z(n14099) );
  NAND U14718 ( .A(n14100), .B(n14099), .Z(n14449) );
  NANDN U14719 ( .A(n2973), .B(o[50]), .Z(n14453) );
  NANDN U14720 ( .A(n14102), .B(n14101), .Z(n14106) );
  NANDN U14721 ( .A(n14104), .B(n14103), .Z(n14105) );
  NAND U14722 ( .A(n14106), .B(n14105), .Z(n14455) );
  NANDN U14723 ( .A(n2975), .B(o[48]), .Z(n14962) );
  NANDN U14724 ( .A(n14108), .B(n14107), .Z(n14112) );
  NANDN U14725 ( .A(n14110), .B(n14109), .Z(n14111) );
  NAND U14726 ( .A(n14112), .B(n14111), .Z(n14964) );
  NANDN U14727 ( .A(n2977), .B(o[46]), .Z(n14944) );
  NANDN U14728 ( .A(n14114), .B(n14113), .Z(n14118) );
  NANDN U14729 ( .A(n14116), .B(n14115), .Z(n14117) );
  NAND U14730 ( .A(n14118), .B(n14117), .Z(n14946) );
  NANDN U14731 ( .A(n16786), .B(o[44]), .Z(n14920) );
  NANDN U14732 ( .A(n14120), .B(n14119), .Z(n14124) );
  NANDN U14733 ( .A(n14122), .B(n14121), .Z(n14123) );
  NAND U14734 ( .A(n14124), .B(n14123), .Z(n14922) );
  NANDN U14735 ( .A(n16712), .B(o[42]), .Z(n14926) );
  NANDN U14736 ( .A(n14126), .B(n14125), .Z(n14130) );
  NANDN U14737 ( .A(n14128), .B(n14127), .Z(n14129) );
  NAND U14738 ( .A(n14130), .B(n14129), .Z(n14928) );
  NANDN U14739 ( .A(n2979), .B(o[40]), .Z(n14909) );
  NANDN U14740 ( .A(n14132), .B(n14131), .Z(n14136) );
  NANDN U14741 ( .A(n14134), .B(n14133), .Z(n14135) );
  NAND U14742 ( .A(n14136), .B(n14135), .Z(n14908) );
  NANDN U14743 ( .A(n2981), .B(o[38]), .Z(n14884) );
  NANDN U14744 ( .A(n14138), .B(n14137), .Z(n14142) );
  NANDN U14745 ( .A(n14140), .B(n14139), .Z(n14141) );
  NAND U14746 ( .A(n14142), .B(n14141), .Z(n14886) );
  NANDN U14747 ( .A(n2983), .B(o[36]), .Z(n14477) );
  NANDN U14748 ( .A(n14144), .B(n14143), .Z(n14148) );
  NANDN U14749 ( .A(n14146), .B(n14145), .Z(n14147) );
  NAND U14750 ( .A(n14148), .B(n14147), .Z(n14479) );
  NANDN U14751 ( .A(n2985), .B(o[34]), .Z(n14866) );
  NANDN U14752 ( .A(n14150), .B(n14149), .Z(n14154) );
  NANDN U14753 ( .A(n14152), .B(n14151), .Z(n14153) );
  NAND U14754 ( .A(n14154), .B(n14153), .Z(n14868) );
  NANDN U14755 ( .A(n2987), .B(o[32]), .Z(n14489) );
  NANDN U14756 ( .A(n14156), .B(n14155), .Z(n14160) );
  NANDN U14757 ( .A(n14158), .B(n14157), .Z(n14159) );
  NAND U14758 ( .A(n14160), .B(n14159), .Z(n14491) );
  NANDN U14759 ( .A(n2989), .B(o[30]), .Z(n14854) );
  OR U14760 ( .A(n14162), .B(n14161), .Z(n14166) );
  OR U14761 ( .A(n14164), .B(n14163), .Z(n14165) );
  NAND U14762 ( .A(n14166), .B(n14165), .Z(n14856) );
  NANDN U14763 ( .A(n3021), .B(\stack[1][34] ), .Z(n14831) );
  OR U14764 ( .A(n14168), .B(n14167), .Z(n14172) );
  NANDN U14765 ( .A(n14170), .B(n14169), .Z(n14171) );
  NAND U14766 ( .A(n14172), .B(n14171), .Z(n14833) );
  NANDN U14767 ( .A(n14174), .B(n14173), .Z(n14178) );
  OR U14768 ( .A(n14176), .B(n14175), .Z(n14177) );
  AND U14769 ( .A(n14178), .B(n14177), .Z(n14814) );
  AND U14770 ( .A(\stack[1][37] ), .B(o[25]), .Z(n14502) );
  NANDN U14771 ( .A(n14180), .B(n14179), .Z(n14184) );
  OR U14772 ( .A(n14182), .B(n14181), .Z(n14183) );
  NAND U14773 ( .A(n14184), .B(n14183), .Z(n14503) );
  XNOR U14774 ( .A(n14502), .B(n14503), .Z(n14501) );
  ANDN U14775 ( .B(\stack[1][38] ), .A(n3018), .Z(n14820) );
  OR U14776 ( .A(n14186), .B(n14185), .Z(n14190) );
  OR U14777 ( .A(n14188), .B(n14187), .Z(n14189) );
  AND U14778 ( .A(n14190), .B(n14189), .Z(n14819) );
  AND U14779 ( .A(\stack[1][40] ), .B(o[22]), .Z(n14795) );
  AND U14780 ( .A(\stack[1][41] ), .B(o[21]), .Z(n14800) );
  NANDN U14781 ( .A(n3013), .B(\stack[1][43] ), .Z(n14779) );
  OR U14782 ( .A(n14192), .B(n14191), .Z(n14196) );
  NAND U14783 ( .A(n14194), .B(n14193), .Z(n14195) );
  AND U14784 ( .A(n14196), .B(n14195), .Z(n14759) );
  OR U14785 ( .A(n14198), .B(n14197), .Z(n14202) );
  OR U14786 ( .A(n14200), .B(n14199), .Z(n14201) );
  AND U14787 ( .A(n14202), .B(n14201), .Z(n14766) );
  NANDN U14788 ( .A(n3010), .B(\stack[1][46] ), .Z(n14767) );
  XOR U14789 ( .A(n14766), .B(n14767), .Z(n14765) );
  NANDN U14790 ( .A(n3009), .B(\stack[1][47] ), .Z(n14519) );
  NANDN U14791 ( .A(n14204), .B(n14203), .Z(n14208) );
  NANDN U14792 ( .A(n14206), .B(n14205), .Z(n14207) );
  AND U14793 ( .A(n14208), .B(n14207), .Z(n14525) );
  OR U14794 ( .A(n14210), .B(n14209), .Z(n14214) );
  OR U14795 ( .A(n14212), .B(n14211), .Z(n14213) );
  NAND U14796 ( .A(n14214), .B(n14213), .Z(n14747) );
  NANDN U14797 ( .A(n3006), .B(\stack[1][50] ), .Z(n14749) );
  NANDN U14798 ( .A(n15507), .B(o[11]), .Z(n14530) );
  OR U14799 ( .A(n14216), .B(n14215), .Z(n14220) );
  NANDN U14800 ( .A(n14218), .B(n14217), .Z(n14219) );
  AND U14801 ( .A(n14220), .B(n14219), .Z(n14533) );
  NANDN U14802 ( .A(n15468), .B(o[10]), .Z(n14722) );
  ANDN U14803 ( .B(\stack[1][53] ), .A(n3003), .Z(n14728) );
  NANDN U14804 ( .A(n14222), .B(n14221), .Z(n14226) );
  NAND U14805 ( .A(n14224), .B(n14223), .Z(n14225) );
  AND U14806 ( .A(n14226), .B(n14225), .Z(n14711) );
  ANDN U14807 ( .B(\stack[1][57] ), .A(n2999), .Z(n14687) );
  OR U14808 ( .A(n14228), .B(n14227), .Z(n14232) );
  NANDN U14809 ( .A(n14230), .B(n14229), .Z(n14231) );
  AND U14810 ( .A(n14232), .B(n14231), .Z(n14688) );
  AND U14811 ( .A(\stack[1][58] ), .B(o[4]), .Z(n14543) );
  AND U14812 ( .A(\stack[1][59] ), .B(o[3]), .Z(n14693) );
  NANDN U14813 ( .A(n14233), .B(n14679), .Z(n14234) );
  AND U14814 ( .A(n14235), .B(n14234), .Z(n14239) );
  OR U14815 ( .A(n14237), .B(n14236), .Z(n14238) );
  AND U14816 ( .A(n14239), .B(n14238), .Z(n14694) );
  NANDN U14817 ( .A(n2995), .B(\stack[1][62] ), .Z(n14555) );
  NOR U14818 ( .A(n14240), .B(n14555), .Z(n14678) );
  XNOR U14819 ( .A(n14678), .B(n14679), .Z(n14243) );
  NANDN U14820 ( .A(n2994), .B(\stack[1][62] ), .Z(n14241) );
  NAND U14821 ( .A(n14242), .B(n14241), .Z(n14681) );
  NAND U14822 ( .A(n14243), .B(n14681), .Z(n14677) );
  AND U14823 ( .A(\stack[1][60] ), .B(o[2]), .Z(n14676) );
  XNOR U14824 ( .A(n14677), .B(n14676), .Z(n14695) );
  XOR U14825 ( .A(n14694), .B(n14695), .Z(n14692) );
  XOR U14826 ( .A(n14693), .B(n14692), .Z(n14545) );
  OR U14827 ( .A(n14245), .B(n14244), .Z(n14249) );
  NANDN U14828 ( .A(n14247), .B(n14246), .Z(n14248) );
  AND U14829 ( .A(n14249), .B(n14248), .Z(n14544) );
  XOR U14830 ( .A(n14545), .B(n14544), .Z(n14542) );
  XOR U14831 ( .A(n14543), .B(n14542), .Z(n14689) );
  XNOR U14832 ( .A(n14688), .B(n14689), .Z(n14686) );
  OR U14833 ( .A(n14251), .B(n14250), .Z(n14255) );
  OR U14834 ( .A(n14253), .B(n14252), .Z(n14254) );
  NAND U14835 ( .A(n14255), .B(n14254), .Z(n14539) );
  IV U14836 ( .A(\stack[1][56] ), .Z(n15315) );
  ANDN U14837 ( .B(o[6]), .A(n15315), .Z(n14538) );
  XNOR U14838 ( .A(n14539), .B(n14538), .Z(n14537) );
  XNOR U14839 ( .A(n14536), .B(n14537), .Z(n14713) );
  ANDN U14840 ( .B(\stack[1][55] ), .A(n3001), .Z(n14712) );
  XOR U14841 ( .A(n14713), .B(n14712), .Z(n14710) );
  NANDN U14842 ( .A(n14257), .B(n14256), .Z(n14261) );
  OR U14843 ( .A(n14259), .B(n14258), .Z(n14260) );
  AND U14844 ( .A(n14261), .B(n14260), .Z(n14706) );
  XNOR U14845 ( .A(n14707), .B(n14706), .Z(n14705) );
  ANDN U14846 ( .B(\stack[1][54] ), .A(n3002), .Z(n14704) );
  XNOR U14847 ( .A(n14705), .B(n14704), .Z(n14730) );
  OR U14848 ( .A(n14263), .B(n14262), .Z(n14267) );
  NANDN U14849 ( .A(n14265), .B(n14264), .Z(n14266) );
  NAND U14850 ( .A(n14267), .B(n14266), .Z(n14731) );
  XNOR U14851 ( .A(n14730), .B(n14731), .Z(n14729) );
  XNOR U14852 ( .A(n14728), .B(n14729), .Z(n14725) );
  OR U14853 ( .A(n14269), .B(n14268), .Z(n14273) );
  OR U14854 ( .A(n14271), .B(n14270), .Z(n14272) );
  AND U14855 ( .A(n14273), .B(n14272), .Z(n14724) );
  XNOR U14856 ( .A(n14725), .B(n14724), .Z(n14723) );
  XNOR U14857 ( .A(n14722), .B(n14723), .Z(n14532) );
  XOR U14858 ( .A(n14533), .B(n14532), .Z(n14531) );
  XNOR U14859 ( .A(n14530), .B(n14531), .Z(n14748) );
  XNOR U14860 ( .A(n14749), .B(n14748), .Z(n14746) );
  XNOR U14861 ( .A(n14747), .B(n14746), .Z(n14527) );
  ANDN U14862 ( .B(\stack[1][49] ), .A(n3007), .Z(n14526) );
  XOR U14863 ( .A(n14527), .B(n14526), .Z(n14524) );
  NANDN U14864 ( .A(n14275), .B(n14274), .Z(n14279) );
  OR U14865 ( .A(n14277), .B(n14276), .Z(n14278) );
  AND U14866 ( .A(n14279), .B(n14278), .Z(n14742) );
  XNOR U14867 ( .A(n14743), .B(n14742), .Z(n14741) );
  ANDN U14868 ( .B(o[14]), .A(n15623), .Z(n14740) );
  XOR U14869 ( .A(n14741), .B(n14740), .Z(n14521) );
  OR U14870 ( .A(n14281), .B(n14280), .Z(n14285) );
  NANDN U14871 ( .A(n14283), .B(n14282), .Z(n14284) );
  AND U14872 ( .A(n14285), .B(n14284), .Z(n14520) );
  XNOR U14873 ( .A(n14521), .B(n14520), .Z(n14518) );
  XOR U14874 ( .A(n14519), .B(n14518), .Z(n14764) );
  XNOR U14875 ( .A(n14765), .B(n14764), .Z(n14761) );
  ANDN U14876 ( .B(o[17]), .A(n15740), .Z(n14760) );
  XOR U14877 ( .A(n14761), .B(n14760), .Z(n14758) );
  NANDN U14878 ( .A(n14287), .B(n14286), .Z(n14291) );
  OR U14879 ( .A(n14289), .B(n14288), .Z(n14290) );
  AND U14880 ( .A(n14291), .B(n14290), .Z(n14784) );
  XNOR U14881 ( .A(n14785), .B(n14784), .Z(n14783) );
  NANDN U14882 ( .A(n3012), .B(\stack[1][44] ), .Z(n14782) );
  XOR U14883 ( .A(n14783), .B(n14782), .Z(n14778) );
  XOR U14884 ( .A(n14779), .B(n14778), .Z(n14777) );
  OR U14885 ( .A(n14293), .B(n14292), .Z(n14297) );
  NANDN U14886 ( .A(n14295), .B(n14294), .Z(n14296) );
  AND U14887 ( .A(n14297), .B(n14296), .Z(n14776) );
  XNOR U14888 ( .A(n14777), .B(n14776), .Z(n14514) );
  OR U14889 ( .A(n14299), .B(n14298), .Z(n14303) );
  NANDN U14890 ( .A(n14301), .B(n14300), .Z(n14302) );
  AND U14891 ( .A(n14303), .B(n14302), .Z(n14515) );
  AND U14892 ( .A(\stack[1][42] ), .B(o[20]), .Z(n14512) );
  XNOR U14893 ( .A(n14513), .B(n14512), .Z(n14802) );
  OR U14894 ( .A(n14305), .B(n14304), .Z(n14309) );
  NANDN U14895 ( .A(n14307), .B(n14306), .Z(n14308) );
  NAND U14896 ( .A(n14309), .B(n14308), .Z(n14803) );
  XNOR U14897 ( .A(n14802), .B(n14803), .Z(n14801) );
  XNOR U14898 ( .A(n14800), .B(n14801), .Z(n14797) );
  OR U14899 ( .A(n14311), .B(n14310), .Z(n14315) );
  OR U14900 ( .A(n14313), .B(n14312), .Z(n14314) );
  AND U14901 ( .A(n14315), .B(n14314), .Z(n14796) );
  XNOR U14902 ( .A(n14797), .B(n14796), .Z(n14794) );
  NANDN U14903 ( .A(n3017), .B(\stack[1][39] ), .Z(n14509) );
  XOR U14904 ( .A(n14508), .B(n14509), .Z(n14507) );
  OR U14905 ( .A(n14317), .B(n14316), .Z(n14321) );
  NANDN U14906 ( .A(n14319), .B(n14318), .Z(n14320) );
  NAND U14907 ( .A(n14321), .B(n14320), .Z(n14506) );
  XOR U14908 ( .A(n14507), .B(n14506), .Z(n14818) );
  XOR U14909 ( .A(n14819), .B(n14818), .Z(n14821) );
  XOR U14910 ( .A(n14820), .B(n14821), .Z(n14500) );
  XOR U14911 ( .A(n14501), .B(n14500), .Z(n14815) );
  XOR U14912 ( .A(n14814), .B(n14815), .Z(n14813) );
  AND U14913 ( .A(\stack[1][36] ), .B(o[26]), .Z(n14812) );
  XOR U14914 ( .A(n14813), .B(n14812), .Z(n14839) );
  OR U14915 ( .A(n14323), .B(n14322), .Z(n14327) );
  OR U14916 ( .A(n14325), .B(n14324), .Z(n14326) );
  AND U14917 ( .A(n14327), .B(n14326), .Z(n14836) );
  NANDN U14918 ( .A(n2992), .B(o[27]), .Z(n14837) );
  XOR U14919 ( .A(n14836), .B(n14837), .Z(n14838) );
  XOR U14920 ( .A(n14839), .B(n14838), .Z(n14832) );
  XNOR U14921 ( .A(n14833), .B(n14832), .Z(n14830) );
  XNOR U14922 ( .A(n14831), .B(n14830), .Z(n14494) );
  OR U14923 ( .A(n14329), .B(n14328), .Z(n14333) );
  NANDN U14924 ( .A(n14331), .B(n14330), .Z(n14332) );
  AND U14925 ( .A(n14333), .B(n14332), .Z(n14497) );
  NANDN U14926 ( .A(n2990), .B(o[29]), .Z(n14496) );
  XOR U14927 ( .A(n14497), .B(n14496), .Z(n14495) );
  XNOR U14928 ( .A(n14494), .B(n14495), .Z(n14855) );
  XNOR U14929 ( .A(n14856), .B(n14855), .Z(n14853) );
  XNOR U14930 ( .A(n14854), .B(n14853), .Z(n14848) );
  AND U14931 ( .A(o[31]), .B(\stack[1][31] ), .Z(n16283) );
  OR U14932 ( .A(n14335), .B(n14334), .Z(n14339) );
  OR U14933 ( .A(n14337), .B(n14336), .Z(n14338) );
  NAND U14934 ( .A(n14339), .B(n14338), .Z(n14850) );
  XNOR U14935 ( .A(n16283), .B(n14850), .Z(n14849) );
  XNOR U14936 ( .A(n14848), .B(n14849), .Z(n14490) );
  XNOR U14937 ( .A(n14491), .B(n14490), .Z(n14488) );
  XNOR U14938 ( .A(n14489), .B(n14488), .Z(n14871) );
  NANDN U14939 ( .A(n2986), .B(o[33]), .Z(n14873) );
  OR U14940 ( .A(n14341), .B(n14340), .Z(n14345) );
  OR U14941 ( .A(n14343), .B(n14342), .Z(n14344) );
  NAND U14942 ( .A(n14345), .B(n14344), .Z(n14874) );
  XOR U14943 ( .A(n14873), .B(n14874), .Z(n14872) );
  XNOR U14944 ( .A(n14871), .B(n14872), .Z(n14867) );
  XNOR U14945 ( .A(n14868), .B(n14867), .Z(n14865) );
  XNOR U14946 ( .A(n14866), .B(n14865), .Z(n14482) );
  NANDN U14947 ( .A(n2984), .B(o[35]), .Z(n14484) );
  OR U14948 ( .A(n14347), .B(n14346), .Z(n14351) );
  OR U14949 ( .A(n14349), .B(n14348), .Z(n14350) );
  NAND U14950 ( .A(n14351), .B(n14350), .Z(n14485) );
  XOR U14951 ( .A(n14484), .B(n14485), .Z(n14483) );
  XNOR U14952 ( .A(n14482), .B(n14483), .Z(n14478) );
  XNOR U14953 ( .A(n14479), .B(n14478), .Z(n14476) );
  XNOR U14954 ( .A(n14477), .B(n14476), .Z(n14889) );
  NANDN U14955 ( .A(n2982), .B(o[37]), .Z(n14891) );
  OR U14956 ( .A(n14353), .B(n14352), .Z(n14357) );
  OR U14957 ( .A(n14355), .B(n14354), .Z(n14356) );
  NAND U14958 ( .A(n14357), .B(n14356), .Z(n14892) );
  XOR U14959 ( .A(n14891), .B(n14892), .Z(n14890) );
  XNOR U14960 ( .A(n14889), .B(n14890), .Z(n14885) );
  XNOR U14961 ( .A(n14886), .B(n14885), .Z(n14883) );
  XNOR U14962 ( .A(n14884), .B(n14883), .Z(n14470) );
  NANDN U14963 ( .A(n2980), .B(o[39]), .Z(n14472) );
  OR U14964 ( .A(n14359), .B(n14358), .Z(n14363) );
  OR U14965 ( .A(n14361), .B(n14360), .Z(n14362) );
  NAND U14966 ( .A(n14363), .B(n14362), .Z(n14473) );
  XOR U14967 ( .A(n14472), .B(n14473), .Z(n14471) );
  XNOR U14968 ( .A(n14470), .B(n14471), .Z(n14907) );
  XNOR U14969 ( .A(n14908), .B(n14907), .Z(n14910) );
  XNOR U14970 ( .A(n14909), .B(n14910), .Z(n14901) );
  NANDN U14971 ( .A(n2978), .B(o[41]), .Z(n14903) );
  OR U14972 ( .A(n14365), .B(n14364), .Z(n14369) );
  OR U14973 ( .A(n14367), .B(n14366), .Z(n14368) );
  NAND U14974 ( .A(n14369), .B(n14368), .Z(n14904) );
  XOR U14975 ( .A(n14903), .B(n14904), .Z(n14902) );
  XNOR U14976 ( .A(n14901), .B(n14902), .Z(n14927) );
  XNOR U14977 ( .A(n14928), .B(n14927), .Z(n14925) );
  XNOR U14978 ( .A(n14926), .B(n14925), .Z(n14464) );
  NANDN U14979 ( .A(n16746), .B(o[43]), .Z(n14466) );
  OR U14980 ( .A(n14371), .B(n14370), .Z(n14375) );
  OR U14981 ( .A(n14373), .B(n14372), .Z(n14374) );
  NAND U14982 ( .A(n14375), .B(n14374), .Z(n14467) );
  XOR U14983 ( .A(n14466), .B(n14467), .Z(n14465) );
  XNOR U14984 ( .A(n14464), .B(n14465), .Z(n14921) );
  XNOR U14985 ( .A(n14922), .B(n14921), .Z(n14919) );
  XNOR U14986 ( .A(n14920), .B(n14919), .Z(n14458) );
  NANDN U14987 ( .A(n16826), .B(o[45]), .Z(n14460) );
  OR U14988 ( .A(n14377), .B(n14376), .Z(n14381) );
  OR U14989 ( .A(n14379), .B(n14378), .Z(n14380) );
  NAND U14990 ( .A(n14381), .B(n14380), .Z(n14461) );
  XOR U14991 ( .A(n14460), .B(n14461), .Z(n14459) );
  XNOR U14992 ( .A(n14458), .B(n14459), .Z(n14945) );
  XNOR U14993 ( .A(n14946), .B(n14945), .Z(n14943) );
  XNOR U14994 ( .A(n14944), .B(n14943), .Z(n14937) );
  NANDN U14995 ( .A(n2976), .B(o[47]), .Z(n14939) );
  OR U14996 ( .A(n14383), .B(n14382), .Z(n14387) );
  OR U14997 ( .A(n14385), .B(n14384), .Z(n14386) );
  NAND U14998 ( .A(n14387), .B(n14386), .Z(n14940) );
  XOR U14999 ( .A(n14939), .B(n14940), .Z(n14938) );
  XNOR U15000 ( .A(n14937), .B(n14938), .Z(n14963) );
  XNOR U15001 ( .A(n14964), .B(n14963), .Z(n14961) );
  XNOR U15002 ( .A(n14962), .B(n14961), .Z(n14955) );
  NANDN U15003 ( .A(n2974), .B(o[49]), .Z(n14957) );
  OR U15004 ( .A(n14389), .B(n14388), .Z(n14393) );
  OR U15005 ( .A(n14391), .B(n14390), .Z(n14392) );
  NAND U15006 ( .A(n14393), .B(n14392), .Z(n14958) );
  XOR U15007 ( .A(n14957), .B(n14958), .Z(n14956) );
  XNOR U15008 ( .A(n14955), .B(n14956), .Z(n14454) );
  XNOR U15009 ( .A(n14455), .B(n14454), .Z(n14452) );
  XNOR U15010 ( .A(n14453), .B(n14452), .Z(n14979) );
  NANDN U15011 ( .A(n2972), .B(o[51]), .Z(n14981) );
  OR U15012 ( .A(n14395), .B(n14394), .Z(n14399) );
  OR U15013 ( .A(n14397), .B(n14396), .Z(n14398) );
  NAND U15014 ( .A(n14399), .B(n14398), .Z(n14982) );
  XOR U15015 ( .A(n14981), .B(n14982), .Z(n14980) );
  XNOR U15016 ( .A(n14979), .B(n14980), .Z(n14448) );
  XNOR U15017 ( .A(n14449), .B(n14448), .Z(n14446) );
  XNOR U15018 ( .A(n14447), .B(n14446), .Z(n14973) );
  NANDN U15019 ( .A(n17145), .B(o[53]), .Z(n14975) );
  OR U15020 ( .A(n14401), .B(n14400), .Z(n14405) );
  OR U15021 ( .A(n14403), .B(n14402), .Z(n14404) );
  NAND U15022 ( .A(n14405), .B(n14404), .Z(n14976) );
  XOR U15023 ( .A(n14975), .B(n14976), .Z(n14974) );
  XNOR U15024 ( .A(n14973), .B(n14974), .Z(n14442) );
  XNOR U15025 ( .A(n14443), .B(n14442), .Z(n14440) );
  XNOR U15026 ( .A(n14441), .B(n14440), .Z(n15000) );
  NANDN U15027 ( .A(n17219), .B(o[55]), .Z(n14998) );
  OR U15028 ( .A(n14407), .B(n14406), .Z(n14411) );
  OR U15029 ( .A(n14409), .B(n14408), .Z(n14410) );
  NAND U15030 ( .A(n14411), .B(n14410), .Z(n14997) );
  XOR U15031 ( .A(n14998), .B(n14997), .Z(n14999) );
  XNOR U15032 ( .A(n15000), .B(n14999), .Z(n14993) );
  XNOR U15033 ( .A(n14994), .B(n14993), .Z(n14991) );
  XNOR U15034 ( .A(n14992), .B(n14991), .Z(n15015) );
  NANDN U15035 ( .A(n17296), .B(o[57]), .Z(n15017) );
  OR U15036 ( .A(n14413), .B(n14412), .Z(n14417) );
  OR U15037 ( .A(n14415), .B(n14414), .Z(n14416) );
  NAND U15038 ( .A(n14417), .B(n14416), .Z(n15018) );
  XOR U15039 ( .A(n15017), .B(n15018), .Z(n15016) );
  XNOR U15040 ( .A(n15015), .B(n15016), .Z(n14436) );
  XNOR U15041 ( .A(n14437), .B(n14436), .Z(n14434) );
  XNOR U15042 ( .A(n14435), .B(n14434), .Z(n15009) );
  NANDN U15043 ( .A(n17375), .B(o[59]), .Z(n15011) );
  OR U15044 ( .A(n14419), .B(n14418), .Z(n14423) );
  OR U15045 ( .A(n14421), .B(n14420), .Z(n14422) );
  NAND U15046 ( .A(n14423), .B(n14422), .Z(n15012) );
  XOR U15047 ( .A(n15011), .B(n15012), .Z(n15010) );
  XNOR U15048 ( .A(n15009), .B(n15010), .Z(n15033) );
  XNOR U15049 ( .A(n15034), .B(n15033), .Z(n15036) );
  XNOR U15050 ( .A(n15035), .B(n15036), .Z(n15027) );
  AND U15051 ( .A(o[61]), .B(\stack[1][1] ), .Z(n15030) );
  OR U15052 ( .A(n14425), .B(n14424), .Z(n14429) );
  OR U15053 ( .A(n14427), .B(n14426), .Z(n14428) );
  NAND U15054 ( .A(n14429), .B(n14428), .Z(n15029) );
  XNOR U15055 ( .A(n15030), .B(n15029), .Z(n15028) );
  XOR U15056 ( .A(n15027), .B(n15028), .Z(n14431) );
  XNOR U15057 ( .A(n14430), .B(n14431), .Z(n15086) );
  AND U15058 ( .A(o[62]), .B(\stack[1][0] ), .Z(n15087) );
  OR U15059 ( .A(n15086), .B(n15087), .Z(n14433) );
  OR U15060 ( .A(n14431), .B(n14430), .Z(n14432) );
  AND U15061 ( .A(n14433), .B(n14432), .Z(n15044) );
  OR U15062 ( .A(n14435), .B(n14434), .Z(n14439) );
  OR U15063 ( .A(n14437), .B(n14436), .Z(n14438) );
  AND U15064 ( .A(n14439), .B(n14438), .Z(n15026) );
  OR U15065 ( .A(n14441), .B(n14440), .Z(n14445) );
  OR U15066 ( .A(n14443), .B(n14442), .Z(n14444) );
  AND U15067 ( .A(n14445), .B(n14444), .Z(n15008) );
  OR U15068 ( .A(n14447), .B(n14446), .Z(n14451) );
  OR U15069 ( .A(n14449), .B(n14448), .Z(n14450) );
  AND U15070 ( .A(n14451), .B(n14450), .Z(n14990) );
  OR U15071 ( .A(n14453), .B(n14452), .Z(n14457) );
  OR U15072 ( .A(n14455), .B(n14454), .Z(n14456) );
  AND U15073 ( .A(n14457), .B(n14456), .Z(n14972) );
  NANDN U15074 ( .A(n14459), .B(n14458), .Z(n14463) );
  NANDN U15075 ( .A(n14461), .B(n14460), .Z(n14462) );
  AND U15076 ( .A(n14463), .B(n14462), .Z(n14954) );
  NANDN U15077 ( .A(n14465), .B(n14464), .Z(n14469) );
  NANDN U15078 ( .A(n14467), .B(n14466), .Z(n14468) );
  AND U15079 ( .A(n14469), .B(n14468), .Z(n14936) );
  NANDN U15080 ( .A(n14471), .B(n14470), .Z(n14475) );
  NANDN U15081 ( .A(n14473), .B(n14472), .Z(n14474) );
  AND U15082 ( .A(n14475), .B(n14474), .Z(n14918) );
  OR U15083 ( .A(n14477), .B(n14476), .Z(n14481) );
  OR U15084 ( .A(n14479), .B(n14478), .Z(n14480) );
  AND U15085 ( .A(n14481), .B(n14480), .Z(n14900) );
  NANDN U15086 ( .A(n14483), .B(n14482), .Z(n14487) );
  NANDN U15087 ( .A(n14485), .B(n14484), .Z(n14486) );
  AND U15088 ( .A(n14487), .B(n14486), .Z(n14882) );
  OR U15089 ( .A(n14489), .B(n14488), .Z(n14493) );
  OR U15090 ( .A(n14491), .B(n14490), .Z(n14492) );
  AND U15091 ( .A(n14493), .B(n14492), .Z(n14864) );
  NANDN U15092 ( .A(n14495), .B(n14494), .Z(n14499) );
  NANDN U15093 ( .A(n14497), .B(n14496), .Z(n14498) );
  AND U15094 ( .A(n14499), .B(n14498), .Z(n14847) );
  OR U15095 ( .A(n14501), .B(n14500), .Z(n14505) );
  OR U15096 ( .A(n14503), .B(n14502), .Z(n14504) );
  AND U15097 ( .A(n14505), .B(n14504), .Z(n14829) );
  OR U15098 ( .A(n14507), .B(n14506), .Z(n14511) );
  NANDN U15099 ( .A(n14509), .B(n14508), .Z(n14510) );
  AND U15100 ( .A(n14511), .B(n14510), .Z(n14811) );
  NANDN U15101 ( .A(n14513), .B(n14512), .Z(n14517) );
  OR U15102 ( .A(n14515), .B(n14514), .Z(n14516) );
  AND U15103 ( .A(n14517), .B(n14516), .Z(n14793) );
  OR U15104 ( .A(n14519), .B(n14518), .Z(n14523) );
  OR U15105 ( .A(n14521), .B(n14520), .Z(n14522) );
  AND U15106 ( .A(n14523), .B(n14522), .Z(n14775) );
  OR U15107 ( .A(n14525), .B(n14524), .Z(n14529) );
  NANDN U15108 ( .A(n14527), .B(n14526), .Z(n14528) );
  AND U15109 ( .A(n14529), .B(n14528), .Z(n14757) );
  NANDN U15110 ( .A(n14531), .B(n14530), .Z(n14535) );
  NANDN U15111 ( .A(n14533), .B(n14532), .Z(n14534) );
  AND U15112 ( .A(n14535), .B(n14534), .Z(n14739) );
  NAND U15113 ( .A(n14537), .B(n14536), .Z(n14541) );
  NANDN U15114 ( .A(n14539), .B(n14538), .Z(n14540) );
  AND U15115 ( .A(n14541), .B(n14540), .Z(n14721) );
  NANDN U15116 ( .A(n14543), .B(n14542), .Z(n14547) );
  OR U15117 ( .A(n14545), .B(n14544), .Z(n14546) );
  AND U15118 ( .A(n14547), .B(n14546), .Z(n14703) );
  XOR U15119 ( .A(\stack[1][63] ), .B(n14678), .Z(n14549) );
  NANDN U15120 ( .A(o[0]), .B(\stack[1][63] ), .Z(n14548) );
  NAND U15121 ( .A(n14549), .B(n14548), .Z(n14579) );
  ANDN U15122 ( .B(o[59]), .A(n2971), .Z(n14561) );
  ANDN U15123 ( .B(o[61]), .A(n2970), .Z(n14551) );
  NANDN U15124 ( .A(n2969), .B(o[62]), .Z(n14550) );
  XNOR U15125 ( .A(n14551), .B(n14550), .Z(n14559) );
  ANDN U15126 ( .B(o[63]), .A(n2968), .Z(n14557) );
  ANDN U15127 ( .B(o[56]), .A(n17219), .Z(n14553) );
  NANDN U15128 ( .A(n17256), .B(o[57]), .Z(n14552) );
  XNOR U15129 ( .A(n14553), .B(n14552), .Z(n14554) );
  XOR U15130 ( .A(n14555), .B(n14554), .Z(n14556) );
  XNOR U15131 ( .A(n14557), .B(n14556), .Z(n14558) );
  XNOR U15132 ( .A(n14559), .B(n14558), .Z(n14560) );
  XNOR U15133 ( .A(n14561), .B(n14560), .Z(n14577) );
  ANDN U15134 ( .B(o[50]), .A(n2974), .Z(n14563) );
  NANDN U15135 ( .A(n17296), .B(o[58]), .Z(n14562) );
  XNOR U15136 ( .A(n14563), .B(n14562), .Z(n14567) );
  ANDN U15137 ( .B(o[47]), .A(n2977), .Z(n14565) );
  NANDN U15138 ( .A(n2975), .B(o[49]), .Z(n14564) );
  XNOR U15139 ( .A(n14565), .B(n14564), .Z(n14566) );
  XOR U15140 ( .A(n14567), .B(n14566), .Z(n14575) );
  ANDN U15141 ( .B(o[45]), .A(n16786), .Z(n14569) );
  NANDN U15142 ( .A(n2973), .B(o[51]), .Z(n14568) );
  XNOR U15143 ( .A(n14569), .B(n14568), .Z(n14573) );
  ANDN U15144 ( .B(o[33]), .A(n2987), .Z(n14571) );
  NANDN U15145 ( .A(n2983), .B(o[37]), .Z(n14570) );
  XNOR U15146 ( .A(n14571), .B(n14570), .Z(n14572) );
  XNOR U15147 ( .A(n14573), .B(n14572), .Z(n14574) );
  XNOR U15148 ( .A(n14575), .B(n14574), .Z(n14576) );
  XOR U15149 ( .A(n14577), .B(n14576), .Z(n14578) );
  XNOR U15150 ( .A(n14579), .B(n14578), .Z(n14643) );
  ANDN U15151 ( .B(o[23]), .A(n15935), .Z(n14581) );
  NANDN U15152 ( .A(n3016), .B(\stack[1][41] ), .Z(n14580) );
  XNOR U15153 ( .A(n14581), .B(n14580), .Z(n14585) );
  ANDN U15154 ( .B(\stack[1][49] ), .A(n3008), .Z(n14583) );
  NANDN U15155 ( .A(n2997), .B(\stack[1][60] ), .Z(n14582) );
  XNOR U15156 ( .A(n14583), .B(n14582), .Z(n14584) );
  XOR U15157 ( .A(n14585), .B(n14584), .Z(n14593) );
  ANDN U15158 ( .B(o[29]), .A(n2991), .Z(n14587) );
  NANDN U15159 ( .A(n3020), .B(\stack[1][37] ), .Z(n14586) );
  XNOR U15160 ( .A(n14587), .B(n14586), .Z(n14591) );
  ANDN U15161 ( .B(\stack[1][38] ), .A(n3019), .Z(n14589) );
  NANDN U15162 ( .A(n3015), .B(\stack[1][42] ), .Z(n14588) );
  XNOR U15163 ( .A(n14589), .B(n14588), .Z(n14590) );
  XNOR U15164 ( .A(n14591), .B(n14590), .Z(n14592) );
  XNOR U15165 ( .A(n14593), .B(n14592), .Z(n14609) );
  ANDN U15166 ( .B(\stack[1][57] ), .A(n3000), .Z(n14595) );
  NANDN U15167 ( .A(n2998), .B(\stack[1][59] ), .Z(n14594) );
  XNOR U15168 ( .A(n14595), .B(n14594), .Z(n14599) );
  ANDN U15169 ( .B(\stack[1][55] ), .A(n3002), .Z(n14597) );
  NANDN U15170 ( .A(n3001), .B(\stack[1][56] ), .Z(n14596) );
  XNOR U15171 ( .A(n14597), .B(n14596), .Z(n14598) );
  XOR U15172 ( .A(n14599), .B(n14598), .Z(n14607) );
  ANDN U15173 ( .B(\stack[1][53] ), .A(n3004), .Z(n14601) );
  NANDN U15174 ( .A(n2999), .B(\stack[1][58] ), .Z(n14600) );
  XNOR U15175 ( .A(n14601), .B(n14600), .Z(n14605) );
  ANDN U15176 ( .B(\stack[1][54] ), .A(n3003), .Z(n14603) );
  NANDN U15177 ( .A(n2996), .B(\stack[1][61] ), .Z(n14602) );
  XNOR U15178 ( .A(n14603), .B(n14602), .Z(n14604) );
  XNOR U15179 ( .A(n14605), .B(n14604), .Z(n14606) );
  XNOR U15180 ( .A(n14607), .B(n14606), .Z(n14608) );
  XOR U15181 ( .A(n14609), .B(n14608), .Z(n14641) );
  ANDN U15182 ( .B(o[48]), .A(n2976), .Z(n14611) );
  NANDN U15183 ( .A(n2972), .B(o[52]), .Z(n14610) );
  XNOR U15184 ( .A(n14611), .B(n14610), .Z(n14615) );
  ANDN U15185 ( .B(o[42]), .A(n2978), .Z(n14613) );
  NANDN U15186 ( .A(n16826), .B(o[46]), .Z(n14612) );
  XNOR U15187 ( .A(n14613), .B(n14612), .Z(n14614) );
  XOR U15188 ( .A(n14615), .B(n14614), .Z(n14623) );
  ANDN U15189 ( .B(o[54]), .A(n17145), .Z(n14617) );
  NANDN U15190 ( .A(n17375), .B(o[60]), .Z(n14616) );
  XNOR U15191 ( .A(n14617), .B(n14616), .Z(n14621) );
  ANDN U15192 ( .B(o[53]), .A(n17101), .Z(n14619) );
  NANDN U15193 ( .A(n17179), .B(o[55]), .Z(n14618) );
  XNOR U15194 ( .A(n14619), .B(n14618), .Z(n14620) );
  XNOR U15195 ( .A(n14621), .B(n14620), .Z(n14622) );
  XNOR U15196 ( .A(n14623), .B(n14622), .Z(n14639) );
  ANDN U15197 ( .B(o[38]), .A(n2982), .Z(n14625) );
  NANDN U15198 ( .A(n2980), .B(o[40]), .Z(n14624) );
  XNOR U15199 ( .A(n14625), .B(n14624), .Z(n14629) );
  ANDN U15200 ( .B(o[31]), .A(n2989), .Z(n14627) );
  NANDN U15201 ( .A(n2984), .B(o[36]), .Z(n14626) );
  XNOR U15202 ( .A(n14627), .B(n14626), .Z(n14628) );
  XOR U15203 ( .A(n14629), .B(n14628), .Z(n14637) );
  ANDN U15204 ( .B(o[43]), .A(n16712), .Z(n14631) );
  NANDN U15205 ( .A(n16746), .B(o[44]), .Z(n14630) );
  XNOR U15206 ( .A(n14631), .B(n14630), .Z(n14635) );
  ANDN U15207 ( .B(o[39]), .A(n2981), .Z(n14633) );
  NANDN U15208 ( .A(n2979), .B(o[41]), .Z(n14632) );
  XNOR U15209 ( .A(n14633), .B(n14632), .Z(n14634) );
  XNOR U15210 ( .A(n14635), .B(n14634), .Z(n14636) );
  XNOR U15211 ( .A(n14637), .B(n14636), .Z(n14638) );
  XNOR U15212 ( .A(n14639), .B(n14638), .Z(n14640) );
  XNOR U15213 ( .A(n14641), .B(n14640), .Z(n14642) );
  XOR U15214 ( .A(n14643), .B(n14642), .Z(n14675) );
  ANDN U15215 ( .B(o[32]), .A(n2988), .Z(n14645) );
  NANDN U15216 ( .A(n2985), .B(o[35]), .Z(n14644) );
  XNOR U15217 ( .A(n14645), .B(n14644), .Z(n14649) );
  ANDN U15218 ( .B(o[30]), .A(n2990), .Z(n14647) );
  NANDN U15219 ( .A(n2986), .B(o[34]), .Z(n14646) );
  XNOR U15220 ( .A(n14647), .B(n14646), .Z(n14648) );
  XOR U15221 ( .A(n14649), .B(n14648), .Z(n14657) );
  ANDN U15222 ( .B(o[28]), .A(n2992), .Z(n14651) );
  NANDN U15223 ( .A(n3018), .B(\stack[1][39] ), .Z(n14650) );
  XNOR U15224 ( .A(n14651), .B(n14650), .Z(n14655) );
  ANDN U15225 ( .B(o[27]), .A(n2993), .Z(n14653) );
  NANDN U15226 ( .A(n3011), .B(\stack[1][46] ), .Z(n14652) );
  XNOR U15227 ( .A(n14653), .B(n14652), .Z(n14654) );
  XNOR U15228 ( .A(n14655), .B(n14654), .Z(n14656) );
  XNOR U15229 ( .A(n14657), .B(n14656), .Z(n14673) );
  ANDN U15230 ( .B(o[20]), .A(n15818), .Z(n14659) );
  NANDN U15231 ( .A(n3012), .B(\stack[1][45] ), .Z(n14658) );
  XNOR U15232 ( .A(n14659), .B(n14658), .Z(n14663) );
  ANDN U15233 ( .B(o[19]), .A(n15779), .Z(n14661) );
  NANDN U15234 ( .A(n3006), .B(\stack[1][51] ), .Z(n14660) );
  XNOR U15235 ( .A(n14661), .B(n14660), .Z(n14662) );
  XOR U15236 ( .A(n14663), .B(n14662), .Z(n14671) );
  ANDN U15237 ( .B(o[16]), .A(n15662), .Z(n14665) );
  NANDN U15238 ( .A(n3005), .B(\stack[1][52] ), .Z(n14664) );
  XNOR U15239 ( .A(n14665), .B(n14664), .Z(n14669) );
  ANDN U15240 ( .B(o[15]), .A(n15623), .Z(n14667) );
  NANDN U15241 ( .A(n3007), .B(\stack[1][50] ), .Z(n14666) );
  XNOR U15242 ( .A(n14667), .B(n14666), .Z(n14668) );
  XNOR U15243 ( .A(n14669), .B(n14668), .Z(n14670) );
  XNOR U15244 ( .A(n14671), .B(n14670), .Z(n14672) );
  XNOR U15245 ( .A(n14673), .B(n14672), .Z(n14674) );
  XNOR U15246 ( .A(n14675), .B(n14674), .Z(n14685) );
  OR U15247 ( .A(n14677), .B(n14676), .Z(n14683) );
  NANDN U15248 ( .A(n14679), .B(n14678), .Z(n14680) );
  AND U15249 ( .A(n14681), .B(n14680), .Z(n14682) );
  NAND U15250 ( .A(n14683), .B(n14682), .Z(n14684) );
  XNOR U15251 ( .A(n14685), .B(n14684), .Z(n14701) );
  OR U15252 ( .A(n14687), .B(n14686), .Z(n14691) );
  OR U15253 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15254 ( .A(n14691), .B(n14690), .Z(n14699) );
  NANDN U15255 ( .A(n14693), .B(n14692), .Z(n14697) );
  OR U15256 ( .A(n14695), .B(n14694), .Z(n14696) );
  NAND U15257 ( .A(n14697), .B(n14696), .Z(n14698) );
  XNOR U15258 ( .A(n14699), .B(n14698), .Z(n14700) );
  XNOR U15259 ( .A(n14701), .B(n14700), .Z(n14702) );
  XNOR U15260 ( .A(n14703), .B(n14702), .Z(n14719) );
  NANDN U15261 ( .A(n14705), .B(n14704), .Z(n14709) );
  OR U15262 ( .A(n14707), .B(n14706), .Z(n14708) );
  AND U15263 ( .A(n14709), .B(n14708), .Z(n14717) );
  OR U15264 ( .A(n14711), .B(n14710), .Z(n14715) );
  NANDN U15265 ( .A(n14713), .B(n14712), .Z(n14714) );
  NAND U15266 ( .A(n14715), .B(n14714), .Z(n14716) );
  XNOR U15267 ( .A(n14717), .B(n14716), .Z(n14718) );
  XNOR U15268 ( .A(n14719), .B(n14718), .Z(n14720) );
  XNOR U15269 ( .A(n14721), .B(n14720), .Z(n14737) );
  NANDN U15270 ( .A(n14723), .B(n14722), .Z(n14727) );
  OR U15271 ( .A(n14725), .B(n14724), .Z(n14726) );
  AND U15272 ( .A(n14727), .B(n14726), .Z(n14735) );
  OR U15273 ( .A(n14729), .B(n14728), .Z(n14733) );
  OR U15274 ( .A(n14731), .B(n14730), .Z(n14732) );
  NAND U15275 ( .A(n14733), .B(n14732), .Z(n14734) );
  XNOR U15276 ( .A(n14735), .B(n14734), .Z(n14736) );
  XNOR U15277 ( .A(n14737), .B(n14736), .Z(n14738) );
  XNOR U15278 ( .A(n14739), .B(n14738), .Z(n14755) );
  NANDN U15279 ( .A(n14741), .B(n14740), .Z(n14745) );
  OR U15280 ( .A(n14743), .B(n14742), .Z(n14744) );
  AND U15281 ( .A(n14745), .B(n14744), .Z(n14753) );
  OR U15282 ( .A(n14747), .B(n14746), .Z(n14751) );
  OR U15283 ( .A(n14749), .B(n14748), .Z(n14750) );
  NAND U15284 ( .A(n14751), .B(n14750), .Z(n14752) );
  XNOR U15285 ( .A(n14753), .B(n14752), .Z(n14754) );
  XNOR U15286 ( .A(n14755), .B(n14754), .Z(n14756) );
  XNOR U15287 ( .A(n14757), .B(n14756), .Z(n14773) );
  OR U15288 ( .A(n14759), .B(n14758), .Z(n14763) );
  NANDN U15289 ( .A(n14761), .B(n14760), .Z(n14762) );
  AND U15290 ( .A(n14763), .B(n14762), .Z(n14771) );
  NAND U15291 ( .A(n14765), .B(n14764), .Z(n14769) );
  OR U15292 ( .A(n14767), .B(n14766), .Z(n14768) );
  NAND U15293 ( .A(n14769), .B(n14768), .Z(n14770) );
  XNOR U15294 ( .A(n14771), .B(n14770), .Z(n14772) );
  XNOR U15295 ( .A(n14773), .B(n14772), .Z(n14774) );
  XNOR U15296 ( .A(n14775), .B(n14774), .Z(n14791) );
  OR U15297 ( .A(n14777), .B(n14776), .Z(n14781) );
  NANDN U15298 ( .A(n14779), .B(n14778), .Z(n14780) );
  AND U15299 ( .A(n14781), .B(n14780), .Z(n14789) );
  OR U15300 ( .A(n14783), .B(n14782), .Z(n14787) );
  OR U15301 ( .A(n14785), .B(n14784), .Z(n14786) );
  NAND U15302 ( .A(n14787), .B(n14786), .Z(n14788) );
  XNOR U15303 ( .A(n14789), .B(n14788), .Z(n14790) );
  XNOR U15304 ( .A(n14791), .B(n14790), .Z(n14792) );
  XNOR U15305 ( .A(n14793), .B(n14792), .Z(n14809) );
  OR U15306 ( .A(n14795), .B(n14794), .Z(n14799) );
  OR U15307 ( .A(n14797), .B(n14796), .Z(n14798) );
  AND U15308 ( .A(n14799), .B(n14798), .Z(n14807) );
  OR U15309 ( .A(n14801), .B(n14800), .Z(n14805) );
  OR U15310 ( .A(n14803), .B(n14802), .Z(n14804) );
  NAND U15311 ( .A(n14805), .B(n14804), .Z(n14806) );
  XNOR U15312 ( .A(n14807), .B(n14806), .Z(n14808) );
  XNOR U15313 ( .A(n14809), .B(n14808), .Z(n14810) );
  XNOR U15314 ( .A(n14811), .B(n14810), .Z(n14827) );
  NAND U15315 ( .A(n14813), .B(n14812), .Z(n14817) );
  OR U15316 ( .A(n14815), .B(n14814), .Z(n14816) );
  AND U15317 ( .A(n14817), .B(n14816), .Z(n14825) );
  NOR U15318 ( .A(n14819), .B(n14818), .Z(n14823) );
  ANDN U15319 ( .B(n14821), .A(n14820), .Z(n14822) );
  OR U15320 ( .A(n14823), .B(n14822), .Z(n14824) );
  XNOR U15321 ( .A(n14825), .B(n14824), .Z(n14826) );
  XNOR U15322 ( .A(n14827), .B(n14826), .Z(n14828) );
  XNOR U15323 ( .A(n14829), .B(n14828), .Z(n14845) );
  OR U15324 ( .A(n14831), .B(n14830), .Z(n14835) );
  NOR U15325 ( .A(n14833), .B(n14832), .Z(n14834) );
  ANDN U15326 ( .B(n14835), .A(n14834), .Z(n14843) );
  ANDN U15327 ( .B(n14837), .A(n14836), .Z(n14841) );
  NOR U15328 ( .A(n14839), .B(n14838), .Z(n14840) );
  OR U15329 ( .A(n14841), .B(n14840), .Z(n14842) );
  XNOR U15330 ( .A(n14843), .B(n14842), .Z(n14844) );
  XNOR U15331 ( .A(n14845), .B(n14844), .Z(n14846) );
  XNOR U15332 ( .A(n14847), .B(n14846), .Z(n14862) );
  NANDN U15333 ( .A(n14849), .B(n14848), .Z(n14852) );
  OR U15334 ( .A(n14850), .B(n16283), .Z(n14851) );
  AND U15335 ( .A(n14852), .B(n14851), .Z(n14860) );
  OR U15336 ( .A(n14854), .B(n14853), .Z(n14858) );
  OR U15337 ( .A(n14856), .B(n14855), .Z(n14857) );
  NAND U15338 ( .A(n14858), .B(n14857), .Z(n14859) );
  XNOR U15339 ( .A(n14860), .B(n14859), .Z(n14861) );
  XNOR U15340 ( .A(n14862), .B(n14861), .Z(n14863) );
  XNOR U15341 ( .A(n14864), .B(n14863), .Z(n14880) );
  OR U15342 ( .A(n14866), .B(n14865), .Z(n14870) );
  OR U15343 ( .A(n14868), .B(n14867), .Z(n14869) );
  AND U15344 ( .A(n14870), .B(n14869), .Z(n14878) );
  NANDN U15345 ( .A(n14872), .B(n14871), .Z(n14876) );
  NANDN U15346 ( .A(n14874), .B(n14873), .Z(n14875) );
  NAND U15347 ( .A(n14876), .B(n14875), .Z(n14877) );
  XNOR U15348 ( .A(n14878), .B(n14877), .Z(n14879) );
  XNOR U15349 ( .A(n14880), .B(n14879), .Z(n14881) );
  XNOR U15350 ( .A(n14882), .B(n14881), .Z(n14898) );
  OR U15351 ( .A(n14884), .B(n14883), .Z(n14888) );
  OR U15352 ( .A(n14886), .B(n14885), .Z(n14887) );
  AND U15353 ( .A(n14888), .B(n14887), .Z(n14896) );
  NANDN U15354 ( .A(n14890), .B(n14889), .Z(n14894) );
  NANDN U15355 ( .A(n14892), .B(n14891), .Z(n14893) );
  NAND U15356 ( .A(n14894), .B(n14893), .Z(n14895) );
  XNOR U15357 ( .A(n14896), .B(n14895), .Z(n14897) );
  XNOR U15358 ( .A(n14898), .B(n14897), .Z(n14899) );
  XNOR U15359 ( .A(n14900), .B(n14899), .Z(n14916) );
  NANDN U15360 ( .A(n14902), .B(n14901), .Z(n14906) );
  NANDN U15361 ( .A(n14904), .B(n14903), .Z(n14905) );
  AND U15362 ( .A(n14906), .B(n14905), .Z(n14914) );
  NOR U15363 ( .A(n14908), .B(n14907), .Z(n14912) );
  NOR U15364 ( .A(n14910), .B(n14909), .Z(n14911) );
  OR U15365 ( .A(n14912), .B(n14911), .Z(n14913) );
  XNOR U15366 ( .A(n14914), .B(n14913), .Z(n14915) );
  XNOR U15367 ( .A(n14916), .B(n14915), .Z(n14917) );
  XNOR U15368 ( .A(n14918), .B(n14917), .Z(n14934) );
  OR U15369 ( .A(n14920), .B(n14919), .Z(n14924) );
  OR U15370 ( .A(n14922), .B(n14921), .Z(n14923) );
  AND U15371 ( .A(n14924), .B(n14923), .Z(n14932) );
  OR U15372 ( .A(n14926), .B(n14925), .Z(n14930) );
  OR U15373 ( .A(n14928), .B(n14927), .Z(n14929) );
  NAND U15374 ( .A(n14930), .B(n14929), .Z(n14931) );
  XNOR U15375 ( .A(n14932), .B(n14931), .Z(n14933) );
  XNOR U15376 ( .A(n14934), .B(n14933), .Z(n14935) );
  XNOR U15377 ( .A(n14936), .B(n14935), .Z(n14952) );
  NANDN U15378 ( .A(n14938), .B(n14937), .Z(n14942) );
  NANDN U15379 ( .A(n14940), .B(n14939), .Z(n14941) );
  AND U15380 ( .A(n14942), .B(n14941), .Z(n14950) );
  OR U15381 ( .A(n14944), .B(n14943), .Z(n14948) );
  OR U15382 ( .A(n14946), .B(n14945), .Z(n14947) );
  NAND U15383 ( .A(n14948), .B(n14947), .Z(n14949) );
  XNOR U15384 ( .A(n14950), .B(n14949), .Z(n14951) );
  XNOR U15385 ( .A(n14952), .B(n14951), .Z(n14953) );
  XNOR U15386 ( .A(n14954), .B(n14953), .Z(n14970) );
  NANDN U15387 ( .A(n14956), .B(n14955), .Z(n14960) );
  NANDN U15388 ( .A(n14958), .B(n14957), .Z(n14959) );
  AND U15389 ( .A(n14960), .B(n14959), .Z(n14968) );
  OR U15390 ( .A(n14962), .B(n14961), .Z(n14966) );
  OR U15391 ( .A(n14964), .B(n14963), .Z(n14965) );
  NAND U15392 ( .A(n14966), .B(n14965), .Z(n14967) );
  XNOR U15393 ( .A(n14968), .B(n14967), .Z(n14969) );
  XNOR U15394 ( .A(n14970), .B(n14969), .Z(n14971) );
  XNOR U15395 ( .A(n14972), .B(n14971), .Z(n14988) );
  NANDN U15396 ( .A(n14974), .B(n14973), .Z(n14978) );
  NANDN U15397 ( .A(n14976), .B(n14975), .Z(n14977) );
  AND U15398 ( .A(n14978), .B(n14977), .Z(n14986) );
  NANDN U15399 ( .A(n14980), .B(n14979), .Z(n14984) );
  NANDN U15400 ( .A(n14982), .B(n14981), .Z(n14983) );
  NAND U15401 ( .A(n14984), .B(n14983), .Z(n14985) );
  XNOR U15402 ( .A(n14986), .B(n14985), .Z(n14987) );
  XNOR U15403 ( .A(n14988), .B(n14987), .Z(n14989) );
  XNOR U15404 ( .A(n14990), .B(n14989), .Z(n15006) );
  OR U15405 ( .A(n14992), .B(n14991), .Z(n14996) );
  OR U15406 ( .A(n14994), .B(n14993), .Z(n14995) );
  AND U15407 ( .A(n14996), .B(n14995), .Z(n15004) );
  ANDN U15408 ( .B(n14998), .A(n14997), .Z(n15002) );
  ANDN U15409 ( .B(n15000), .A(n14999), .Z(n15001) );
  OR U15410 ( .A(n15002), .B(n15001), .Z(n15003) );
  XNOR U15411 ( .A(n15004), .B(n15003), .Z(n15005) );
  XNOR U15412 ( .A(n15006), .B(n15005), .Z(n15007) );
  XNOR U15413 ( .A(n15008), .B(n15007), .Z(n15024) );
  NANDN U15414 ( .A(n15010), .B(n15009), .Z(n15014) );
  NANDN U15415 ( .A(n15012), .B(n15011), .Z(n15013) );
  AND U15416 ( .A(n15014), .B(n15013), .Z(n15022) );
  NANDN U15417 ( .A(n15016), .B(n15015), .Z(n15020) );
  NANDN U15418 ( .A(n15018), .B(n15017), .Z(n15019) );
  NAND U15419 ( .A(n15020), .B(n15019), .Z(n15021) );
  XNOR U15420 ( .A(n15022), .B(n15021), .Z(n15023) );
  XNOR U15421 ( .A(n15024), .B(n15023), .Z(n15025) );
  XNOR U15422 ( .A(n15026), .B(n15025), .Z(n15042) );
  NANDN U15423 ( .A(n15028), .B(n15027), .Z(n15032) );
  NOR U15424 ( .A(n15030), .B(n15029), .Z(n15031) );
  ANDN U15425 ( .B(n15032), .A(n15031), .Z(n15040) );
  NOR U15426 ( .A(n15034), .B(n15033), .Z(n15038) );
  NOR U15427 ( .A(n15036), .B(n15035), .Z(n15037) );
  OR U15428 ( .A(n15038), .B(n15037), .Z(n15039) );
  XNOR U15429 ( .A(n15040), .B(n15039), .Z(n15041) );
  XNOR U15430 ( .A(n15042), .B(n15041), .Z(n15043) );
  XNOR U15431 ( .A(n15044), .B(n15043), .Z(n15045) );
  NAND U15432 ( .A(opcode[0]), .B(opcode[1]), .Z(n17478) );
  NOR U15433 ( .A(opcode[2]), .B(n17478), .Z(n17458) );
  NANDN U15434 ( .A(n15045), .B(n17458), .Z(n15046) );
  NANDN U15435 ( .A(n2967), .B(x[63]), .Z(n15048) );
  ANDN U15436 ( .B(opcode[2]), .A(n17478), .Z(n17461) );
  IV U15437 ( .A(n17461), .Z(n17483) );
  NANDN U15438 ( .A(n17483), .B(\stack[1][63] ), .Z(n15047) );
  NAND U15439 ( .A(n15048), .B(n15047), .Z(n15049) );
  ANDN U15440 ( .B(n15050), .A(n15049), .Z(n15057) );
  ANDN U15441 ( .B(opcode[2]), .A(n15051), .Z(n17479) );
  NAND U15442 ( .A(\stack[1][63] ), .B(n17479), .Z(n15054) );
  XOR U15443 ( .A(n3221), .B(opcode[2]), .Z(n15053) );
  XOR U15444 ( .A(n3220), .B(opcode[1]), .Z(n15052) );
  NAND U15445 ( .A(n15053), .B(n15052), .Z(n17481) );
  IV U15446 ( .A(n17481), .Z(n17467) );
  ANDN U15447 ( .B(n15054), .A(n17467), .Z(n15055) );
  NANDN U15448 ( .A(n15055), .B(o[63]), .Z(n15056) );
  NAND U15449 ( .A(n15057), .B(n15056), .Z(n2134) );
  NANDN U15450 ( .A(n2967), .B(\stack[6][62] ), .Z(n15059) );
  NANDN U15451 ( .A(n17471), .B(\stack[7][62] ), .Z(n15058) );
  NAND U15452 ( .A(n15059), .B(n15058), .Z(n2135) );
  NANDN U15453 ( .A(n2967), .B(\stack[5][62] ), .Z(n15061) );
  NANDN U15454 ( .A(n17472), .B(\stack[7][62] ), .Z(n15060) );
  AND U15455 ( .A(n15061), .B(n15060), .Z(n15063) );
  NANDN U15456 ( .A(n17475), .B(\stack[6][62] ), .Z(n15062) );
  NAND U15457 ( .A(n15063), .B(n15062), .Z(n2136) );
  NANDN U15458 ( .A(n2967), .B(\stack[4][62] ), .Z(n15065) );
  NANDN U15459 ( .A(n17472), .B(\stack[6][62] ), .Z(n15064) );
  AND U15460 ( .A(n15065), .B(n15064), .Z(n15067) );
  NANDN U15461 ( .A(n17475), .B(\stack[5][62] ), .Z(n15066) );
  NAND U15462 ( .A(n15067), .B(n15066), .Z(n2137) );
  NANDN U15463 ( .A(n2967), .B(\stack[3][62] ), .Z(n15069) );
  NANDN U15464 ( .A(n17472), .B(\stack[5][62] ), .Z(n15068) );
  AND U15465 ( .A(n15069), .B(n15068), .Z(n15071) );
  NANDN U15466 ( .A(n17475), .B(\stack[4][62] ), .Z(n15070) );
  NAND U15467 ( .A(n15071), .B(n15070), .Z(n2138) );
  NANDN U15468 ( .A(n2967), .B(\stack[2][62] ), .Z(n15073) );
  NANDN U15469 ( .A(n17472), .B(\stack[4][62] ), .Z(n15072) );
  AND U15470 ( .A(n15073), .B(n15072), .Z(n15075) );
  NANDN U15471 ( .A(n17475), .B(\stack[3][62] ), .Z(n15074) );
  NAND U15472 ( .A(n15075), .B(n15074), .Z(n2139) );
  NANDN U15473 ( .A(n2967), .B(\stack[1][62] ), .Z(n15077) );
  NANDN U15474 ( .A(n17472), .B(\stack[3][62] ), .Z(n15076) );
  AND U15475 ( .A(n15077), .B(n15076), .Z(n15079) );
  NANDN U15476 ( .A(n17475), .B(\stack[2][62] ), .Z(n15078) );
  NAND U15477 ( .A(n15079), .B(n15078), .Z(n2140) );
  NANDN U15478 ( .A(n2967), .B(o[62]), .Z(n15081) );
  NANDN U15479 ( .A(n17472), .B(\stack[2][62] ), .Z(n15080) );
  AND U15480 ( .A(n15081), .B(n15080), .Z(n15083) );
  NANDN U15481 ( .A(n17475), .B(\stack[1][62] ), .Z(n15082) );
  NAND U15482 ( .A(n15083), .B(n15082), .Z(n2141) );
  NAND U15483 ( .A(\stack[1][62] ), .B(n17479), .Z(n15084) );
  NANDN U15484 ( .A(n17467), .B(n15084), .Z(n15085) );
  AND U15485 ( .A(n15085), .B(o[62]), .Z(n15094) );
  XNOR U15486 ( .A(n15087), .B(n15086), .Z(n15088) );
  NAND U15487 ( .A(n15088), .B(n17458), .Z(n15092) );
  NANDN U15488 ( .A(n2967), .B(x[62]), .Z(n15090) );
  NANDN U15489 ( .A(n17483), .B(\stack[1][62] ), .Z(n15089) );
  AND U15490 ( .A(n15090), .B(n15089), .Z(n15091) );
  NAND U15491 ( .A(n15092), .B(n15091), .Z(n15093) );
  NOR U15492 ( .A(n15094), .B(n15093), .Z(n15095) );
  NANDN U15493 ( .A(n2967), .B(\stack[6][61] ), .Z(n15097) );
  NANDN U15494 ( .A(n17471), .B(\stack[7][61] ), .Z(n15096) );
  NAND U15495 ( .A(n15097), .B(n15096), .Z(n2143) );
  NANDN U15496 ( .A(n2967), .B(\stack[5][61] ), .Z(n15099) );
  NANDN U15497 ( .A(n17472), .B(\stack[7][61] ), .Z(n15098) );
  AND U15498 ( .A(n15099), .B(n15098), .Z(n15101) );
  NANDN U15499 ( .A(n17475), .B(\stack[6][61] ), .Z(n15100) );
  NAND U15500 ( .A(n15101), .B(n15100), .Z(n2144) );
  NANDN U15501 ( .A(n2967), .B(\stack[4][61] ), .Z(n15103) );
  NANDN U15502 ( .A(n17472), .B(\stack[6][61] ), .Z(n15102) );
  AND U15503 ( .A(n15103), .B(n15102), .Z(n15105) );
  NANDN U15504 ( .A(n17475), .B(\stack[5][61] ), .Z(n15104) );
  NAND U15505 ( .A(n15105), .B(n15104), .Z(n2145) );
  NANDN U15506 ( .A(n2967), .B(\stack[3][61] ), .Z(n15107) );
  NANDN U15507 ( .A(n17472), .B(\stack[5][61] ), .Z(n15106) );
  AND U15508 ( .A(n15107), .B(n15106), .Z(n15109) );
  NANDN U15509 ( .A(n17475), .B(\stack[4][61] ), .Z(n15108) );
  NAND U15510 ( .A(n15109), .B(n15108), .Z(n2146) );
  NANDN U15511 ( .A(n2967), .B(\stack[2][61] ), .Z(n15111) );
  NANDN U15512 ( .A(n17472), .B(\stack[4][61] ), .Z(n15110) );
  AND U15513 ( .A(n15111), .B(n15110), .Z(n15113) );
  NANDN U15514 ( .A(n17475), .B(\stack[3][61] ), .Z(n15112) );
  NAND U15515 ( .A(n15113), .B(n15112), .Z(n2147) );
  NANDN U15516 ( .A(n2967), .B(\stack[1][61] ), .Z(n15115) );
  NANDN U15517 ( .A(n17472), .B(\stack[3][61] ), .Z(n15114) );
  AND U15518 ( .A(n15115), .B(n15114), .Z(n15117) );
  NANDN U15519 ( .A(n17475), .B(\stack[2][61] ), .Z(n15116) );
  NAND U15520 ( .A(n15117), .B(n15116), .Z(n2148) );
  NANDN U15521 ( .A(n2967), .B(o[61]), .Z(n15119) );
  NANDN U15522 ( .A(n17472), .B(\stack[2][61] ), .Z(n15118) );
  AND U15523 ( .A(n15119), .B(n15118), .Z(n15121) );
  NANDN U15524 ( .A(n17475), .B(\stack[1][61] ), .Z(n15120) );
  NAND U15525 ( .A(n15121), .B(n15120), .Z(n2149) );
  NAND U15526 ( .A(\stack[1][61] ), .B(n17479), .Z(n15122) );
  NANDN U15527 ( .A(n17467), .B(n15122), .Z(n15123) );
  AND U15528 ( .A(n15123), .B(o[61]), .Z(n15132) );
  XNOR U15529 ( .A(n15125), .B(n15124), .Z(n15126) );
  NAND U15530 ( .A(n15126), .B(n17458), .Z(n15130) );
  NANDN U15531 ( .A(n2967), .B(x[61]), .Z(n15128) );
  NANDN U15532 ( .A(n17483), .B(\stack[1][61] ), .Z(n15127) );
  AND U15533 ( .A(n15128), .B(n15127), .Z(n15129) );
  NAND U15534 ( .A(n15130), .B(n15129), .Z(n15131) );
  NOR U15535 ( .A(n15132), .B(n15131), .Z(n15133) );
  NANDN U15536 ( .A(n2967), .B(\stack[6][60] ), .Z(n15135) );
  NANDN U15537 ( .A(n17471), .B(\stack[7][60] ), .Z(n15134) );
  NAND U15538 ( .A(n15135), .B(n15134), .Z(n2151) );
  NANDN U15539 ( .A(n2967), .B(\stack[5][60] ), .Z(n15137) );
  NANDN U15540 ( .A(n17472), .B(\stack[7][60] ), .Z(n15136) );
  AND U15541 ( .A(n15137), .B(n15136), .Z(n15139) );
  NANDN U15542 ( .A(n17475), .B(\stack[6][60] ), .Z(n15138) );
  NAND U15543 ( .A(n15139), .B(n15138), .Z(n2152) );
  NANDN U15544 ( .A(n2967), .B(\stack[4][60] ), .Z(n15141) );
  NANDN U15545 ( .A(n17472), .B(\stack[6][60] ), .Z(n15140) );
  AND U15546 ( .A(n15141), .B(n15140), .Z(n15143) );
  NANDN U15547 ( .A(n17475), .B(\stack[5][60] ), .Z(n15142) );
  NAND U15548 ( .A(n15143), .B(n15142), .Z(n2153) );
  NANDN U15549 ( .A(n2967), .B(\stack[3][60] ), .Z(n15145) );
  NANDN U15550 ( .A(n17472), .B(\stack[5][60] ), .Z(n15144) );
  AND U15551 ( .A(n15145), .B(n15144), .Z(n15147) );
  NANDN U15552 ( .A(n17475), .B(\stack[4][60] ), .Z(n15146) );
  NAND U15553 ( .A(n15147), .B(n15146), .Z(n2154) );
  NANDN U15554 ( .A(n2967), .B(\stack[2][60] ), .Z(n15149) );
  NANDN U15555 ( .A(n17472), .B(\stack[4][60] ), .Z(n15148) );
  AND U15556 ( .A(n15149), .B(n15148), .Z(n15151) );
  NANDN U15557 ( .A(n17475), .B(\stack[3][60] ), .Z(n15150) );
  NAND U15558 ( .A(n15151), .B(n15150), .Z(n2155) );
  IV U15559 ( .A(\stack[1][60] ), .Z(n15160) );
  NANDN U15560 ( .A(n15160), .B(n17471), .Z(n15153) );
  NANDN U15561 ( .A(n17472), .B(\stack[3][60] ), .Z(n15152) );
  AND U15562 ( .A(n15153), .B(n15152), .Z(n15155) );
  NANDN U15563 ( .A(n17475), .B(\stack[2][60] ), .Z(n15154) );
  NAND U15564 ( .A(n15155), .B(n15154), .Z(n2156) );
  NANDN U15565 ( .A(n2967), .B(o[60]), .Z(n15157) );
  NANDN U15566 ( .A(n17472), .B(\stack[2][60] ), .Z(n15156) );
  AND U15567 ( .A(n15157), .B(n15156), .Z(n15159) );
  OR U15568 ( .A(n17475), .B(n15160), .Z(n15158) );
  NAND U15569 ( .A(n15159), .B(n15158), .Z(n2157) );
  NANDN U15570 ( .A(n15160), .B(n17479), .Z(n15161) );
  NANDN U15571 ( .A(n17467), .B(n15161), .Z(n15162) );
  AND U15572 ( .A(n15162), .B(o[60]), .Z(n15171) );
  XNOR U15573 ( .A(n15164), .B(n15163), .Z(n15165) );
  NAND U15574 ( .A(n15165), .B(n17458), .Z(n15169) );
  NANDN U15575 ( .A(n2967), .B(x[60]), .Z(n15167) );
  NANDN U15576 ( .A(n17483), .B(\stack[1][60] ), .Z(n15166) );
  AND U15577 ( .A(n15167), .B(n15166), .Z(n15168) );
  NAND U15578 ( .A(n15169), .B(n15168), .Z(n15170) );
  NOR U15579 ( .A(n15171), .B(n15170), .Z(n15172) );
  NANDN U15580 ( .A(n2967), .B(\stack[6][59] ), .Z(n15174) );
  NANDN U15581 ( .A(n17471), .B(\stack[7][59] ), .Z(n15173) );
  NAND U15582 ( .A(n15174), .B(n15173), .Z(n2159) );
  NANDN U15583 ( .A(n2967), .B(\stack[5][59] ), .Z(n15176) );
  NANDN U15584 ( .A(n17472), .B(\stack[7][59] ), .Z(n15175) );
  AND U15585 ( .A(n15176), .B(n15175), .Z(n15178) );
  NANDN U15586 ( .A(n17475), .B(\stack[6][59] ), .Z(n15177) );
  NAND U15587 ( .A(n15178), .B(n15177), .Z(n2160) );
  NANDN U15588 ( .A(n2967), .B(\stack[4][59] ), .Z(n15180) );
  NANDN U15589 ( .A(n17472), .B(\stack[6][59] ), .Z(n15179) );
  AND U15590 ( .A(n15180), .B(n15179), .Z(n15182) );
  NANDN U15591 ( .A(n17475), .B(\stack[5][59] ), .Z(n15181) );
  NAND U15592 ( .A(n15182), .B(n15181), .Z(n2161) );
  NANDN U15593 ( .A(n2967), .B(\stack[3][59] ), .Z(n15184) );
  NANDN U15594 ( .A(n17472), .B(\stack[5][59] ), .Z(n15183) );
  AND U15595 ( .A(n15184), .B(n15183), .Z(n15186) );
  NANDN U15596 ( .A(n17475), .B(\stack[4][59] ), .Z(n15185) );
  NAND U15597 ( .A(n15186), .B(n15185), .Z(n2162) );
  NANDN U15598 ( .A(n2967), .B(\stack[2][59] ), .Z(n15188) );
  NANDN U15599 ( .A(n17472), .B(\stack[4][59] ), .Z(n15187) );
  AND U15600 ( .A(n15188), .B(n15187), .Z(n15190) );
  NANDN U15601 ( .A(n17475), .B(\stack[3][59] ), .Z(n15189) );
  NAND U15602 ( .A(n15190), .B(n15189), .Z(n2163) );
  IV U15603 ( .A(\stack[1][59] ), .Z(n15199) );
  NANDN U15604 ( .A(n15199), .B(n17471), .Z(n15192) );
  NANDN U15605 ( .A(n17472), .B(\stack[3][59] ), .Z(n15191) );
  AND U15606 ( .A(n15192), .B(n15191), .Z(n15194) );
  NANDN U15607 ( .A(n17475), .B(\stack[2][59] ), .Z(n15193) );
  NAND U15608 ( .A(n15194), .B(n15193), .Z(n2164) );
  NANDN U15609 ( .A(n2967), .B(o[59]), .Z(n15196) );
  NANDN U15610 ( .A(n17472), .B(\stack[2][59] ), .Z(n15195) );
  AND U15611 ( .A(n15196), .B(n15195), .Z(n15198) );
  OR U15612 ( .A(n17475), .B(n15199), .Z(n15197) );
  NAND U15613 ( .A(n15198), .B(n15197), .Z(n2165) );
  NANDN U15614 ( .A(n15199), .B(n17479), .Z(n15200) );
  NANDN U15615 ( .A(n17467), .B(n15200), .Z(n15201) );
  AND U15616 ( .A(n15201), .B(o[59]), .Z(n15210) );
  XNOR U15617 ( .A(n15203), .B(n15202), .Z(n15204) );
  NAND U15618 ( .A(n15204), .B(n17458), .Z(n15208) );
  NANDN U15619 ( .A(n2967), .B(x[59]), .Z(n15206) );
  NANDN U15620 ( .A(n17483), .B(\stack[1][59] ), .Z(n15205) );
  AND U15621 ( .A(n15206), .B(n15205), .Z(n15207) );
  NAND U15622 ( .A(n15208), .B(n15207), .Z(n15209) );
  NOR U15623 ( .A(n15210), .B(n15209), .Z(n15211) );
  NANDN U15624 ( .A(n2967), .B(\stack[6][58] ), .Z(n15213) );
  NANDN U15625 ( .A(n17471), .B(\stack[7][58] ), .Z(n15212) );
  NAND U15626 ( .A(n15213), .B(n15212), .Z(n2167) );
  NANDN U15627 ( .A(n2967), .B(\stack[5][58] ), .Z(n15215) );
  NANDN U15628 ( .A(n17472), .B(\stack[7][58] ), .Z(n15214) );
  AND U15629 ( .A(n15215), .B(n15214), .Z(n15217) );
  NANDN U15630 ( .A(n17475), .B(\stack[6][58] ), .Z(n15216) );
  NAND U15631 ( .A(n15217), .B(n15216), .Z(n2168) );
  NANDN U15632 ( .A(n2967), .B(\stack[4][58] ), .Z(n15219) );
  NANDN U15633 ( .A(n17472), .B(\stack[6][58] ), .Z(n15218) );
  AND U15634 ( .A(n15219), .B(n15218), .Z(n15221) );
  NANDN U15635 ( .A(n17475), .B(\stack[5][58] ), .Z(n15220) );
  NAND U15636 ( .A(n15221), .B(n15220), .Z(n2169) );
  NANDN U15637 ( .A(n2967), .B(\stack[3][58] ), .Z(n15223) );
  NANDN U15638 ( .A(n17472), .B(\stack[5][58] ), .Z(n15222) );
  AND U15639 ( .A(n15223), .B(n15222), .Z(n15225) );
  NANDN U15640 ( .A(n17475), .B(\stack[4][58] ), .Z(n15224) );
  NAND U15641 ( .A(n15225), .B(n15224), .Z(n2170) );
  NANDN U15642 ( .A(n2967), .B(\stack[2][58] ), .Z(n15227) );
  NANDN U15643 ( .A(n17472), .B(\stack[4][58] ), .Z(n15226) );
  AND U15644 ( .A(n15227), .B(n15226), .Z(n15229) );
  NANDN U15645 ( .A(n17475), .B(\stack[3][58] ), .Z(n15228) );
  NAND U15646 ( .A(n15229), .B(n15228), .Z(n2171) );
  IV U15647 ( .A(\stack[1][58] ), .Z(n15238) );
  NANDN U15648 ( .A(n15238), .B(n17471), .Z(n15231) );
  NANDN U15649 ( .A(n17472), .B(\stack[3][58] ), .Z(n15230) );
  AND U15650 ( .A(n15231), .B(n15230), .Z(n15233) );
  NANDN U15651 ( .A(n17475), .B(\stack[2][58] ), .Z(n15232) );
  NAND U15652 ( .A(n15233), .B(n15232), .Z(n2172) );
  NANDN U15653 ( .A(n2967), .B(o[58]), .Z(n15235) );
  NANDN U15654 ( .A(n17472), .B(\stack[2][58] ), .Z(n15234) );
  AND U15655 ( .A(n15235), .B(n15234), .Z(n15237) );
  OR U15656 ( .A(n17475), .B(n15238), .Z(n15236) );
  NAND U15657 ( .A(n15237), .B(n15236), .Z(n2173) );
  NANDN U15658 ( .A(n15238), .B(n17479), .Z(n15239) );
  NANDN U15659 ( .A(n17467), .B(n15239), .Z(n15240) );
  AND U15660 ( .A(n15240), .B(o[58]), .Z(n15249) );
  XNOR U15661 ( .A(n15242), .B(n15241), .Z(n15243) );
  NAND U15662 ( .A(n15243), .B(n17458), .Z(n15247) );
  NANDN U15663 ( .A(n2967), .B(x[58]), .Z(n15245) );
  NANDN U15664 ( .A(n17483), .B(\stack[1][58] ), .Z(n15244) );
  AND U15665 ( .A(n15245), .B(n15244), .Z(n15246) );
  NAND U15666 ( .A(n15247), .B(n15246), .Z(n15248) );
  NOR U15667 ( .A(n15249), .B(n15248), .Z(n15250) );
  NANDN U15668 ( .A(n2967), .B(\stack[6][57] ), .Z(n15252) );
  NANDN U15669 ( .A(n17471), .B(\stack[7][57] ), .Z(n15251) );
  NAND U15670 ( .A(n15252), .B(n15251), .Z(n2175) );
  NANDN U15671 ( .A(n2967), .B(\stack[5][57] ), .Z(n15254) );
  NANDN U15672 ( .A(n17472), .B(\stack[7][57] ), .Z(n15253) );
  AND U15673 ( .A(n15254), .B(n15253), .Z(n15256) );
  NANDN U15674 ( .A(n17475), .B(\stack[6][57] ), .Z(n15255) );
  NAND U15675 ( .A(n15256), .B(n15255), .Z(n2176) );
  NANDN U15676 ( .A(n2967), .B(\stack[4][57] ), .Z(n15258) );
  NANDN U15677 ( .A(n17472), .B(\stack[6][57] ), .Z(n15257) );
  AND U15678 ( .A(n15258), .B(n15257), .Z(n15260) );
  NANDN U15679 ( .A(n17475), .B(\stack[5][57] ), .Z(n15259) );
  NAND U15680 ( .A(n15260), .B(n15259), .Z(n2177) );
  NANDN U15681 ( .A(n2967), .B(\stack[3][57] ), .Z(n15262) );
  NANDN U15682 ( .A(n17472), .B(\stack[5][57] ), .Z(n15261) );
  AND U15683 ( .A(n15262), .B(n15261), .Z(n15264) );
  NANDN U15684 ( .A(n17475), .B(\stack[4][57] ), .Z(n15263) );
  NAND U15685 ( .A(n15264), .B(n15263), .Z(n2178) );
  NANDN U15686 ( .A(n2967), .B(\stack[2][57] ), .Z(n15266) );
  NANDN U15687 ( .A(n17472), .B(\stack[4][57] ), .Z(n15265) );
  AND U15688 ( .A(n15266), .B(n15265), .Z(n15268) );
  NANDN U15689 ( .A(n17475), .B(\stack[3][57] ), .Z(n15267) );
  NAND U15690 ( .A(n15268), .B(n15267), .Z(n2179) );
  NANDN U15691 ( .A(n2967), .B(\stack[1][57] ), .Z(n15270) );
  NANDN U15692 ( .A(n17472), .B(\stack[3][57] ), .Z(n15269) );
  AND U15693 ( .A(n15270), .B(n15269), .Z(n15272) );
  NANDN U15694 ( .A(n17475), .B(\stack[2][57] ), .Z(n15271) );
  NAND U15695 ( .A(n15272), .B(n15271), .Z(n2180) );
  NANDN U15696 ( .A(n2967), .B(o[57]), .Z(n15274) );
  NANDN U15697 ( .A(n17472), .B(\stack[2][57] ), .Z(n15273) );
  AND U15698 ( .A(n15274), .B(n15273), .Z(n15276) );
  NANDN U15699 ( .A(n17475), .B(\stack[1][57] ), .Z(n15275) );
  NAND U15700 ( .A(n15276), .B(n15275), .Z(n2181) );
  NAND U15701 ( .A(\stack[1][57] ), .B(n17479), .Z(n15277) );
  NANDN U15702 ( .A(n17467), .B(n15277), .Z(n15278) );
  AND U15703 ( .A(n15278), .B(o[57]), .Z(n15287) );
  XNOR U15704 ( .A(n15280), .B(n15279), .Z(n15281) );
  NAND U15705 ( .A(n15281), .B(n17458), .Z(n15285) );
  NANDN U15706 ( .A(n2967), .B(x[57]), .Z(n15283) );
  NANDN U15707 ( .A(n17483), .B(\stack[1][57] ), .Z(n15282) );
  AND U15708 ( .A(n15283), .B(n15282), .Z(n15284) );
  NAND U15709 ( .A(n15285), .B(n15284), .Z(n15286) );
  NOR U15710 ( .A(n15287), .B(n15286), .Z(n15288) );
  NANDN U15711 ( .A(n2967), .B(\stack[6][56] ), .Z(n15290) );
  NANDN U15712 ( .A(n17471), .B(\stack[7][56] ), .Z(n15289) );
  NAND U15713 ( .A(n15290), .B(n15289), .Z(n2183) );
  NANDN U15714 ( .A(n2967), .B(\stack[5][56] ), .Z(n15292) );
  NANDN U15715 ( .A(n17472), .B(\stack[7][56] ), .Z(n15291) );
  AND U15716 ( .A(n15292), .B(n15291), .Z(n15294) );
  NANDN U15717 ( .A(n17475), .B(\stack[6][56] ), .Z(n15293) );
  NAND U15718 ( .A(n15294), .B(n15293), .Z(n2184) );
  NANDN U15719 ( .A(n2967), .B(\stack[4][56] ), .Z(n15296) );
  NANDN U15720 ( .A(n17472), .B(\stack[6][56] ), .Z(n15295) );
  AND U15721 ( .A(n15296), .B(n15295), .Z(n15298) );
  NANDN U15722 ( .A(n17475), .B(\stack[5][56] ), .Z(n15297) );
  NAND U15723 ( .A(n15298), .B(n15297), .Z(n2185) );
  NANDN U15724 ( .A(n2967), .B(\stack[3][56] ), .Z(n15300) );
  NANDN U15725 ( .A(n17472), .B(\stack[5][56] ), .Z(n15299) );
  AND U15726 ( .A(n15300), .B(n15299), .Z(n15302) );
  NANDN U15727 ( .A(n17475), .B(\stack[4][56] ), .Z(n15301) );
  NAND U15728 ( .A(n15302), .B(n15301), .Z(n2186) );
  NANDN U15729 ( .A(n2967), .B(\stack[2][56] ), .Z(n15304) );
  NANDN U15730 ( .A(n17472), .B(\stack[4][56] ), .Z(n15303) );
  AND U15731 ( .A(n15304), .B(n15303), .Z(n15306) );
  NANDN U15732 ( .A(n17475), .B(\stack[3][56] ), .Z(n15305) );
  NAND U15733 ( .A(n15306), .B(n15305), .Z(n2187) );
  NANDN U15734 ( .A(n15315), .B(n17471), .Z(n15308) );
  NANDN U15735 ( .A(n17472), .B(\stack[3][56] ), .Z(n15307) );
  AND U15736 ( .A(n15308), .B(n15307), .Z(n15310) );
  NANDN U15737 ( .A(n17475), .B(\stack[2][56] ), .Z(n15309) );
  NAND U15738 ( .A(n15310), .B(n15309), .Z(n2188) );
  NANDN U15739 ( .A(n2967), .B(o[56]), .Z(n15312) );
  NANDN U15740 ( .A(n17472), .B(\stack[2][56] ), .Z(n15311) );
  AND U15741 ( .A(n15312), .B(n15311), .Z(n15314) );
  OR U15742 ( .A(n17475), .B(n15315), .Z(n15313) );
  NAND U15743 ( .A(n15314), .B(n15313), .Z(n2189) );
  NANDN U15744 ( .A(n15315), .B(n17479), .Z(n15316) );
  NANDN U15745 ( .A(n17467), .B(n15316), .Z(n15317) );
  AND U15746 ( .A(n15317), .B(o[56]), .Z(n15326) );
  XNOR U15747 ( .A(n15319), .B(n15318), .Z(n15320) );
  NAND U15748 ( .A(n15320), .B(n17458), .Z(n15324) );
  NANDN U15749 ( .A(n2967), .B(x[56]), .Z(n15322) );
  NANDN U15750 ( .A(n17483), .B(\stack[1][56] ), .Z(n15321) );
  AND U15751 ( .A(n15322), .B(n15321), .Z(n15323) );
  NAND U15752 ( .A(n15324), .B(n15323), .Z(n15325) );
  NOR U15753 ( .A(n15326), .B(n15325), .Z(n15327) );
  NANDN U15754 ( .A(n2967), .B(\stack[6][55] ), .Z(n15329) );
  NANDN U15755 ( .A(n17471), .B(\stack[7][55] ), .Z(n15328) );
  NAND U15756 ( .A(n15329), .B(n15328), .Z(n2191) );
  NANDN U15757 ( .A(n2967), .B(\stack[5][55] ), .Z(n15331) );
  NANDN U15758 ( .A(n17472), .B(\stack[7][55] ), .Z(n15330) );
  AND U15759 ( .A(n15331), .B(n15330), .Z(n15333) );
  NANDN U15760 ( .A(n17475), .B(\stack[6][55] ), .Z(n15332) );
  NAND U15761 ( .A(n15333), .B(n15332), .Z(n2192) );
  NANDN U15762 ( .A(n2967), .B(\stack[4][55] ), .Z(n15335) );
  NANDN U15763 ( .A(n17472), .B(\stack[6][55] ), .Z(n15334) );
  AND U15764 ( .A(n15335), .B(n15334), .Z(n15337) );
  NANDN U15765 ( .A(n17475), .B(\stack[5][55] ), .Z(n15336) );
  NAND U15766 ( .A(n15337), .B(n15336), .Z(n2193) );
  NANDN U15767 ( .A(n2967), .B(\stack[3][55] ), .Z(n15339) );
  NANDN U15768 ( .A(n17472), .B(\stack[5][55] ), .Z(n15338) );
  AND U15769 ( .A(n15339), .B(n15338), .Z(n15341) );
  NANDN U15770 ( .A(n17475), .B(\stack[4][55] ), .Z(n15340) );
  NAND U15771 ( .A(n15341), .B(n15340), .Z(n2194) );
  NANDN U15772 ( .A(n2967), .B(\stack[2][55] ), .Z(n15343) );
  NANDN U15773 ( .A(n17472), .B(\stack[4][55] ), .Z(n15342) );
  AND U15774 ( .A(n15343), .B(n15342), .Z(n15345) );
  NANDN U15775 ( .A(n17475), .B(\stack[3][55] ), .Z(n15344) );
  NAND U15776 ( .A(n15345), .B(n15344), .Z(n2195) );
  NANDN U15777 ( .A(n2967), .B(\stack[1][55] ), .Z(n15347) );
  NANDN U15778 ( .A(n17472), .B(\stack[3][55] ), .Z(n15346) );
  AND U15779 ( .A(n15347), .B(n15346), .Z(n15349) );
  NANDN U15780 ( .A(n17475), .B(\stack[2][55] ), .Z(n15348) );
  NAND U15781 ( .A(n15349), .B(n15348), .Z(n2196) );
  NANDN U15782 ( .A(n2967), .B(o[55]), .Z(n15351) );
  NANDN U15783 ( .A(n17472), .B(\stack[2][55] ), .Z(n15350) );
  AND U15784 ( .A(n15351), .B(n15350), .Z(n15353) );
  NANDN U15785 ( .A(n17475), .B(\stack[1][55] ), .Z(n15352) );
  NAND U15786 ( .A(n15353), .B(n15352), .Z(n2197) );
  NAND U15787 ( .A(\stack[1][55] ), .B(n17479), .Z(n15354) );
  NANDN U15788 ( .A(n17467), .B(n15354), .Z(n15355) );
  AND U15789 ( .A(n15355), .B(o[55]), .Z(n15364) );
  XNOR U15790 ( .A(n15357), .B(n15356), .Z(n15358) );
  NAND U15791 ( .A(n15358), .B(n17458), .Z(n15362) );
  NANDN U15792 ( .A(n2967), .B(x[55]), .Z(n15360) );
  NANDN U15793 ( .A(n17483), .B(\stack[1][55] ), .Z(n15359) );
  AND U15794 ( .A(n15360), .B(n15359), .Z(n15361) );
  NAND U15795 ( .A(n15362), .B(n15361), .Z(n15363) );
  NOR U15796 ( .A(n15364), .B(n15363), .Z(n15365) );
  NANDN U15797 ( .A(n2967), .B(\stack[6][54] ), .Z(n15367) );
  NANDN U15798 ( .A(n17471), .B(\stack[7][54] ), .Z(n15366) );
  NAND U15799 ( .A(n15367), .B(n15366), .Z(n2199) );
  NANDN U15800 ( .A(n2967), .B(\stack[5][54] ), .Z(n15369) );
  NANDN U15801 ( .A(n17472), .B(\stack[7][54] ), .Z(n15368) );
  AND U15802 ( .A(n15369), .B(n15368), .Z(n15371) );
  NANDN U15803 ( .A(n17475), .B(\stack[6][54] ), .Z(n15370) );
  NAND U15804 ( .A(n15371), .B(n15370), .Z(n2200) );
  NANDN U15805 ( .A(n2967), .B(\stack[4][54] ), .Z(n15373) );
  NANDN U15806 ( .A(n17472), .B(\stack[6][54] ), .Z(n15372) );
  AND U15807 ( .A(n15373), .B(n15372), .Z(n15375) );
  NANDN U15808 ( .A(n17475), .B(\stack[5][54] ), .Z(n15374) );
  NAND U15809 ( .A(n15375), .B(n15374), .Z(n2201) );
  NANDN U15810 ( .A(n2967), .B(\stack[3][54] ), .Z(n15377) );
  NANDN U15811 ( .A(n17472), .B(\stack[5][54] ), .Z(n15376) );
  AND U15812 ( .A(n15377), .B(n15376), .Z(n15379) );
  NANDN U15813 ( .A(n17475), .B(\stack[4][54] ), .Z(n15378) );
  NAND U15814 ( .A(n15379), .B(n15378), .Z(n2202) );
  NANDN U15815 ( .A(n2967), .B(\stack[2][54] ), .Z(n15381) );
  NANDN U15816 ( .A(n17472), .B(\stack[4][54] ), .Z(n15380) );
  AND U15817 ( .A(n15381), .B(n15380), .Z(n15383) );
  NANDN U15818 ( .A(n17475), .B(\stack[3][54] ), .Z(n15382) );
  NAND U15819 ( .A(n15383), .B(n15382), .Z(n2203) );
  NANDN U15820 ( .A(n2967), .B(\stack[1][54] ), .Z(n15385) );
  NANDN U15821 ( .A(n17472), .B(\stack[3][54] ), .Z(n15384) );
  AND U15822 ( .A(n15385), .B(n15384), .Z(n15387) );
  NANDN U15823 ( .A(n17475), .B(\stack[2][54] ), .Z(n15386) );
  NAND U15824 ( .A(n15387), .B(n15386), .Z(n2204) );
  NANDN U15825 ( .A(n2967), .B(o[54]), .Z(n15389) );
  NANDN U15826 ( .A(n17472), .B(\stack[2][54] ), .Z(n15388) );
  AND U15827 ( .A(n15389), .B(n15388), .Z(n15391) );
  NANDN U15828 ( .A(n17475), .B(\stack[1][54] ), .Z(n15390) );
  NAND U15829 ( .A(n15391), .B(n15390), .Z(n2205) );
  NAND U15830 ( .A(\stack[1][54] ), .B(n17479), .Z(n15392) );
  NANDN U15831 ( .A(n17467), .B(n15392), .Z(n15393) );
  AND U15832 ( .A(n15393), .B(o[54]), .Z(n15402) );
  XNOR U15833 ( .A(n15395), .B(n15394), .Z(n15396) );
  NAND U15834 ( .A(n15396), .B(n17458), .Z(n15400) );
  NANDN U15835 ( .A(n2967), .B(x[54]), .Z(n15398) );
  NANDN U15836 ( .A(n17483), .B(\stack[1][54] ), .Z(n15397) );
  AND U15837 ( .A(n15398), .B(n15397), .Z(n15399) );
  NAND U15838 ( .A(n15400), .B(n15399), .Z(n15401) );
  NOR U15839 ( .A(n15402), .B(n15401), .Z(n15403) );
  NANDN U15840 ( .A(n2967), .B(\stack[6][53] ), .Z(n15405) );
  NANDN U15841 ( .A(n17471), .B(\stack[7][53] ), .Z(n15404) );
  NAND U15842 ( .A(n15405), .B(n15404), .Z(n2207) );
  NANDN U15843 ( .A(n2967), .B(\stack[5][53] ), .Z(n15407) );
  NANDN U15844 ( .A(n17472), .B(\stack[7][53] ), .Z(n15406) );
  AND U15845 ( .A(n15407), .B(n15406), .Z(n15409) );
  NANDN U15846 ( .A(n17475), .B(\stack[6][53] ), .Z(n15408) );
  NAND U15847 ( .A(n15409), .B(n15408), .Z(n2208) );
  NANDN U15848 ( .A(n2967), .B(\stack[4][53] ), .Z(n15411) );
  NANDN U15849 ( .A(n17472), .B(\stack[6][53] ), .Z(n15410) );
  AND U15850 ( .A(n15411), .B(n15410), .Z(n15413) );
  NANDN U15851 ( .A(n17475), .B(\stack[5][53] ), .Z(n15412) );
  NAND U15852 ( .A(n15413), .B(n15412), .Z(n2209) );
  NANDN U15853 ( .A(n2967), .B(\stack[3][53] ), .Z(n15415) );
  NANDN U15854 ( .A(n17472), .B(\stack[5][53] ), .Z(n15414) );
  AND U15855 ( .A(n15415), .B(n15414), .Z(n15417) );
  NANDN U15856 ( .A(n17475), .B(\stack[4][53] ), .Z(n15416) );
  NAND U15857 ( .A(n15417), .B(n15416), .Z(n2210) );
  NANDN U15858 ( .A(n2967), .B(\stack[2][53] ), .Z(n15419) );
  NANDN U15859 ( .A(n17472), .B(\stack[4][53] ), .Z(n15418) );
  AND U15860 ( .A(n15419), .B(n15418), .Z(n15421) );
  NANDN U15861 ( .A(n17475), .B(\stack[3][53] ), .Z(n15420) );
  NAND U15862 ( .A(n15421), .B(n15420), .Z(n2211) );
  NANDN U15863 ( .A(n2967), .B(\stack[1][53] ), .Z(n15423) );
  NANDN U15864 ( .A(n17472), .B(\stack[3][53] ), .Z(n15422) );
  AND U15865 ( .A(n15423), .B(n15422), .Z(n15425) );
  NANDN U15866 ( .A(n17475), .B(\stack[2][53] ), .Z(n15424) );
  NAND U15867 ( .A(n15425), .B(n15424), .Z(n2212) );
  NANDN U15868 ( .A(n2967), .B(o[53]), .Z(n15427) );
  NANDN U15869 ( .A(n17472), .B(\stack[2][53] ), .Z(n15426) );
  AND U15870 ( .A(n15427), .B(n15426), .Z(n15429) );
  NANDN U15871 ( .A(n17475), .B(\stack[1][53] ), .Z(n15428) );
  NAND U15872 ( .A(n15429), .B(n15428), .Z(n2213) );
  NAND U15873 ( .A(\stack[1][53] ), .B(n17479), .Z(n15430) );
  NANDN U15874 ( .A(n17467), .B(n15430), .Z(n15431) );
  AND U15875 ( .A(n15431), .B(o[53]), .Z(n15440) );
  XNOR U15876 ( .A(n15433), .B(n15432), .Z(n15434) );
  NAND U15877 ( .A(n15434), .B(n17458), .Z(n15438) );
  NANDN U15878 ( .A(n2967), .B(x[53]), .Z(n15436) );
  NANDN U15879 ( .A(n17483), .B(\stack[1][53] ), .Z(n15435) );
  AND U15880 ( .A(n15436), .B(n15435), .Z(n15437) );
  NAND U15881 ( .A(n15438), .B(n15437), .Z(n15439) );
  NOR U15882 ( .A(n15440), .B(n15439), .Z(n15441) );
  NANDN U15883 ( .A(n2967), .B(\stack[6][52] ), .Z(n15443) );
  NANDN U15884 ( .A(n17471), .B(\stack[7][52] ), .Z(n15442) );
  NAND U15885 ( .A(n15443), .B(n15442), .Z(n2215) );
  NANDN U15886 ( .A(n2967), .B(\stack[5][52] ), .Z(n15445) );
  NANDN U15887 ( .A(n17472), .B(\stack[7][52] ), .Z(n15444) );
  AND U15888 ( .A(n15445), .B(n15444), .Z(n15447) );
  NANDN U15889 ( .A(n17475), .B(\stack[6][52] ), .Z(n15446) );
  NAND U15890 ( .A(n15447), .B(n15446), .Z(n2216) );
  NANDN U15891 ( .A(n2967), .B(\stack[4][52] ), .Z(n15449) );
  NANDN U15892 ( .A(n17472), .B(\stack[6][52] ), .Z(n15448) );
  AND U15893 ( .A(n15449), .B(n15448), .Z(n15451) );
  NANDN U15894 ( .A(n17475), .B(\stack[5][52] ), .Z(n15450) );
  NAND U15895 ( .A(n15451), .B(n15450), .Z(n2217) );
  NANDN U15896 ( .A(n2967), .B(\stack[3][52] ), .Z(n15453) );
  NANDN U15897 ( .A(n17472), .B(\stack[5][52] ), .Z(n15452) );
  AND U15898 ( .A(n15453), .B(n15452), .Z(n15455) );
  NANDN U15899 ( .A(n17475), .B(\stack[4][52] ), .Z(n15454) );
  NAND U15900 ( .A(n15455), .B(n15454), .Z(n2218) );
  NANDN U15901 ( .A(n2967), .B(\stack[2][52] ), .Z(n15457) );
  NANDN U15902 ( .A(n17472), .B(\stack[4][52] ), .Z(n15456) );
  AND U15903 ( .A(n15457), .B(n15456), .Z(n15459) );
  NANDN U15904 ( .A(n17475), .B(\stack[3][52] ), .Z(n15458) );
  NAND U15905 ( .A(n15459), .B(n15458), .Z(n2219) );
  NANDN U15906 ( .A(n15468), .B(n17471), .Z(n15461) );
  NANDN U15907 ( .A(n17472), .B(\stack[3][52] ), .Z(n15460) );
  AND U15908 ( .A(n15461), .B(n15460), .Z(n15463) );
  NANDN U15909 ( .A(n17475), .B(\stack[2][52] ), .Z(n15462) );
  NAND U15910 ( .A(n15463), .B(n15462), .Z(n2220) );
  NANDN U15911 ( .A(n2967), .B(o[52]), .Z(n15465) );
  NANDN U15912 ( .A(n17472), .B(\stack[2][52] ), .Z(n15464) );
  AND U15913 ( .A(n15465), .B(n15464), .Z(n15467) );
  OR U15914 ( .A(n17475), .B(n15468), .Z(n15466) );
  NAND U15915 ( .A(n15467), .B(n15466), .Z(n2221) );
  NANDN U15916 ( .A(n15468), .B(n17479), .Z(n15469) );
  NANDN U15917 ( .A(n17467), .B(n15469), .Z(n15470) );
  AND U15918 ( .A(n15470), .B(o[52]), .Z(n15479) );
  XNOR U15919 ( .A(n15472), .B(n15471), .Z(n15473) );
  NAND U15920 ( .A(n15473), .B(n17458), .Z(n15477) );
  NANDN U15921 ( .A(n2967), .B(x[52]), .Z(n15475) );
  NANDN U15922 ( .A(n17483), .B(\stack[1][52] ), .Z(n15474) );
  AND U15923 ( .A(n15475), .B(n15474), .Z(n15476) );
  NAND U15924 ( .A(n15477), .B(n15476), .Z(n15478) );
  NOR U15925 ( .A(n15479), .B(n15478), .Z(n15480) );
  NANDN U15926 ( .A(n2967), .B(\stack[6][51] ), .Z(n15482) );
  NANDN U15927 ( .A(n17471), .B(\stack[7][51] ), .Z(n15481) );
  NAND U15928 ( .A(n15482), .B(n15481), .Z(n2223) );
  NANDN U15929 ( .A(n2967), .B(\stack[5][51] ), .Z(n15484) );
  NANDN U15930 ( .A(n17472), .B(\stack[7][51] ), .Z(n15483) );
  AND U15931 ( .A(n15484), .B(n15483), .Z(n15486) );
  NANDN U15932 ( .A(n17475), .B(\stack[6][51] ), .Z(n15485) );
  NAND U15933 ( .A(n15486), .B(n15485), .Z(n2224) );
  NANDN U15934 ( .A(n2967), .B(\stack[4][51] ), .Z(n15488) );
  NANDN U15935 ( .A(n17472), .B(\stack[6][51] ), .Z(n15487) );
  AND U15936 ( .A(n15488), .B(n15487), .Z(n15490) );
  NANDN U15937 ( .A(n17475), .B(\stack[5][51] ), .Z(n15489) );
  NAND U15938 ( .A(n15490), .B(n15489), .Z(n2225) );
  NANDN U15939 ( .A(n2967), .B(\stack[3][51] ), .Z(n15492) );
  NANDN U15940 ( .A(n17472), .B(\stack[5][51] ), .Z(n15491) );
  AND U15941 ( .A(n15492), .B(n15491), .Z(n15494) );
  NANDN U15942 ( .A(n17475), .B(\stack[4][51] ), .Z(n15493) );
  NAND U15943 ( .A(n15494), .B(n15493), .Z(n2226) );
  NANDN U15944 ( .A(n2967), .B(\stack[2][51] ), .Z(n15496) );
  NANDN U15945 ( .A(n17472), .B(\stack[4][51] ), .Z(n15495) );
  AND U15946 ( .A(n15496), .B(n15495), .Z(n15498) );
  NANDN U15947 ( .A(n17475), .B(\stack[3][51] ), .Z(n15497) );
  NAND U15948 ( .A(n15498), .B(n15497), .Z(n2227) );
  NANDN U15949 ( .A(n15507), .B(n17471), .Z(n15500) );
  NANDN U15950 ( .A(n17472), .B(\stack[3][51] ), .Z(n15499) );
  AND U15951 ( .A(n15500), .B(n15499), .Z(n15502) );
  NANDN U15952 ( .A(n17475), .B(\stack[2][51] ), .Z(n15501) );
  NAND U15953 ( .A(n15502), .B(n15501), .Z(n2228) );
  NANDN U15954 ( .A(n2967), .B(o[51]), .Z(n15504) );
  NANDN U15955 ( .A(n17472), .B(\stack[2][51] ), .Z(n15503) );
  AND U15956 ( .A(n15504), .B(n15503), .Z(n15506) );
  OR U15957 ( .A(n17475), .B(n15507), .Z(n15505) );
  NAND U15958 ( .A(n15506), .B(n15505), .Z(n2229) );
  NANDN U15959 ( .A(n15507), .B(n17479), .Z(n15508) );
  NANDN U15960 ( .A(n17467), .B(n15508), .Z(n15509) );
  AND U15961 ( .A(n15509), .B(o[51]), .Z(n15518) );
  XNOR U15962 ( .A(n15511), .B(n15510), .Z(n15512) );
  NAND U15963 ( .A(n15512), .B(n17458), .Z(n15516) );
  NANDN U15964 ( .A(n2967), .B(x[51]), .Z(n15514) );
  NANDN U15965 ( .A(n17483), .B(\stack[1][51] ), .Z(n15513) );
  AND U15966 ( .A(n15514), .B(n15513), .Z(n15515) );
  NAND U15967 ( .A(n15516), .B(n15515), .Z(n15517) );
  NOR U15968 ( .A(n15518), .B(n15517), .Z(n15519) );
  NANDN U15969 ( .A(n2967), .B(\stack[6][50] ), .Z(n15521) );
  NANDN U15970 ( .A(n17471), .B(\stack[7][50] ), .Z(n15520) );
  NAND U15971 ( .A(n15521), .B(n15520), .Z(n2231) );
  NANDN U15972 ( .A(n2967), .B(\stack[5][50] ), .Z(n15523) );
  NANDN U15973 ( .A(n17472), .B(\stack[7][50] ), .Z(n15522) );
  AND U15974 ( .A(n15523), .B(n15522), .Z(n15525) );
  NANDN U15975 ( .A(n17475), .B(\stack[6][50] ), .Z(n15524) );
  NAND U15976 ( .A(n15525), .B(n15524), .Z(n2232) );
  NANDN U15977 ( .A(n2967), .B(\stack[4][50] ), .Z(n15527) );
  NANDN U15978 ( .A(n17472), .B(\stack[6][50] ), .Z(n15526) );
  AND U15979 ( .A(n15527), .B(n15526), .Z(n15529) );
  NANDN U15980 ( .A(n17475), .B(\stack[5][50] ), .Z(n15528) );
  NAND U15981 ( .A(n15529), .B(n15528), .Z(n2233) );
  NANDN U15982 ( .A(n2967), .B(\stack[3][50] ), .Z(n15531) );
  NANDN U15983 ( .A(n17472), .B(\stack[5][50] ), .Z(n15530) );
  AND U15984 ( .A(n15531), .B(n15530), .Z(n15533) );
  NANDN U15985 ( .A(n17475), .B(\stack[4][50] ), .Z(n15532) );
  NAND U15986 ( .A(n15533), .B(n15532), .Z(n2234) );
  NANDN U15987 ( .A(n2967), .B(\stack[2][50] ), .Z(n15535) );
  NANDN U15988 ( .A(n17472), .B(\stack[4][50] ), .Z(n15534) );
  AND U15989 ( .A(n15535), .B(n15534), .Z(n15537) );
  NANDN U15990 ( .A(n17475), .B(\stack[3][50] ), .Z(n15536) );
  NAND U15991 ( .A(n15537), .B(n15536), .Z(n2235) );
  NANDN U15992 ( .A(n15546), .B(n17471), .Z(n15539) );
  NANDN U15993 ( .A(n17472), .B(\stack[3][50] ), .Z(n15538) );
  AND U15994 ( .A(n15539), .B(n15538), .Z(n15541) );
  NANDN U15995 ( .A(n17475), .B(\stack[2][50] ), .Z(n15540) );
  NAND U15996 ( .A(n15541), .B(n15540), .Z(n2236) );
  NANDN U15997 ( .A(n2967), .B(o[50]), .Z(n15543) );
  NANDN U15998 ( .A(n17472), .B(\stack[2][50] ), .Z(n15542) );
  AND U15999 ( .A(n15543), .B(n15542), .Z(n15545) );
  OR U16000 ( .A(n17475), .B(n15546), .Z(n15544) );
  NAND U16001 ( .A(n15545), .B(n15544), .Z(n2237) );
  NANDN U16002 ( .A(n15546), .B(n17479), .Z(n15547) );
  NANDN U16003 ( .A(n17467), .B(n15547), .Z(n15548) );
  AND U16004 ( .A(n15548), .B(o[50]), .Z(n15557) );
  XNOR U16005 ( .A(n15550), .B(n15549), .Z(n15551) );
  NAND U16006 ( .A(n15551), .B(n17458), .Z(n15555) );
  NANDN U16007 ( .A(n2967), .B(x[50]), .Z(n15553) );
  NANDN U16008 ( .A(n17483), .B(\stack[1][50] ), .Z(n15552) );
  AND U16009 ( .A(n15553), .B(n15552), .Z(n15554) );
  NAND U16010 ( .A(n15555), .B(n15554), .Z(n15556) );
  NOR U16011 ( .A(n15557), .B(n15556), .Z(n15558) );
  NANDN U16012 ( .A(n2967), .B(\stack[6][49] ), .Z(n15560) );
  NANDN U16013 ( .A(n17471), .B(\stack[7][49] ), .Z(n15559) );
  NAND U16014 ( .A(n15560), .B(n15559), .Z(n2239) );
  NANDN U16015 ( .A(n2967), .B(\stack[5][49] ), .Z(n15562) );
  NANDN U16016 ( .A(n17472), .B(\stack[7][49] ), .Z(n15561) );
  AND U16017 ( .A(n15562), .B(n15561), .Z(n15564) );
  NANDN U16018 ( .A(n17475), .B(\stack[6][49] ), .Z(n15563) );
  NAND U16019 ( .A(n15564), .B(n15563), .Z(n2240) );
  NANDN U16020 ( .A(n2967), .B(\stack[4][49] ), .Z(n15566) );
  NANDN U16021 ( .A(n17472), .B(\stack[6][49] ), .Z(n15565) );
  AND U16022 ( .A(n15566), .B(n15565), .Z(n15568) );
  NANDN U16023 ( .A(n17475), .B(\stack[5][49] ), .Z(n15567) );
  NAND U16024 ( .A(n15568), .B(n15567), .Z(n2241) );
  NANDN U16025 ( .A(n2967), .B(\stack[3][49] ), .Z(n15570) );
  NANDN U16026 ( .A(n17472), .B(\stack[5][49] ), .Z(n15569) );
  AND U16027 ( .A(n15570), .B(n15569), .Z(n15572) );
  NANDN U16028 ( .A(n17475), .B(\stack[4][49] ), .Z(n15571) );
  NAND U16029 ( .A(n15572), .B(n15571), .Z(n2242) );
  NANDN U16030 ( .A(n2967), .B(\stack[2][49] ), .Z(n15574) );
  NANDN U16031 ( .A(n17472), .B(\stack[4][49] ), .Z(n15573) );
  AND U16032 ( .A(n15574), .B(n15573), .Z(n15576) );
  NANDN U16033 ( .A(n17475), .B(\stack[3][49] ), .Z(n15575) );
  NAND U16034 ( .A(n15576), .B(n15575), .Z(n2243) );
  NANDN U16035 ( .A(n2967), .B(\stack[1][49] ), .Z(n15578) );
  NANDN U16036 ( .A(n17472), .B(\stack[3][49] ), .Z(n15577) );
  AND U16037 ( .A(n15578), .B(n15577), .Z(n15580) );
  NANDN U16038 ( .A(n17475), .B(\stack[2][49] ), .Z(n15579) );
  NAND U16039 ( .A(n15580), .B(n15579), .Z(n2244) );
  NANDN U16040 ( .A(n2967), .B(o[49]), .Z(n15582) );
  NANDN U16041 ( .A(n17472), .B(\stack[2][49] ), .Z(n15581) );
  AND U16042 ( .A(n15582), .B(n15581), .Z(n15584) );
  NANDN U16043 ( .A(n17475), .B(\stack[1][49] ), .Z(n15583) );
  NAND U16044 ( .A(n15584), .B(n15583), .Z(n2245) );
  NAND U16045 ( .A(\stack[1][49] ), .B(n17479), .Z(n15585) );
  NANDN U16046 ( .A(n17467), .B(n15585), .Z(n15586) );
  AND U16047 ( .A(n15586), .B(o[49]), .Z(n15595) );
  XNOR U16048 ( .A(n15588), .B(n15587), .Z(n15589) );
  NAND U16049 ( .A(n15589), .B(n17458), .Z(n15593) );
  NANDN U16050 ( .A(n2967), .B(x[49]), .Z(n15591) );
  NANDN U16051 ( .A(n17483), .B(\stack[1][49] ), .Z(n15590) );
  AND U16052 ( .A(n15591), .B(n15590), .Z(n15592) );
  NAND U16053 ( .A(n15593), .B(n15592), .Z(n15594) );
  NOR U16054 ( .A(n15595), .B(n15594), .Z(n15596) );
  NANDN U16055 ( .A(n2967), .B(\stack[6][48] ), .Z(n15598) );
  NANDN U16056 ( .A(n17471), .B(\stack[7][48] ), .Z(n15597) );
  NAND U16057 ( .A(n15598), .B(n15597), .Z(n2247) );
  NANDN U16058 ( .A(n2967), .B(\stack[5][48] ), .Z(n15600) );
  NANDN U16059 ( .A(n17472), .B(\stack[7][48] ), .Z(n15599) );
  AND U16060 ( .A(n15600), .B(n15599), .Z(n15602) );
  NANDN U16061 ( .A(n17475), .B(\stack[6][48] ), .Z(n15601) );
  NAND U16062 ( .A(n15602), .B(n15601), .Z(n2248) );
  NANDN U16063 ( .A(n2967), .B(\stack[4][48] ), .Z(n15604) );
  NANDN U16064 ( .A(n17472), .B(\stack[6][48] ), .Z(n15603) );
  AND U16065 ( .A(n15604), .B(n15603), .Z(n15606) );
  NANDN U16066 ( .A(n17475), .B(\stack[5][48] ), .Z(n15605) );
  NAND U16067 ( .A(n15606), .B(n15605), .Z(n2249) );
  NANDN U16068 ( .A(n2967), .B(\stack[3][48] ), .Z(n15608) );
  NANDN U16069 ( .A(n17472), .B(\stack[5][48] ), .Z(n15607) );
  AND U16070 ( .A(n15608), .B(n15607), .Z(n15610) );
  NANDN U16071 ( .A(n17475), .B(\stack[4][48] ), .Z(n15609) );
  NAND U16072 ( .A(n15610), .B(n15609), .Z(n2250) );
  NANDN U16073 ( .A(n2967), .B(\stack[2][48] ), .Z(n15612) );
  NANDN U16074 ( .A(n17472), .B(\stack[4][48] ), .Z(n15611) );
  AND U16075 ( .A(n15612), .B(n15611), .Z(n15614) );
  NANDN U16076 ( .A(n17475), .B(\stack[3][48] ), .Z(n15613) );
  NAND U16077 ( .A(n15614), .B(n15613), .Z(n2251) );
  NANDN U16078 ( .A(n15623), .B(n17471), .Z(n15616) );
  NANDN U16079 ( .A(n17472), .B(\stack[3][48] ), .Z(n15615) );
  AND U16080 ( .A(n15616), .B(n15615), .Z(n15618) );
  NANDN U16081 ( .A(n17475), .B(\stack[2][48] ), .Z(n15617) );
  NAND U16082 ( .A(n15618), .B(n15617), .Z(n2252) );
  NANDN U16083 ( .A(n2967), .B(o[48]), .Z(n15620) );
  NANDN U16084 ( .A(n17472), .B(\stack[2][48] ), .Z(n15619) );
  AND U16085 ( .A(n15620), .B(n15619), .Z(n15622) );
  OR U16086 ( .A(n17475), .B(n15623), .Z(n15621) );
  NAND U16087 ( .A(n15622), .B(n15621), .Z(n2253) );
  NANDN U16088 ( .A(n15623), .B(n17479), .Z(n15624) );
  NANDN U16089 ( .A(n17467), .B(n15624), .Z(n15625) );
  AND U16090 ( .A(n15625), .B(o[48]), .Z(n15634) );
  XNOR U16091 ( .A(n15627), .B(n15626), .Z(n15628) );
  NAND U16092 ( .A(n15628), .B(n17458), .Z(n15632) );
  NANDN U16093 ( .A(n2967), .B(x[48]), .Z(n15630) );
  NANDN U16094 ( .A(n17483), .B(\stack[1][48] ), .Z(n15629) );
  AND U16095 ( .A(n15630), .B(n15629), .Z(n15631) );
  NAND U16096 ( .A(n15632), .B(n15631), .Z(n15633) );
  NOR U16097 ( .A(n15634), .B(n15633), .Z(n15635) );
  NANDN U16098 ( .A(n2967), .B(\stack[6][47] ), .Z(n15637) );
  NANDN U16099 ( .A(n17471), .B(\stack[7][47] ), .Z(n15636) );
  NAND U16100 ( .A(n15637), .B(n15636), .Z(n2255) );
  NANDN U16101 ( .A(n2967), .B(\stack[5][47] ), .Z(n15639) );
  NANDN U16102 ( .A(n17472), .B(\stack[7][47] ), .Z(n15638) );
  AND U16103 ( .A(n15639), .B(n15638), .Z(n15641) );
  NANDN U16104 ( .A(n17475), .B(\stack[6][47] ), .Z(n15640) );
  NAND U16105 ( .A(n15641), .B(n15640), .Z(n2256) );
  NANDN U16106 ( .A(n2967), .B(\stack[4][47] ), .Z(n15643) );
  NANDN U16107 ( .A(n17472), .B(\stack[6][47] ), .Z(n15642) );
  AND U16108 ( .A(n15643), .B(n15642), .Z(n15645) );
  NANDN U16109 ( .A(n17475), .B(\stack[5][47] ), .Z(n15644) );
  NAND U16110 ( .A(n15645), .B(n15644), .Z(n2257) );
  NANDN U16111 ( .A(n2967), .B(\stack[3][47] ), .Z(n15647) );
  NANDN U16112 ( .A(n17472), .B(\stack[5][47] ), .Z(n15646) );
  AND U16113 ( .A(n15647), .B(n15646), .Z(n15649) );
  NANDN U16114 ( .A(n17475), .B(\stack[4][47] ), .Z(n15648) );
  NAND U16115 ( .A(n15649), .B(n15648), .Z(n2258) );
  NANDN U16116 ( .A(n2967), .B(\stack[2][47] ), .Z(n15651) );
  NANDN U16117 ( .A(n17472), .B(\stack[4][47] ), .Z(n15650) );
  AND U16118 ( .A(n15651), .B(n15650), .Z(n15653) );
  NANDN U16119 ( .A(n17475), .B(\stack[3][47] ), .Z(n15652) );
  NAND U16120 ( .A(n15653), .B(n15652), .Z(n2259) );
  NANDN U16121 ( .A(n15662), .B(n17471), .Z(n15655) );
  NANDN U16122 ( .A(n17472), .B(\stack[3][47] ), .Z(n15654) );
  AND U16123 ( .A(n15655), .B(n15654), .Z(n15657) );
  NANDN U16124 ( .A(n17475), .B(\stack[2][47] ), .Z(n15656) );
  NAND U16125 ( .A(n15657), .B(n15656), .Z(n2260) );
  NANDN U16126 ( .A(n2967), .B(o[47]), .Z(n15659) );
  NANDN U16127 ( .A(n17472), .B(\stack[2][47] ), .Z(n15658) );
  AND U16128 ( .A(n15659), .B(n15658), .Z(n15661) );
  OR U16129 ( .A(n17475), .B(n15662), .Z(n15660) );
  NAND U16130 ( .A(n15661), .B(n15660), .Z(n2261) );
  NANDN U16131 ( .A(n15662), .B(n17479), .Z(n15663) );
  NANDN U16132 ( .A(n17467), .B(n15663), .Z(n15664) );
  AND U16133 ( .A(n15664), .B(o[47]), .Z(n15673) );
  XNOR U16134 ( .A(n15666), .B(n15665), .Z(n15667) );
  NAND U16135 ( .A(n15667), .B(n17458), .Z(n15671) );
  NANDN U16136 ( .A(n2967), .B(x[47]), .Z(n15669) );
  NANDN U16137 ( .A(n17483), .B(\stack[1][47] ), .Z(n15668) );
  AND U16138 ( .A(n15669), .B(n15668), .Z(n15670) );
  NAND U16139 ( .A(n15671), .B(n15670), .Z(n15672) );
  NOR U16140 ( .A(n15673), .B(n15672), .Z(n15674) );
  NANDN U16141 ( .A(n2967), .B(\stack[6][46] ), .Z(n15676) );
  NANDN U16142 ( .A(n17471), .B(\stack[7][46] ), .Z(n15675) );
  NAND U16143 ( .A(n15676), .B(n15675), .Z(n2263) );
  NANDN U16144 ( .A(n2967), .B(\stack[5][46] ), .Z(n15678) );
  NANDN U16145 ( .A(n17472), .B(\stack[7][46] ), .Z(n15677) );
  AND U16146 ( .A(n15678), .B(n15677), .Z(n15680) );
  NANDN U16147 ( .A(n17475), .B(\stack[6][46] ), .Z(n15679) );
  NAND U16148 ( .A(n15680), .B(n15679), .Z(n2264) );
  NANDN U16149 ( .A(n2967), .B(\stack[4][46] ), .Z(n15682) );
  NANDN U16150 ( .A(n17472), .B(\stack[6][46] ), .Z(n15681) );
  AND U16151 ( .A(n15682), .B(n15681), .Z(n15684) );
  NANDN U16152 ( .A(n17475), .B(\stack[5][46] ), .Z(n15683) );
  NAND U16153 ( .A(n15684), .B(n15683), .Z(n2265) );
  NANDN U16154 ( .A(n2967), .B(\stack[3][46] ), .Z(n15686) );
  NANDN U16155 ( .A(n17472), .B(\stack[5][46] ), .Z(n15685) );
  AND U16156 ( .A(n15686), .B(n15685), .Z(n15688) );
  NANDN U16157 ( .A(n17475), .B(\stack[4][46] ), .Z(n15687) );
  NAND U16158 ( .A(n15688), .B(n15687), .Z(n2266) );
  NANDN U16159 ( .A(n2967), .B(\stack[2][46] ), .Z(n15690) );
  NANDN U16160 ( .A(n17472), .B(\stack[4][46] ), .Z(n15689) );
  AND U16161 ( .A(n15690), .B(n15689), .Z(n15692) );
  NANDN U16162 ( .A(n17475), .B(\stack[3][46] ), .Z(n15691) );
  NAND U16163 ( .A(n15692), .B(n15691), .Z(n2267) );
  NANDN U16164 ( .A(n15701), .B(n17471), .Z(n15694) );
  NANDN U16165 ( .A(n17472), .B(\stack[3][46] ), .Z(n15693) );
  AND U16166 ( .A(n15694), .B(n15693), .Z(n15696) );
  NANDN U16167 ( .A(n17475), .B(\stack[2][46] ), .Z(n15695) );
  NAND U16168 ( .A(n15696), .B(n15695), .Z(n2268) );
  NANDN U16169 ( .A(n2967), .B(o[46]), .Z(n15698) );
  NANDN U16170 ( .A(n17472), .B(\stack[2][46] ), .Z(n15697) );
  AND U16171 ( .A(n15698), .B(n15697), .Z(n15700) );
  OR U16172 ( .A(n17475), .B(n15701), .Z(n15699) );
  NAND U16173 ( .A(n15700), .B(n15699), .Z(n2269) );
  NANDN U16174 ( .A(n15701), .B(n17479), .Z(n15702) );
  NANDN U16175 ( .A(n17467), .B(n15702), .Z(n15703) );
  AND U16176 ( .A(n15703), .B(o[46]), .Z(n15712) );
  XNOR U16177 ( .A(n15705), .B(n15704), .Z(n15706) );
  NAND U16178 ( .A(n15706), .B(n17458), .Z(n15710) );
  NANDN U16179 ( .A(n2967), .B(x[46]), .Z(n15708) );
  NANDN U16180 ( .A(n17483), .B(\stack[1][46] ), .Z(n15707) );
  AND U16181 ( .A(n15708), .B(n15707), .Z(n15709) );
  NAND U16182 ( .A(n15710), .B(n15709), .Z(n15711) );
  NOR U16183 ( .A(n15712), .B(n15711), .Z(n15713) );
  NANDN U16184 ( .A(n2967), .B(\stack[6][45] ), .Z(n15715) );
  NANDN U16185 ( .A(n17471), .B(\stack[7][45] ), .Z(n15714) );
  NAND U16186 ( .A(n15715), .B(n15714), .Z(n2271) );
  NANDN U16187 ( .A(n2967), .B(\stack[5][45] ), .Z(n15717) );
  NANDN U16188 ( .A(n17472), .B(\stack[7][45] ), .Z(n15716) );
  AND U16189 ( .A(n15717), .B(n15716), .Z(n15719) );
  NANDN U16190 ( .A(n17475), .B(\stack[6][45] ), .Z(n15718) );
  NAND U16191 ( .A(n15719), .B(n15718), .Z(n2272) );
  NANDN U16192 ( .A(n2967), .B(\stack[4][45] ), .Z(n15721) );
  NANDN U16193 ( .A(n17472), .B(\stack[6][45] ), .Z(n15720) );
  AND U16194 ( .A(n15721), .B(n15720), .Z(n15723) );
  NANDN U16195 ( .A(n17475), .B(\stack[5][45] ), .Z(n15722) );
  NAND U16196 ( .A(n15723), .B(n15722), .Z(n2273) );
  NANDN U16197 ( .A(n2967), .B(\stack[3][45] ), .Z(n15725) );
  NANDN U16198 ( .A(n17472), .B(\stack[5][45] ), .Z(n15724) );
  AND U16199 ( .A(n15725), .B(n15724), .Z(n15727) );
  NANDN U16200 ( .A(n17475), .B(\stack[4][45] ), .Z(n15726) );
  NAND U16201 ( .A(n15727), .B(n15726), .Z(n2274) );
  NANDN U16202 ( .A(n2967), .B(\stack[2][45] ), .Z(n15729) );
  NANDN U16203 ( .A(n17472), .B(\stack[4][45] ), .Z(n15728) );
  AND U16204 ( .A(n15729), .B(n15728), .Z(n15731) );
  NANDN U16205 ( .A(n17475), .B(\stack[3][45] ), .Z(n15730) );
  NAND U16206 ( .A(n15731), .B(n15730), .Z(n2275) );
  NANDN U16207 ( .A(n15740), .B(n17471), .Z(n15733) );
  NANDN U16208 ( .A(n17472), .B(\stack[3][45] ), .Z(n15732) );
  AND U16209 ( .A(n15733), .B(n15732), .Z(n15735) );
  NANDN U16210 ( .A(n17475), .B(\stack[2][45] ), .Z(n15734) );
  NAND U16211 ( .A(n15735), .B(n15734), .Z(n2276) );
  NANDN U16212 ( .A(n2967), .B(o[45]), .Z(n15737) );
  NANDN U16213 ( .A(n17472), .B(\stack[2][45] ), .Z(n15736) );
  AND U16214 ( .A(n15737), .B(n15736), .Z(n15739) );
  OR U16215 ( .A(n17475), .B(n15740), .Z(n15738) );
  NAND U16216 ( .A(n15739), .B(n15738), .Z(n2277) );
  NANDN U16217 ( .A(n15740), .B(n17479), .Z(n15741) );
  NANDN U16218 ( .A(n17467), .B(n15741), .Z(n15742) );
  AND U16219 ( .A(n15742), .B(o[45]), .Z(n15751) );
  XNOR U16220 ( .A(n15744), .B(n15743), .Z(n15745) );
  NAND U16221 ( .A(n15745), .B(n17458), .Z(n15749) );
  NANDN U16222 ( .A(n2967), .B(x[45]), .Z(n15747) );
  NANDN U16223 ( .A(n17483), .B(\stack[1][45] ), .Z(n15746) );
  AND U16224 ( .A(n15747), .B(n15746), .Z(n15748) );
  NAND U16225 ( .A(n15749), .B(n15748), .Z(n15750) );
  NOR U16226 ( .A(n15751), .B(n15750), .Z(n15752) );
  NANDN U16227 ( .A(n2967), .B(\stack[6][44] ), .Z(n15754) );
  NANDN U16228 ( .A(n17471), .B(\stack[7][44] ), .Z(n15753) );
  NAND U16229 ( .A(n15754), .B(n15753), .Z(n2279) );
  NANDN U16230 ( .A(n2967), .B(\stack[5][44] ), .Z(n15756) );
  NANDN U16231 ( .A(n17472), .B(\stack[7][44] ), .Z(n15755) );
  AND U16232 ( .A(n15756), .B(n15755), .Z(n15758) );
  NANDN U16233 ( .A(n17475), .B(\stack[6][44] ), .Z(n15757) );
  NAND U16234 ( .A(n15758), .B(n15757), .Z(n2280) );
  NANDN U16235 ( .A(n2967), .B(\stack[4][44] ), .Z(n15760) );
  NANDN U16236 ( .A(n17472), .B(\stack[6][44] ), .Z(n15759) );
  AND U16237 ( .A(n15760), .B(n15759), .Z(n15762) );
  NANDN U16238 ( .A(n17475), .B(\stack[5][44] ), .Z(n15761) );
  NAND U16239 ( .A(n15762), .B(n15761), .Z(n2281) );
  NANDN U16240 ( .A(n2967), .B(\stack[3][44] ), .Z(n15764) );
  NANDN U16241 ( .A(n17472), .B(\stack[5][44] ), .Z(n15763) );
  AND U16242 ( .A(n15764), .B(n15763), .Z(n15766) );
  NANDN U16243 ( .A(n17475), .B(\stack[4][44] ), .Z(n15765) );
  NAND U16244 ( .A(n15766), .B(n15765), .Z(n2282) );
  NANDN U16245 ( .A(n2967), .B(\stack[2][44] ), .Z(n15768) );
  NANDN U16246 ( .A(n17472), .B(\stack[4][44] ), .Z(n15767) );
  AND U16247 ( .A(n15768), .B(n15767), .Z(n15770) );
  NANDN U16248 ( .A(n17475), .B(\stack[3][44] ), .Z(n15769) );
  NAND U16249 ( .A(n15770), .B(n15769), .Z(n2283) );
  NANDN U16250 ( .A(n15779), .B(n17471), .Z(n15772) );
  NANDN U16251 ( .A(n17472), .B(\stack[3][44] ), .Z(n15771) );
  AND U16252 ( .A(n15772), .B(n15771), .Z(n15774) );
  NANDN U16253 ( .A(n17475), .B(\stack[2][44] ), .Z(n15773) );
  NAND U16254 ( .A(n15774), .B(n15773), .Z(n2284) );
  NANDN U16255 ( .A(n2967), .B(o[44]), .Z(n15776) );
  NANDN U16256 ( .A(n17472), .B(\stack[2][44] ), .Z(n15775) );
  AND U16257 ( .A(n15776), .B(n15775), .Z(n15778) );
  OR U16258 ( .A(n17475), .B(n15779), .Z(n15777) );
  NAND U16259 ( .A(n15778), .B(n15777), .Z(n2285) );
  NANDN U16260 ( .A(n15779), .B(n17479), .Z(n15780) );
  NANDN U16261 ( .A(n17467), .B(n15780), .Z(n15781) );
  AND U16262 ( .A(n15781), .B(o[44]), .Z(n15790) );
  XNOR U16263 ( .A(n15783), .B(n15782), .Z(n15784) );
  NAND U16264 ( .A(n15784), .B(n17458), .Z(n15788) );
  NANDN U16265 ( .A(n2967), .B(x[44]), .Z(n15786) );
  NANDN U16266 ( .A(n17483), .B(\stack[1][44] ), .Z(n15785) );
  AND U16267 ( .A(n15786), .B(n15785), .Z(n15787) );
  NAND U16268 ( .A(n15788), .B(n15787), .Z(n15789) );
  NOR U16269 ( .A(n15790), .B(n15789), .Z(n15791) );
  NANDN U16270 ( .A(n2967), .B(\stack[6][43] ), .Z(n15793) );
  NANDN U16271 ( .A(n17471), .B(\stack[7][43] ), .Z(n15792) );
  NAND U16272 ( .A(n15793), .B(n15792), .Z(n2287) );
  NANDN U16273 ( .A(n2967), .B(\stack[5][43] ), .Z(n15795) );
  NANDN U16274 ( .A(n17472), .B(\stack[7][43] ), .Z(n15794) );
  AND U16275 ( .A(n15795), .B(n15794), .Z(n15797) );
  NANDN U16276 ( .A(n17475), .B(\stack[6][43] ), .Z(n15796) );
  NAND U16277 ( .A(n15797), .B(n15796), .Z(n2288) );
  NANDN U16278 ( .A(n2967), .B(\stack[4][43] ), .Z(n15799) );
  NANDN U16279 ( .A(n17472), .B(\stack[6][43] ), .Z(n15798) );
  AND U16280 ( .A(n15799), .B(n15798), .Z(n15801) );
  NANDN U16281 ( .A(n17475), .B(\stack[5][43] ), .Z(n15800) );
  NAND U16282 ( .A(n15801), .B(n15800), .Z(n2289) );
  NANDN U16283 ( .A(n2967), .B(\stack[3][43] ), .Z(n15803) );
  NANDN U16284 ( .A(n17472), .B(\stack[5][43] ), .Z(n15802) );
  AND U16285 ( .A(n15803), .B(n15802), .Z(n15805) );
  NANDN U16286 ( .A(n17475), .B(\stack[4][43] ), .Z(n15804) );
  NAND U16287 ( .A(n15805), .B(n15804), .Z(n2290) );
  NANDN U16288 ( .A(n2967), .B(\stack[2][43] ), .Z(n15807) );
  NANDN U16289 ( .A(n17472), .B(\stack[4][43] ), .Z(n15806) );
  AND U16290 ( .A(n15807), .B(n15806), .Z(n15809) );
  NANDN U16291 ( .A(n17475), .B(\stack[3][43] ), .Z(n15808) );
  NAND U16292 ( .A(n15809), .B(n15808), .Z(n2291) );
  NANDN U16293 ( .A(n15818), .B(n17471), .Z(n15811) );
  NANDN U16294 ( .A(n17472), .B(\stack[3][43] ), .Z(n15810) );
  AND U16295 ( .A(n15811), .B(n15810), .Z(n15813) );
  NANDN U16296 ( .A(n17475), .B(\stack[2][43] ), .Z(n15812) );
  NAND U16297 ( .A(n15813), .B(n15812), .Z(n2292) );
  NANDN U16298 ( .A(n2967), .B(o[43]), .Z(n15815) );
  NANDN U16299 ( .A(n17472), .B(\stack[2][43] ), .Z(n15814) );
  AND U16300 ( .A(n15815), .B(n15814), .Z(n15817) );
  OR U16301 ( .A(n17475), .B(n15818), .Z(n15816) );
  NAND U16302 ( .A(n15817), .B(n15816), .Z(n2293) );
  NANDN U16303 ( .A(n15818), .B(n17479), .Z(n15819) );
  NANDN U16304 ( .A(n17467), .B(n15819), .Z(n15820) );
  AND U16305 ( .A(n15820), .B(o[43]), .Z(n15829) );
  XNOR U16306 ( .A(n15822), .B(n15821), .Z(n15823) );
  NAND U16307 ( .A(n15823), .B(n17458), .Z(n15827) );
  NANDN U16308 ( .A(n2967), .B(x[43]), .Z(n15825) );
  NANDN U16309 ( .A(n17483), .B(\stack[1][43] ), .Z(n15824) );
  AND U16310 ( .A(n15825), .B(n15824), .Z(n15826) );
  NAND U16311 ( .A(n15827), .B(n15826), .Z(n15828) );
  NOR U16312 ( .A(n15829), .B(n15828), .Z(n15830) );
  NANDN U16313 ( .A(n2967), .B(\stack[6][42] ), .Z(n15832) );
  NANDN U16314 ( .A(n17471), .B(\stack[7][42] ), .Z(n15831) );
  NAND U16315 ( .A(n15832), .B(n15831), .Z(n2295) );
  NANDN U16316 ( .A(n2967), .B(\stack[5][42] ), .Z(n15834) );
  NANDN U16317 ( .A(n17472), .B(\stack[7][42] ), .Z(n15833) );
  AND U16318 ( .A(n15834), .B(n15833), .Z(n15836) );
  NANDN U16319 ( .A(n17475), .B(\stack[6][42] ), .Z(n15835) );
  NAND U16320 ( .A(n15836), .B(n15835), .Z(n2296) );
  NANDN U16321 ( .A(n2967), .B(\stack[4][42] ), .Z(n15838) );
  NANDN U16322 ( .A(n17472), .B(\stack[6][42] ), .Z(n15837) );
  AND U16323 ( .A(n15838), .B(n15837), .Z(n15840) );
  NANDN U16324 ( .A(n17475), .B(\stack[5][42] ), .Z(n15839) );
  NAND U16325 ( .A(n15840), .B(n15839), .Z(n2297) );
  NANDN U16326 ( .A(n2967), .B(\stack[3][42] ), .Z(n15842) );
  NANDN U16327 ( .A(n17472), .B(\stack[5][42] ), .Z(n15841) );
  AND U16328 ( .A(n15842), .B(n15841), .Z(n15844) );
  NANDN U16329 ( .A(n17475), .B(\stack[4][42] ), .Z(n15843) );
  NAND U16330 ( .A(n15844), .B(n15843), .Z(n2298) );
  NANDN U16331 ( .A(n2967), .B(\stack[2][42] ), .Z(n15846) );
  NANDN U16332 ( .A(n17472), .B(\stack[4][42] ), .Z(n15845) );
  AND U16333 ( .A(n15846), .B(n15845), .Z(n15848) );
  NANDN U16334 ( .A(n17475), .B(\stack[3][42] ), .Z(n15847) );
  NAND U16335 ( .A(n15848), .B(n15847), .Z(n2299) );
  NANDN U16336 ( .A(n15857), .B(n17471), .Z(n15850) );
  NANDN U16337 ( .A(n17472), .B(\stack[3][42] ), .Z(n15849) );
  AND U16338 ( .A(n15850), .B(n15849), .Z(n15852) );
  NANDN U16339 ( .A(n17475), .B(\stack[2][42] ), .Z(n15851) );
  NAND U16340 ( .A(n15852), .B(n15851), .Z(n2300) );
  NANDN U16341 ( .A(n2967), .B(o[42]), .Z(n15854) );
  NANDN U16342 ( .A(n17472), .B(\stack[2][42] ), .Z(n15853) );
  AND U16343 ( .A(n15854), .B(n15853), .Z(n15856) );
  OR U16344 ( .A(n17475), .B(n15857), .Z(n15855) );
  NAND U16345 ( .A(n15856), .B(n15855), .Z(n2301) );
  NANDN U16346 ( .A(n15857), .B(n17479), .Z(n15858) );
  NANDN U16347 ( .A(n17467), .B(n15858), .Z(n15859) );
  AND U16348 ( .A(n15859), .B(o[42]), .Z(n15868) );
  XNOR U16349 ( .A(n15861), .B(n15860), .Z(n15862) );
  NAND U16350 ( .A(n15862), .B(n17458), .Z(n15866) );
  NANDN U16351 ( .A(n2967), .B(x[42]), .Z(n15864) );
  NANDN U16352 ( .A(n17483), .B(\stack[1][42] ), .Z(n15863) );
  AND U16353 ( .A(n15864), .B(n15863), .Z(n15865) );
  NAND U16354 ( .A(n15866), .B(n15865), .Z(n15867) );
  NOR U16355 ( .A(n15868), .B(n15867), .Z(n15869) );
  NANDN U16356 ( .A(n2967), .B(\stack[6][41] ), .Z(n15871) );
  NANDN U16357 ( .A(n17471), .B(\stack[7][41] ), .Z(n15870) );
  NAND U16358 ( .A(n15871), .B(n15870), .Z(n2303) );
  NANDN U16359 ( .A(n2967), .B(\stack[5][41] ), .Z(n15873) );
  NANDN U16360 ( .A(n17472), .B(\stack[7][41] ), .Z(n15872) );
  AND U16361 ( .A(n15873), .B(n15872), .Z(n15875) );
  NANDN U16362 ( .A(n17475), .B(\stack[6][41] ), .Z(n15874) );
  NAND U16363 ( .A(n15875), .B(n15874), .Z(n2304) );
  NANDN U16364 ( .A(n2967), .B(\stack[4][41] ), .Z(n15877) );
  NANDN U16365 ( .A(n17472), .B(\stack[6][41] ), .Z(n15876) );
  AND U16366 ( .A(n15877), .B(n15876), .Z(n15879) );
  NANDN U16367 ( .A(n17475), .B(\stack[5][41] ), .Z(n15878) );
  NAND U16368 ( .A(n15879), .B(n15878), .Z(n2305) );
  NANDN U16369 ( .A(n2967), .B(\stack[3][41] ), .Z(n15881) );
  NANDN U16370 ( .A(n17472), .B(\stack[5][41] ), .Z(n15880) );
  AND U16371 ( .A(n15881), .B(n15880), .Z(n15883) );
  NANDN U16372 ( .A(n17475), .B(\stack[4][41] ), .Z(n15882) );
  NAND U16373 ( .A(n15883), .B(n15882), .Z(n2306) );
  NANDN U16374 ( .A(n2967), .B(\stack[2][41] ), .Z(n15885) );
  NANDN U16375 ( .A(n17472), .B(\stack[4][41] ), .Z(n15884) );
  AND U16376 ( .A(n15885), .B(n15884), .Z(n15887) );
  NANDN U16377 ( .A(n17475), .B(\stack[3][41] ), .Z(n15886) );
  NAND U16378 ( .A(n15887), .B(n15886), .Z(n2307) );
  NANDN U16379 ( .A(n15896), .B(n17471), .Z(n15889) );
  NANDN U16380 ( .A(n17472), .B(\stack[3][41] ), .Z(n15888) );
  AND U16381 ( .A(n15889), .B(n15888), .Z(n15891) );
  NANDN U16382 ( .A(n17475), .B(\stack[2][41] ), .Z(n15890) );
  NAND U16383 ( .A(n15891), .B(n15890), .Z(n2308) );
  NANDN U16384 ( .A(n2967), .B(o[41]), .Z(n15893) );
  NANDN U16385 ( .A(n17472), .B(\stack[2][41] ), .Z(n15892) );
  AND U16386 ( .A(n15893), .B(n15892), .Z(n15895) );
  OR U16387 ( .A(n17475), .B(n15896), .Z(n15894) );
  NAND U16388 ( .A(n15895), .B(n15894), .Z(n2309) );
  NANDN U16389 ( .A(n15896), .B(n17479), .Z(n15897) );
  NANDN U16390 ( .A(n17467), .B(n15897), .Z(n15898) );
  AND U16391 ( .A(n15898), .B(o[41]), .Z(n15907) );
  XNOR U16392 ( .A(n15900), .B(n15899), .Z(n15901) );
  NAND U16393 ( .A(n15901), .B(n17458), .Z(n15905) );
  NANDN U16394 ( .A(n2967), .B(x[41]), .Z(n15903) );
  NANDN U16395 ( .A(n17483), .B(\stack[1][41] ), .Z(n15902) );
  AND U16396 ( .A(n15903), .B(n15902), .Z(n15904) );
  NAND U16397 ( .A(n15905), .B(n15904), .Z(n15906) );
  NOR U16398 ( .A(n15907), .B(n15906), .Z(n15908) );
  NANDN U16399 ( .A(n2967), .B(\stack[6][40] ), .Z(n15910) );
  NANDN U16400 ( .A(n17471), .B(\stack[7][40] ), .Z(n15909) );
  NAND U16401 ( .A(n15910), .B(n15909), .Z(n2311) );
  NANDN U16402 ( .A(n2967), .B(\stack[5][40] ), .Z(n15912) );
  NANDN U16403 ( .A(n17472), .B(\stack[7][40] ), .Z(n15911) );
  AND U16404 ( .A(n15912), .B(n15911), .Z(n15914) );
  NANDN U16405 ( .A(n17475), .B(\stack[6][40] ), .Z(n15913) );
  NAND U16406 ( .A(n15914), .B(n15913), .Z(n2312) );
  NANDN U16407 ( .A(n2967), .B(\stack[4][40] ), .Z(n15916) );
  NANDN U16408 ( .A(n17472), .B(\stack[6][40] ), .Z(n15915) );
  AND U16409 ( .A(n15916), .B(n15915), .Z(n15918) );
  NANDN U16410 ( .A(n17475), .B(\stack[5][40] ), .Z(n15917) );
  NAND U16411 ( .A(n15918), .B(n15917), .Z(n2313) );
  NANDN U16412 ( .A(n2967), .B(\stack[3][40] ), .Z(n15920) );
  NANDN U16413 ( .A(n17472), .B(\stack[5][40] ), .Z(n15919) );
  AND U16414 ( .A(n15920), .B(n15919), .Z(n15922) );
  NANDN U16415 ( .A(n17475), .B(\stack[4][40] ), .Z(n15921) );
  NAND U16416 ( .A(n15922), .B(n15921), .Z(n2314) );
  NANDN U16417 ( .A(n2967), .B(\stack[2][40] ), .Z(n15924) );
  NANDN U16418 ( .A(n17472), .B(\stack[4][40] ), .Z(n15923) );
  AND U16419 ( .A(n15924), .B(n15923), .Z(n15926) );
  NANDN U16420 ( .A(n17475), .B(\stack[3][40] ), .Z(n15925) );
  NAND U16421 ( .A(n15926), .B(n15925), .Z(n2315) );
  NANDN U16422 ( .A(n15935), .B(n17471), .Z(n15928) );
  NANDN U16423 ( .A(n17472), .B(\stack[3][40] ), .Z(n15927) );
  AND U16424 ( .A(n15928), .B(n15927), .Z(n15930) );
  NANDN U16425 ( .A(n17475), .B(\stack[2][40] ), .Z(n15929) );
  NAND U16426 ( .A(n15930), .B(n15929), .Z(n2316) );
  NANDN U16427 ( .A(n2967), .B(o[40]), .Z(n15932) );
  NANDN U16428 ( .A(n17472), .B(\stack[2][40] ), .Z(n15931) );
  AND U16429 ( .A(n15932), .B(n15931), .Z(n15934) );
  OR U16430 ( .A(n17475), .B(n15935), .Z(n15933) );
  NAND U16431 ( .A(n15934), .B(n15933), .Z(n2317) );
  NANDN U16432 ( .A(n15935), .B(n17479), .Z(n15936) );
  NANDN U16433 ( .A(n17467), .B(n15936), .Z(n15937) );
  AND U16434 ( .A(n15937), .B(o[40]), .Z(n15946) );
  XNOR U16435 ( .A(n15939), .B(n15938), .Z(n15940) );
  NAND U16436 ( .A(n15940), .B(n17458), .Z(n15944) );
  NANDN U16437 ( .A(n2967), .B(x[40]), .Z(n15942) );
  NANDN U16438 ( .A(n17483), .B(\stack[1][40] ), .Z(n15941) );
  AND U16439 ( .A(n15942), .B(n15941), .Z(n15943) );
  NAND U16440 ( .A(n15944), .B(n15943), .Z(n15945) );
  NOR U16441 ( .A(n15946), .B(n15945), .Z(n15947) );
  NANDN U16442 ( .A(n2967), .B(\stack[6][39] ), .Z(n15949) );
  NANDN U16443 ( .A(n17471), .B(\stack[7][39] ), .Z(n15948) );
  NAND U16444 ( .A(n15949), .B(n15948), .Z(n2319) );
  NANDN U16445 ( .A(n2967), .B(\stack[5][39] ), .Z(n15951) );
  NANDN U16446 ( .A(n17472), .B(\stack[7][39] ), .Z(n15950) );
  AND U16447 ( .A(n15951), .B(n15950), .Z(n15953) );
  NANDN U16448 ( .A(n17475), .B(\stack[6][39] ), .Z(n15952) );
  NAND U16449 ( .A(n15953), .B(n15952), .Z(n2320) );
  NANDN U16450 ( .A(n2967), .B(\stack[4][39] ), .Z(n15955) );
  NANDN U16451 ( .A(n17472), .B(\stack[6][39] ), .Z(n15954) );
  AND U16452 ( .A(n15955), .B(n15954), .Z(n15957) );
  NANDN U16453 ( .A(n17475), .B(\stack[5][39] ), .Z(n15956) );
  NAND U16454 ( .A(n15957), .B(n15956), .Z(n2321) );
  NANDN U16455 ( .A(n2967), .B(\stack[3][39] ), .Z(n15959) );
  NANDN U16456 ( .A(n17472), .B(\stack[5][39] ), .Z(n15958) );
  AND U16457 ( .A(n15959), .B(n15958), .Z(n15961) );
  NANDN U16458 ( .A(n17475), .B(\stack[4][39] ), .Z(n15960) );
  NAND U16459 ( .A(n15961), .B(n15960), .Z(n2322) );
  NANDN U16460 ( .A(n2967), .B(\stack[2][39] ), .Z(n15963) );
  NANDN U16461 ( .A(n17472), .B(\stack[4][39] ), .Z(n15962) );
  AND U16462 ( .A(n15963), .B(n15962), .Z(n15965) );
  NANDN U16463 ( .A(n17475), .B(\stack[3][39] ), .Z(n15964) );
  NAND U16464 ( .A(n15965), .B(n15964), .Z(n2323) );
  NANDN U16465 ( .A(n2967), .B(\stack[1][39] ), .Z(n15967) );
  NANDN U16466 ( .A(n17472), .B(\stack[3][39] ), .Z(n15966) );
  AND U16467 ( .A(n15967), .B(n15966), .Z(n15969) );
  NANDN U16468 ( .A(n17475), .B(\stack[2][39] ), .Z(n15968) );
  NAND U16469 ( .A(n15969), .B(n15968), .Z(n2324) );
  NANDN U16470 ( .A(n2967), .B(o[39]), .Z(n15971) );
  NANDN U16471 ( .A(n17472), .B(\stack[2][39] ), .Z(n15970) );
  AND U16472 ( .A(n15971), .B(n15970), .Z(n15973) );
  NANDN U16473 ( .A(n17475), .B(\stack[1][39] ), .Z(n15972) );
  NAND U16474 ( .A(n15973), .B(n15972), .Z(n2325) );
  NAND U16475 ( .A(\stack[1][39] ), .B(n17479), .Z(n15974) );
  NANDN U16476 ( .A(n17467), .B(n15974), .Z(n15975) );
  AND U16477 ( .A(n15975), .B(o[39]), .Z(n15984) );
  XNOR U16478 ( .A(n15977), .B(n15976), .Z(n15978) );
  NAND U16479 ( .A(n15978), .B(n17458), .Z(n15982) );
  NANDN U16480 ( .A(n2967), .B(x[39]), .Z(n15980) );
  NANDN U16481 ( .A(n17483), .B(\stack[1][39] ), .Z(n15979) );
  AND U16482 ( .A(n15980), .B(n15979), .Z(n15981) );
  NAND U16483 ( .A(n15982), .B(n15981), .Z(n15983) );
  NOR U16484 ( .A(n15984), .B(n15983), .Z(n15985) );
  NANDN U16485 ( .A(n2967), .B(\stack[6][38] ), .Z(n15987) );
  NANDN U16486 ( .A(n17471), .B(\stack[7][38] ), .Z(n15986) );
  NAND U16487 ( .A(n15987), .B(n15986), .Z(n2327) );
  NANDN U16488 ( .A(n2967), .B(\stack[5][38] ), .Z(n15989) );
  NANDN U16489 ( .A(n17472), .B(\stack[7][38] ), .Z(n15988) );
  AND U16490 ( .A(n15989), .B(n15988), .Z(n15991) );
  NANDN U16491 ( .A(n17475), .B(\stack[6][38] ), .Z(n15990) );
  NAND U16492 ( .A(n15991), .B(n15990), .Z(n2328) );
  NANDN U16493 ( .A(n2967), .B(\stack[4][38] ), .Z(n15993) );
  NANDN U16494 ( .A(n17472), .B(\stack[6][38] ), .Z(n15992) );
  AND U16495 ( .A(n15993), .B(n15992), .Z(n15995) );
  NANDN U16496 ( .A(n17475), .B(\stack[5][38] ), .Z(n15994) );
  NAND U16497 ( .A(n15995), .B(n15994), .Z(n2329) );
  NANDN U16498 ( .A(n2967), .B(\stack[3][38] ), .Z(n15997) );
  NANDN U16499 ( .A(n17472), .B(\stack[5][38] ), .Z(n15996) );
  AND U16500 ( .A(n15997), .B(n15996), .Z(n15999) );
  NANDN U16501 ( .A(n17475), .B(\stack[4][38] ), .Z(n15998) );
  NAND U16502 ( .A(n15999), .B(n15998), .Z(n2330) );
  NANDN U16503 ( .A(n2967), .B(\stack[2][38] ), .Z(n16001) );
  NANDN U16504 ( .A(n17472), .B(\stack[4][38] ), .Z(n16000) );
  AND U16505 ( .A(n16001), .B(n16000), .Z(n16003) );
  NANDN U16506 ( .A(n17475), .B(\stack[3][38] ), .Z(n16002) );
  NAND U16507 ( .A(n16003), .B(n16002), .Z(n2331) );
  NANDN U16508 ( .A(n2967), .B(\stack[1][38] ), .Z(n16005) );
  NANDN U16509 ( .A(n17472), .B(\stack[3][38] ), .Z(n16004) );
  AND U16510 ( .A(n16005), .B(n16004), .Z(n16007) );
  NANDN U16511 ( .A(n17475), .B(\stack[2][38] ), .Z(n16006) );
  NAND U16512 ( .A(n16007), .B(n16006), .Z(n2332) );
  NANDN U16513 ( .A(n2967), .B(o[38]), .Z(n16009) );
  NANDN U16514 ( .A(n17472), .B(\stack[2][38] ), .Z(n16008) );
  AND U16515 ( .A(n16009), .B(n16008), .Z(n16011) );
  NANDN U16516 ( .A(n17475), .B(\stack[1][38] ), .Z(n16010) );
  NAND U16517 ( .A(n16011), .B(n16010), .Z(n2333) );
  NAND U16518 ( .A(\stack[1][38] ), .B(n17479), .Z(n16012) );
  NANDN U16519 ( .A(n17467), .B(n16012), .Z(n16013) );
  AND U16520 ( .A(n16013), .B(o[38]), .Z(n16022) );
  XNOR U16521 ( .A(n16015), .B(n16014), .Z(n16016) );
  NAND U16522 ( .A(n16016), .B(n17458), .Z(n16020) );
  NANDN U16523 ( .A(n2967), .B(x[38]), .Z(n16018) );
  NANDN U16524 ( .A(n17483), .B(\stack[1][38] ), .Z(n16017) );
  AND U16525 ( .A(n16018), .B(n16017), .Z(n16019) );
  NAND U16526 ( .A(n16020), .B(n16019), .Z(n16021) );
  NOR U16527 ( .A(n16022), .B(n16021), .Z(n16023) );
  NANDN U16528 ( .A(n2967), .B(\stack[6][37] ), .Z(n16025) );
  NANDN U16529 ( .A(n17471), .B(\stack[7][37] ), .Z(n16024) );
  NAND U16530 ( .A(n16025), .B(n16024), .Z(n2335) );
  NANDN U16531 ( .A(n2967), .B(\stack[5][37] ), .Z(n16027) );
  NANDN U16532 ( .A(n17472), .B(\stack[7][37] ), .Z(n16026) );
  AND U16533 ( .A(n16027), .B(n16026), .Z(n16029) );
  NANDN U16534 ( .A(n17475), .B(\stack[6][37] ), .Z(n16028) );
  NAND U16535 ( .A(n16029), .B(n16028), .Z(n2336) );
  NANDN U16536 ( .A(n2967), .B(\stack[4][37] ), .Z(n16031) );
  NANDN U16537 ( .A(n17472), .B(\stack[6][37] ), .Z(n16030) );
  AND U16538 ( .A(n16031), .B(n16030), .Z(n16033) );
  NANDN U16539 ( .A(n17475), .B(\stack[5][37] ), .Z(n16032) );
  NAND U16540 ( .A(n16033), .B(n16032), .Z(n2337) );
  NANDN U16541 ( .A(n2967), .B(\stack[3][37] ), .Z(n16035) );
  NANDN U16542 ( .A(n17472), .B(\stack[5][37] ), .Z(n16034) );
  AND U16543 ( .A(n16035), .B(n16034), .Z(n16037) );
  NANDN U16544 ( .A(n17475), .B(\stack[4][37] ), .Z(n16036) );
  NAND U16545 ( .A(n16037), .B(n16036), .Z(n2338) );
  NANDN U16546 ( .A(n2967), .B(\stack[2][37] ), .Z(n16039) );
  NANDN U16547 ( .A(n17472), .B(\stack[4][37] ), .Z(n16038) );
  AND U16548 ( .A(n16039), .B(n16038), .Z(n16041) );
  NANDN U16549 ( .A(n17475), .B(\stack[3][37] ), .Z(n16040) );
  NAND U16550 ( .A(n16041), .B(n16040), .Z(n2339) );
  NANDN U16551 ( .A(n2967), .B(\stack[1][37] ), .Z(n16043) );
  NANDN U16552 ( .A(n17472), .B(\stack[3][37] ), .Z(n16042) );
  AND U16553 ( .A(n16043), .B(n16042), .Z(n16045) );
  NANDN U16554 ( .A(n17475), .B(\stack[2][37] ), .Z(n16044) );
  NAND U16555 ( .A(n16045), .B(n16044), .Z(n2340) );
  NANDN U16556 ( .A(n2967), .B(o[37]), .Z(n16047) );
  NANDN U16557 ( .A(n17472), .B(\stack[2][37] ), .Z(n16046) );
  AND U16558 ( .A(n16047), .B(n16046), .Z(n16049) );
  NANDN U16559 ( .A(n17475), .B(\stack[1][37] ), .Z(n16048) );
  NAND U16560 ( .A(n16049), .B(n16048), .Z(n2341) );
  NAND U16561 ( .A(\stack[1][37] ), .B(n17479), .Z(n16050) );
  NANDN U16562 ( .A(n17467), .B(n16050), .Z(n16051) );
  AND U16563 ( .A(n16051), .B(o[37]), .Z(n16060) );
  XNOR U16564 ( .A(n16053), .B(n16052), .Z(n16054) );
  NAND U16565 ( .A(n16054), .B(n17458), .Z(n16058) );
  NANDN U16566 ( .A(n2967), .B(x[37]), .Z(n16056) );
  NANDN U16567 ( .A(n17483), .B(\stack[1][37] ), .Z(n16055) );
  AND U16568 ( .A(n16056), .B(n16055), .Z(n16057) );
  NAND U16569 ( .A(n16058), .B(n16057), .Z(n16059) );
  NOR U16570 ( .A(n16060), .B(n16059), .Z(n16061) );
  NANDN U16571 ( .A(n2967), .B(\stack[6][36] ), .Z(n16063) );
  NANDN U16572 ( .A(n17471), .B(\stack[7][36] ), .Z(n16062) );
  NAND U16573 ( .A(n16063), .B(n16062), .Z(n2343) );
  NANDN U16574 ( .A(n2967), .B(\stack[5][36] ), .Z(n16065) );
  NANDN U16575 ( .A(n17472), .B(\stack[7][36] ), .Z(n16064) );
  AND U16576 ( .A(n16065), .B(n16064), .Z(n16067) );
  NANDN U16577 ( .A(n17475), .B(\stack[6][36] ), .Z(n16066) );
  NAND U16578 ( .A(n16067), .B(n16066), .Z(n2344) );
  NANDN U16579 ( .A(n2967), .B(\stack[4][36] ), .Z(n16069) );
  NANDN U16580 ( .A(n17472), .B(\stack[6][36] ), .Z(n16068) );
  AND U16581 ( .A(n16069), .B(n16068), .Z(n16071) );
  NANDN U16582 ( .A(n17475), .B(\stack[5][36] ), .Z(n16070) );
  NAND U16583 ( .A(n16071), .B(n16070), .Z(n2345) );
  NANDN U16584 ( .A(n2967), .B(\stack[3][36] ), .Z(n16073) );
  NANDN U16585 ( .A(n17472), .B(\stack[5][36] ), .Z(n16072) );
  AND U16586 ( .A(n16073), .B(n16072), .Z(n16075) );
  NANDN U16587 ( .A(n17475), .B(\stack[4][36] ), .Z(n16074) );
  NAND U16588 ( .A(n16075), .B(n16074), .Z(n2346) );
  NANDN U16589 ( .A(n2967), .B(\stack[2][36] ), .Z(n16077) );
  NANDN U16590 ( .A(n17472), .B(\stack[4][36] ), .Z(n16076) );
  AND U16591 ( .A(n16077), .B(n16076), .Z(n16079) );
  NANDN U16592 ( .A(n17475), .B(\stack[3][36] ), .Z(n16078) );
  NAND U16593 ( .A(n16079), .B(n16078), .Z(n2347) );
  NANDN U16594 ( .A(n2993), .B(n17471), .Z(n16081) );
  NANDN U16595 ( .A(n17472), .B(\stack[3][36] ), .Z(n16080) );
  AND U16596 ( .A(n16081), .B(n16080), .Z(n16083) );
  NANDN U16597 ( .A(n17475), .B(\stack[2][36] ), .Z(n16082) );
  NAND U16598 ( .A(n16083), .B(n16082), .Z(n2348) );
  NANDN U16599 ( .A(n2967), .B(o[36]), .Z(n16085) );
  NANDN U16600 ( .A(n17472), .B(\stack[2][36] ), .Z(n16084) );
  AND U16601 ( .A(n16085), .B(n16084), .Z(n16087) );
  OR U16602 ( .A(n17475), .B(n2993), .Z(n16086) );
  NAND U16603 ( .A(n16087), .B(n16086), .Z(n2349) );
  NAND U16604 ( .A(o[36]), .B(n17479), .Z(n16088) );
  NANDN U16605 ( .A(n17461), .B(n16088), .Z(n16089) );
  ANDN U16606 ( .B(n16089), .A(n2993), .Z(n16097) );
  XNOR U16607 ( .A(n16091), .B(n16090), .Z(n16092) );
  NAND U16608 ( .A(n16092), .B(n17458), .Z(n16095) );
  NANDN U16609 ( .A(n2967), .B(x[36]), .Z(n16093) );
  NAND U16610 ( .A(n16095), .B(n16094), .Z(n16096) );
  NOR U16611 ( .A(n16097), .B(n16096), .Z(n16099) );
  NANDN U16612 ( .A(n17481), .B(o[36]), .Z(n16098) );
  NAND U16613 ( .A(n16099), .B(n16098), .Z(n2350) );
  NANDN U16614 ( .A(n2967), .B(\stack[6][35] ), .Z(n16101) );
  NANDN U16615 ( .A(n17471), .B(\stack[7][35] ), .Z(n16100) );
  NAND U16616 ( .A(n16101), .B(n16100), .Z(n2351) );
  NANDN U16617 ( .A(n2967), .B(\stack[5][35] ), .Z(n16103) );
  NANDN U16618 ( .A(n17472), .B(\stack[7][35] ), .Z(n16102) );
  AND U16619 ( .A(n16103), .B(n16102), .Z(n16105) );
  NANDN U16620 ( .A(n17475), .B(\stack[6][35] ), .Z(n16104) );
  NAND U16621 ( .A(n16105), .B(n16104), .Z(n2352) );
  NANDN U16622 ( .A(n2967), .B(\stack[4][35] ), .Z(n16107) );
  NANDN U16623 ( .A(n17472), .B(\stack[6][35] ), .Z(n16106) );
  AND U16624 ( .A(n16107), .B(n16106), .Z(n16109) );
  NANDN U16625 ( .A(n17475), .B(\stack[5][35] ), .Z(n16108) );
  NAND U16626 ( .A(n16109), .B(n16108), .Z(n2353) );
  NANDN U16627 ( .A(n2967), .B(\stack[3][35] ), .Z(n16111) );
  NANDN U16628 ( .A(n17472), .B(\stack[5][35] ), .Z(n16110) );
  AND U16629 ( .A(n16111), .B(n16110), .Z(n16113) );
  NANDN U16630 ( .A(n17475), .B(\stack[4][35] ), .Z(n16112) );
  NAND U16631 ( .A(n16113), .B(n16112), .Z(n2354) );
  NANDN U16632 ( .A(n2967), .B(\stack[2][35] ), .Z(n16115) );
  NANDN U16633 ( .A(n17472), .B(\stack[4][35] ), .Z(n16114) );
  AND U16634 ( .A(n16115), .B(n16114), .Z(n16117) );
  NANDN U16635 ( .A(n17475), .B(\stack[3][35] ), .Z(n16116) );
  NAND U16636 ( .A(n16117), .B(n16116), .Z(n2355) );
  NANDN U16637 ( .A(n2992), .B(n17471), .Z(n16119) );
  NANDN U16638 ( .A(n17472), .B(\stack[3][35] ), .Z(n16118) );
  AND U16639 ( .A(n16119), .B(n16118), .Z(n16121) );
  NANDN U16640 ( .A(n17475), .B(\stack[2][35] ), .Z(n16120) );
  NAND U16641 ( .A(n16121), .B(n16120), .Z(n2356) );
  NANDN U16642 ( .A(n2967), .B(o[35]), .Z(n16123) );
  NANDN U16643 ( .A(n17472), .B(\stack[2][35] ), .Z(n16122) );
  AND U16644 ( .A(n16123), .B(n16122), .Z(n16125) );
  OR U16645 ( .A(n17475), .B(n2992), .Z(n16124) );
  NAND U16646 ( .A(n16125), .B(n16124), .Z(n2357) );
  NANDN U16647 ( .A(n2992), .B(n17479), .Z(n16126) );
  NANDN U16648 ( .A(n17467), .B(n16126), .Z(n16127) );
  AND U16649 ( .A(n16127), .B(o[35]), .Z(n16136) );
  XNOR U16650 ( .A(n16129), .B(n16128), .Z(n16130) );
  NAND U16651 ( .A(n16130), .B(n17458), .Z(n16134) );
  NANDN U16652 ( .A(n2967), .B(x[35]), .Z(n16132) );
  NANDN U16653 ( .A(n17483), .B(\stack[1][35] ), .Z(n16131) );
  AND U16654 ( .A(n16132), .B(n16131), .Z(n16133) );
  NAND U16655 ( .A(n16134), .B(n16133), .Z(n16135) );
  NOR U16656 ( .A(n16136), .B(n16135), .Z(n16137) );
  NANDN U16657 ( .A(n2967), .B(\stack[6][34] ), .Z(n16139) );
  NANDN U16658 ( .A(n17471), .B(\stack[7][34] ), .Z(n16138) );
  NAND U16659 ( .A(n16139), .B(n16138), .Z(n2359) );
  NANDN U16660 ( .A(n2967), .B(\stack[5][34] ), .Z(n16141) );
  NANDN U16661 ( .A(n17472), .B(\stack[7][34] ), .Z(n16140) );
  AND U16662 ( .A(n16141), .B(n16140), .Z(n16143) );
  NANDN U16663 ( .A(n17475), .B(\stack[6][34] ), .Z(n16142) );
  NAND U16664 ( .A(n16143), .B(n16142), .Z(n2360) );
  NANDN U16665 ( .A(n2967), .B(\stack[4][34] ), .Z(n16145) );
  NANDN U16666 ( .A(n17472), .B(\stack[6][34] ), .Z(n16144) );
  AND U16667 ( .A(n16145), .B(n16144), .Z(n16147) );
  NANDN U16668 ( .A(n17475), .B(\stack[5][34] ), .Z(n16146) );
  NAND U16669 ( .A(n16147), .B(n16146), .Z(n2361) );
  NANDN U16670 ( .A(n2967), .B(\stack[3][34] ), .Z(n16149) );
  NANDN U16671 ( .A(n17472), .B(\stack[5][34] ), .Z(n16148) );
  AND U16672 ( .A(n16149), .B(n16148), .Z(n16151) );
  NANDN U16673 ( .A(n17475), .B(\stack[4][34] ), .Z(n16150) );
  NAND U16674 ( .A(n16151), .B(n16150), .Z(n2362) );
  NANDN U16675 ( .A(n2967), .B(\stack[2][34] ), .Z(n16153) );
  NANDN U16676 ( .A(n17472), .B(\stack[4][34] ), .Z(n16152) );
  AND U16677 ( .A(n16153), .B(n16152), .Z(n16155) );
  NANDN U16678 ( .A(n17475), .B(\stack[3][34] ), .Z(n16154) );
  NAND U16679 ( .A(n16155), .B(n16154), .Z(n2363) );
  NANDN U16680 ( .A(n2991), .B(n17471), .Z(n16157) );
  NANDN U16681 ( .A(n17472), .B(\stack[3][34] ), .Z(n16156) );
  AND U16682 ( .A(n16157), .B(n16156), .Z(n16159) );
  NANDN U16683 ( .A(n17475), .B(\stack[2][34] ), .Z(n16158) );
  NAND U16684 ( .A(n16159), .B(n16158), .Z(n2364) );
  NANDN U16685 ( .A(n2967), .B(o[34]), .Z(n16161) );
  NANDN U16686 ( .A(n17472), .B(\stack[2][34] ), .Z(n16160) );
  AND U16687 ( .A(n16161), .B(n16160), .Z(n16163) );
  OR U16688 ( .A(n17475), .B(n2991), .Z(n16162) );
  NAND U16689 ( .A(n16163), .B(n16162), .Z(n2365) );
  NAND U16690 ( .A(o[34]), .B(n17479), .Z(n16164) );
  NANDN U16691 ( .A(n17461), .B(n16164), .Z(n16165) );
  ANDN U16692 ( .B(n16165), .A(n2991), .Z(n16173) );
  XNOR U16693 ( .A(n16167), .B(n16166), .Z(n16168) );
  NAND U16694 ( .A(n16168), .B(n17458), .Z(n16171) );
  NANDN U16695 ( .A(n2967), .B(x[34]), .Z(n16169) );
  NAND U16696 ( .A(n16171), .B(n16170), .Z(n16172) );
  NOR U16697 ( .A(n16173), .B(n16172), .Z(n16175) );
  NANDN U16698 ( .A(n17481), .B(o[34]), .Z(n16174) );
  NAND U16699 ( .A(n16175), .B(n16174), .Z(n2366) );
  NANDN U16700 ( .A(n2967), .B(\stack[6][33] ), .Z(n16177) );
  NANDN U16701 ( .A(n17471), .B(\stack[7][33] ), .Z(n16176) );
  NAND U16702 ( .A(n16177), .B(n16176), .Z(n2367) );
  NANDN U16703 ( .A(n2967), .B(\stack[5][33] ), .Z(n16179) );
  NANDN U16704 ( .A(n17472), .B(\stack[7][33] ), .Z(n16178) );
  AND U16705 ( .A(n16179), .B(n16178), .Z(n16181) );
  NANDN U16706 ( .A(n17475), .B(\stack[6][33] ), .Z(n16180) );
  NAND U16707 ( .A(n16181), .B(n16180), .Z(n2368) );
  NANDN U16708 ( .A(n2967), .B(\stack[4][33] ), .Z(n16183) );
  NANDN U16709 ( .A(n17472), .B(\stack[6][33] ), .Z(n16182) );
  AND U16710 ( .A(n16183), .B(n16182), .Z(n16185) );
  NANDN U16711 ( .A(n17475), .B(\stack[5][33] ), .Z(n16184) );
  NAND U16712 ( .A(n16185), .B(n16184), .Z(n2369) );
  NANDN U16713 ( .A(n2967), .B(\stack[3][33] ), .Z(n16187) );
  NANDN U16714 ( .A(n17472), .B(\stack[5][33] ), .Z(n16186) );
  AND U16715 ( .A(n16187), .B(n16186), .Z(n16189) );
  NANDN U16716 ( .A(n17475), .B(\stack[4][33] ), .Z(n16188) );
  NAND U16717 ( .A(n16189), .B(n16188), .Z(n2370) );
  NANDN U16718 ( .A(n2967), .B(\stack[2][33] ), .Z(n16191) );
  NANDN U16719 ( .A(n17472), .B(\stack[4][33] ), .Z(n16190) );
  AND U16720 ( .A(n16191), .B(n16190), .Z(n16193) );
  NANDN U16721 ( .A(n17475), .B(\stack[3][33] ), .Z(n16192) );
  NAND U16722 ( .A(n16193), .B(n16192), .Z(n2371) );
  NANDN U16723 ( .A(n2990), .B(n17471), .Z(n16195) );
  NANDN U16724 ( .A(n17472), .B(\stack[3][33] ), .Z(n16194) );
  AND U16725 ( .A(n16195), .B(n16194), .Z(n16197) );
  NANDN U16726 ( .A(n17475), .B(\stack[2][33] ), .Z(n16196) );
  NAND U16727 ( .A(n16197), .B(n16196), .Z(n2372) );
  NANDN U16728 ( .A(n2967), .B(o[33]), .Z(n16199) );
  NANDN U16729 ( .A(n17472), .B(\stack[2][33] ), .Z(n16198) );
  AND U16730 ( .A(n16199), .B(n16198), .Z(n16201) );
  OR U16731 ( .A(n17475), .B(n2990), .Z(n16200) );
  NAND U16732 ( .A(n16201), .B(n16200), .Z(n2373) );
  NANDN U16733 ( .A(n2990), .B(n17479), .Z(n16202) );
  NANDN U16734 ( .A(n17467), .B(n16202), .Z(n16203) );
  AND U16735 ( .A(n16203), .B(o[33]), .Z(n16212) );
  XNOR U16736 ( .A(n16205), .B(n16204), .Z(n16206) );
  NAND U16737 ( .A(n16206), .B(n17458), .Z(n16210) );
  NANDN U16738 ( .A(n2967), .B(x[33]), .Z(n16208) );
  NANDN U16739 ( .A(n17483), .B(\stack[1][33] ), .Z(n16207) );
  AND U16740 ( .A(n16208), .B(n16207), .Z(n16209) );
  NAND U16741 ( .A(n16210), .B(n16209), .Z(n16211) );
  NOR U16742 ( .A(n16212), .B(n16211), .Z(n16213) );
  NANDN U16743 ( .A(n2967), .B(\stack[6][32] ), .Z(n16215) );
  NANDN U16744 ( .A(n17471), .B(\stack[7][32] ), .Z(n16214) );
  NAND U16745 ( .A(n16215), .B(n16214), .Z(n2375) );
  NANDN U16746 ( .A(n2967), .B(\stack[5][32] ), .Z(n16217) );
  NANDN U16747 ( .A(n17472), .B(\stack[7][32] ), .Z(n16216) );
  AND U16748 ( .A(n16217), .B(n16216), .Z(n16219) );
  NANDN U16749 ( .A(n17475), .B(\stack[6][32] ), .Z(n16218) );
  NAND U16750 ( .A(n16219), .B(n16218), .Z(n2376) );
  NANDN U16751 ( .A(n2967), .B(\stack[4][32] ), .Z(n16221) );
  NANDN U16752 ( .A(n17472), .B(\stack[6][32] ), .Z(n16220) );
  AND U16753 ( .A(n16221), .B(n16220), .Z(n16223) );
  NANDN U16754 ( .A(n17475), .B(\stack[5][32] ), .Z(n16222) );
  NAND U16755 ( .A(n16223), .B(n16222), .Z(n2377) );
  NANDN U16756 ( .A(n2967), .B(\stack[3][32] ), .Z(n16225) );
  NANDN U16757 ( .A(n17472), .B(\stack[5][32] ), .Z(n16224) );
  AND U16758 ( .A(n16225), .B(n16224), .Z(n16227) );
  NANDN U16759 ( .A(n17475), .B(\stack[4][32] ), .Z(n16226) );
  NAND U16760 ( .A(n16227), .B(n16226), .Z(n2378) );
  NANDN U16761 ( .A(n2967), .B(\stack[2][32] ), .Z(n16229) );
  NANDN U16762 ( .A(n17472), .B(\stack[4][32] ), .Z(n16228) );
  AND U16763 ( .A(n16229), .B(n16228), .Z(n16231) );
  NANDN U16764 ( .A(n17475), .B(\stack[3][32] ), .Z(n16230) );
  NAND U16765 ( .A(n16231), .B(n16230), .Z(n2379) );
  NANDN U16766 ( .A(n2989), .B(n17471), .Z(n16233) );
  NANDN U16767 ( .A(n17472), .B(\stack[3][32] ), .Z(n16232) );
  AND U16768 ( .A(n16233), .B(n16232), .Z(n16235) );
  NANDN U16769 ( .A(n17475), .B(\stack[2][32] ), .Z(n16234) );
  NAND U16770 ( .A(n16235), .B(n16234), .Z(n2380) );
  NANDN U16771 ( .A(n2967), .B(o[32]), .Z(n16237) );
  NANDN U16772 ( .A(n17472), .B(\stack[2][32] ), .Z(n16236) );
  AND U16773 ( .A(n16237), .B(n16236), .Z(n16239) );
  OR U16774 ( .A(n17475), .B(n2989), .Z(n16238) );
  NAND U16775 ( .A(n16239), .B(n16238), .Z(n2381) );
  NAND U16776 ( .A(o[32]), .B(n17479), .Z(n16240) );
  NANDN U16777 ( .A(n17461), .B(n16240), .Z(n16241) );
  ANDN U16778 ( .B(n16241), .A(n2989), .Z(n16249) );
  XNOR U16779 ( .A(n16243), .B(n16242), .Z(n16244) );
  NAND U16780 ( .A(n16244), .B(n17458), .Z(n16247) );
  NANDN U16781 ( .A(n2967), .B(x[32]), .Z(n16245) );
  NAND U16782 ( .A(n16247), .B(n16246), .Z(n16248) );
  NOR U16783 ( .A(n16249), .B(n16248), .Z(n16251) );
  NANDN U16784 ( .A(n17481), .B(o[32]), .Z(n16250) );
  NAND U16785 ( .A(n16251), .B(n16250), .Z(n2382) );
  NANDN U16786 ( .A(n2967), .B(\stack[6][31] ), .Z(n16253) );
  NANDN U16787 ( .A(n17471), .B(\stack[7][31] ), .Z(n16252) );
  NAND U16788 ( .A(n16253), .B(n16252), .Z(n2383) );
  NANDN U16789 ( .A(n2967), .B(\stack[5][31] ), .Z(n16255) );
  NANDN U16790 ( .A(n17472), .B(\stack[7][31] ), .Z(n16254) );
  AND U16791 ( .A(n16255), .B(n16254), .Z(n16257) );
  NANDN U16792 ( .A(n17475), .B(\stack[6][31] ), .Z(n16256) );
  NAND U16793 ( .A(n16257), .B(n16256), .Z(n2384) );
  NANDN U16794 ( .A(n2967), .B(\stack[4][31] ), .Z(n16259) );
  NANDN U16795 ( .A(n17472), .B(\stack[6][31] ), .Z(n16258) );
  AND U16796 ( .A(n16259), .B(n16258), .Z(n16261) );
  NANDN U16797 ( .A(n17475), .B(\stack[5][31] ), .Z(n16260) );
  NAND U16798 ( .A(n16261), .B(n16260), .Z(n2385) );
  NANDN U16799 ( .A(n2967), .B(\stack[3][31] ), .Z(n16263) );
  NANDN U16800 ( .A(n17472), .B(\stack[5][31] ), .Z(n16262) );
  AND U16801 ( .A(n16263), .B(n16262), .Z(n16265) );
  NANDN U16802 ( .A(n17475), .B(\stack[4][31] ), .Z(n16264) );
  NAND U16803 ( .A(n16265), .B(n16264), .Z(n2386) );
  NANDN U16804 ( .A(n2967), .B(\stack[2][31] ), .Z(n16267) );
  NANDN U16805 ( .A(n17472), .B(\stack[4][31] ), .Z(n16266) );
  AND U16806 ( .A(n16267), .B(n16266), .Z(n16269) );
  NANDN U16807 ( .A(n17475), .B(\stack[3][31] ), .Z(n16268) );
  NAND U16808 ( .A(n16269), .B(n16268), .Z(n2387) );
  NANDN U16809 ( .A(n2988), .B(n17471), .Z(n16271) );
  NANDN U16810 ( .A(n17472), .B(\stack[3][31] ), .Z(n16270) );
  AND U16811 ( .A(n16271), .B(n16270), .Z(n16273) );
  NANDN U16812 ( .A(n17475), .B(\stack[2][31] ), .Z(n16272) );
  NAND U16813 ( .A(n16273), .B(n16272), .Z(n2388) );
  NANDN U16814 ( .A(n2967), .B(o[31]), .Z(n16275) );
  NANDN U16815 ( .A(n17472), .B(\stack[2][31] ), .Z(n16274) );
  AND U16816 ( .A(n16275), .B(n16274), .Z(n16277) );
  OR U16817 ( .A(n17475), .B(n2988), .Z(n16276) );
  NAND U16818 ( .A(n16277), .B(n16276), .Z(n2389) );
  NANDN U16819 ( .A(n2967), .B(x[31]), .Z(n16279) );
  NANDN U16820 ( .A(n17483), .B(\stack[1][31] ), .Z(n16278) );
  NAND U16821 ( .A(n16279), .B(n16278), .Z(n16288) );
  XNOR U16822 ( .A(n16281), .B(n16280), .Z(n16282) );
  NAND U16823 ( .A(n16282), .B(n17458), .Z(n16286) );
  NAND U16824 ( .A(n16283), .B(n17479), .Z(n16284) );
  NAND U16825 ( .A(n16286), .B(n16285), .Z(n16287) );
  NOR U16826 ( .A(n16288), .B(n16287), .Z(n16290) );
  NANDN U16827 ( .A(n17481), .B(o[31]), .Z(n16289) );
  NAND U16828 ( .A(n16290), .B(n16289), .Z(n2390) );
  NANDN U16829 ( .A(n2967), .B(\stack[6][30] ), .Z(n16292) );
  NANDN U16830 ( .A(n17471), .B(\stack[7][30] ), .Z(n16291) );
  NAND U16831 ( .A(n16292), .B(n16291), .Z(n2391) );
  NANDN U16832 ( .A(n2967), .B(\stack[5][30] ), .Z(n16294) );
  NANDN U16833 ( .A(n17472), .B(\stack[7][30] ), .Z(n16293) );
  AND U16834 ( .A(n16294), .B(n16293), .Z(n16296) );
  NANDN U16835 ( .A(n17475), .B(\stack[6][30] ), .Z(n16295) );
  NAND U16836 ( .A(n16296), .B(n16295), .Z(n2392) );
  NANDN U16837 ( .A(n2967), .B(\stack[4][30] ), .Z(n16298) );
  NANDN U16838 ( .A(n17472), .B(\stack[6][30] ), .Z(n16297) );
  AND U16839 ( .A(n16298), .B(n16297), .Z(n16300) );
  NANDN U16840 ( .A(n17475), .B(\stack[5][30] ), .Z(n16299) );
  NAND U16841 ( .A(n16300), .B(n16299), .Z(n2393) );
  NANDN U16842 ( .A(n2967), .B(\stack[3][30] ), .Z(n16302) );
  NANDN U16843 ( .A(n17472), .B(\stack[5][30] ), .Z(n16301) );
  AND U16844 ( .A(n16302), .B(n16301), .Z(n16304) );
  NANDN U16845 ( .A(n17475), .B(\stack[4][30] ), .Z(n16303) );
  NAND U16846 ( .A(n16304), .B(n16303), .Z(n2394) );
  NANDN U16847 ( .A(n2967), .B(\stack[2][30] ), .Z(n16306) );
  NANDN U16848 ( .A(n17472), .B(\stack[4][30] ), .Z(n16305) );
  AND U16849 ( .A(n16306), .B(n16305), .Z(n16308) );
  NANDN U16850 ( .A(n17475), .B(\stack[3][30] ), .Z(n16307) );
  NAND U16851 ( .A(n16308), .B(n16307), .Z(n2395) );
  NANDN U16852 ( .A(n2987), .B(n17471), .Z(n16310) );
  NANDN U16853 ( .A(n17472), .B(\stack[3][30] ), .Z(n16309) );
  AND U16854 ( .A(n16310), .B(n16309), .Z(n16312) );
  NANDN U16855 ( .A(n17475), .B(\stack[2][30] ), .Z(n16311) );
  NAND U16856 ( .A(n16312), .B(n16311), .Z(n2396) );
  NANDN U16857 ( .A(n2967), .B(o[30]), .Z(n16314) );
  NANDN U16858 ( .A(n17472), .B(\stack[2][30] ), .Z(n16313) );
  AND U16859 ( .A(n16314), .B(n16313), .Z(n16316) );
  OR U16860 ( .A(n17475), .B(n2987), .Z(n16315) );
  NAND U16861 ( .A(n16316), .B(n16315), .Z(n2397) );
  NANDN U16862 ( .A(n2967), .B(x[30]), .Z(n16319) );
  NANDN U16863 ( .A(n16317), .B(n17479), .Z(n16318) );
  NAND U16864 ( .A(n16319), .B(n16318), .Z(n16327) );
  XNOR U16865 ( .A(n16321), .B(n16320), .Z(n16322) );
  NAND U16866 ( .A(n16322), .B(n17458), .Z(n16325) );
  NANDN U16867 ( .A(n2987), .B(n17461), .Z(n16323) );
  NAND U16868 ( .A(n16325), .B(n16324), .Z(n16326) );
  NOR U16869 ( .A(n16327), .B(n16326), .Z(n16329) );
  NANDN U16870 ( .A(n17481), .B(o[30]), .Z(n16328) );
  NAND U16871 ( .A(n16329), .B(n16328), .Z(n2398) );
  NANDN U16872 ( .A(n2967), .B(\stack[6][29] ), .Z(n16331) );
  NANDN U16873 ( .A(n17471), .B(\stack[7][29] ), .Z(n16330) );
  NAND U16874 ( .A(n16331), .B(n16330), .Z(n2399) );
  NANDN U16875 ( .A(n2967), .B(\stack[5][29] ), .Z(n16333) );
  NANDN U16876 ( .A(n17472), .B(\stack[7][29] ), .Z(n16332) );
  AND U16877 ( .A(n16333), .B(n16332), .Z(n16335) );
  NANDN U16878 ( .A(n17475), .B(\stack[6][29] ), .Z(n16334) );
  NAND U16879 ( .A(n16335), .B(n16334), .Z(n2400) );
  NANDN U16880 ( .A(n2967), .B(\stack[4][29] ), .Z(n16337) );
  NANDN U16881 ( .A(n17472), .B(\stack[6][29] ), .Z(n16336) );
  AND U16882 ( .A(n16337), .B(n16336), .Z(n16339) );
  NANDN U16883 ( .A(n17475), .B(\stack[5][29] ), .Z(n16338) );
  NAND U16884 ( .A(n16339), .B(n16338), .Z(n2401) );
  NANDN U16885 ( .A(n2967), .B(\stack[3][29] ), .Z(n16341) );
  NANDN U16886 ( .A(n17472), .B(\stack[5][29] ), .Z(n16340) );
  AND U16887 ( .A(n16341), .B(n16340), .Z(n16343) );
  NANDN U16888 ( .A(n17475), .B(\stack[4][29] ), .Z(n16342) );
  NAND U16889 ( .A(n16343), .B(n16342), .Z(n2402) );
  NANDN U16890 ( .A(n2967), .B(\stack[2][29] ), .Z(n16345) );
  NANDN U16891 ( .A(n17472), .B(\stack[4][29] ), .Z(n16344) );
  AND U16892 ( .A(n16345), .B(n16344), .Z(n16347) );
  NANDN U16893 ( .A(n17475), .B(\stack[3][29] ), .Z(n16346) );
  NAND U16894 ( .A(n16347), .B(n16346), .Z(n2403) );
  NANDN U16895 ( .A(n2986), .B(n17471), .Z(n16349) );
  NANDN U16896 ( .A(n17472), .B(\stack[3][29] ), .Z(n16348) );
  AND U16897 ( .A(n16349), .B(n16348), .Z(n16351) );
  NANDN U16898 ( .A(n17475), .B(\stack[2][29] ), .Z(n16350) );
  NAND U16899 ( .A(n16351), .B(n16350), .Z(n2404) );
  NANDN U16900 ( .A(n2967), .B(o[29]), .Z(n16353) );
  NANDN U16901 ( .A(n17472), .B(\stack[2][29] ), .Z(n16352) );
  AND U16902 ( .A(n16353), .B(n16352), .Z(n16355) );
  OR U16903 ( .A(n17475), .B(n2986), .Z(n16354) );
  NAND U16904 ( .A(n16355), .B(n16354), .Z(n2405) );
  NANDN U16905 ( .A(n2986), .B(n17479), .Z(n16356) );
  NANDN U16906 ( .A(n17467), .B(n16356), .Z(n16357) );
  AND U16907 ( .A(n16357), .B(o[29]), .Z(n16366) );
  NANDN U16908 ( .A(n2967), .B(x[29]), .Z(n16359) );
  NANDN U16909 ( .A(n17483), .B(\stack[1][29] ), .Z(n16358) );
  NAND U16910 ( .A(n16359), .B(n16358), .Z(n16364) );
  XNOR U16911 ( .A(n16361), .B(n16360), .Z(n16362) );
  NAND U16912 ( .A(n16362), .B(n17458), .Z(n16363) );
  NANDN U16913 ( .A(n16364), .B(n16363), .Z(n16365) );
  NOR U16914 ( .A(n16366), .B(n16365), .Z(n16367) );
  NANDN U16915 ( .A(n2967), .B(\stack[6][28] ), .Z(n16369) );
  NANDN U16916 ( .A(n17471), .B(\stack[7][28] ), .Z(n16368) );
  NAND U16917 ( .A(n16369), .B(n16368), .Z(n2407) );
  NANDN U16918 ( .A(n2967), .B(\stack[5][28] ), .Z(n16371) );
  NANDN U16919 ( .A(n17472), .B(\stack[7][28] ), .Z(n16370) );
  AND U16920 ( .A(n16371), .B(n16370), .Z(n16373) );
  NANDN U16921 ( .A(n17475), .B(\stack[6][28] ), .Z(n16372) );
  NAND U16922 ( .A(n16373), .B(n16372), .Z(n2408) );
  NANDN U16923 ( .A(n2967), .B(\stack[4][28] ), .Z(n16375) );
  NANDN U16924 ( .A(n17472), .B(\stack[6][28] ), .Z(n16374) );
  AND U16925 ( .A(n16375), .B(n16374), .Z(n16377) );
  NANDN U16926 ( .A(n17475), .B(\stack[5][28] ), .Z(n16376) );
  NAND U16927 ( .A(n16377), .B(n16376), .Z(n2409) );
  NANDN U16928 ( .A(n2967), .B(\stack[3][28] ), .Z(n16379) );
  NANDN U16929 ( .A(n17472), .B(\stack[5][28] ), .Z(n16378) );
  AND U16930 ( .A(n16379), .B(n16378), .Z(n16381) );
  NANDN U16931 ( .A(n17475), .B(\stack[4][28] ), .Z(n16380) );
  NAND U16932 ( .A(n16381), .B(n16380), .Z(n2410) );
  NANDN U16933 ( .A(n2967), .B(\stack[2][28] ), .Z(n16383) );
  NANDN U16934 ( .A(n17472), .B(\stack[4][28] ), .Z(n16382) );
  AND U16935 ( .A(n16383), .B(n16382), .Z(n16385) );
  NANDN U16936 ( .A(n17475), .B(\stack[3][28] ), .Z(n16384) );
  NAND U16937 ( .A(n16385), .B(n16384), .Z(n2411) );
  NANDN U16938 ( .A(n2985), .B(n17471), .Z(n16387) );
  NANDN U16939 ( .A(n17472), .B(\stack[3][28] ), .Z(n16386) );
  AND U16940 ( .A(n16387), .B(n16386), .Z(n16389) );
  NANDN U16941 ( .A(n17475), .B(\stack[2][28] ), .Z(n16388) );
  NAND U16942 ( .A(n16389), .B(n16388), .Z(n2412) );
  NANDN U16943 ( .A(n3021), .B(n17471), .Z(n16391) );
  NANDN U16944 ( .A(n17472), .B(\stack[2][28] ), .Z(n16390) );
  AND U16945 ( .A(n16391), .B(n16390), .Z(n16393) );
  OR U16946 ( .A(n17475), .B(n2985), .Z(n16392) );
  NAND U16947 ( .A(n16393), .B(n16392), .Z(n2413) );
  NANDN U16948 ( .A(n2967), .B(x[28]), .Z(n16395) );
  NANDN U16949 ( .A(n17483), .B(\stack[1][28] ), .Z(n16394) );
  NAND U16950 ( .A(n16395), .B(n16394), .Z(n16404) );
  XNOR U16951 ( .A(n16397), .B(n16396), .Z(n16398) );
  NAND U16952 ( .A(n16398), .B(n17458), .Z(n16402) );
  NANDN U16953 ( .A(n16399), .B(n17479), .Z(n16400) );
  NAND U16954 ( .A(n16402), .B(n16401), .Z(n16403) );
  NOR U16955 ( .A(n16404), .B(n16403), .Z(n16406) );
  NANDN U16956 ( .A(n3021), .B(n17467), .Z(n16405) );
  NAND U16957 ( .A(n16406), .B(n16405), .Z(n2414) );
  NANDN U16958 ( .A(n2967), .B(\stack[6][27] ), .Z(n16408) );
  NANDN U16959 ( .A(n17471), .B(\stack[7][27] ), .Z(n16407) );
  NAND U16960 ( .A(n16408), .B(n16407), .Z(n2415) );
  NANDN U16961 ( .A(n2967), .B(\stack[5][27] ), .Z(n16410) );
  NANDN U16962 ( .A(n17472), .B(\stack[7][27] ), .Z(n16409) );
  AND U16963 ( .A(n16410), .B(n16409), .Z(n16412) );
  NANDN U16964 ( .A(n17475), .B(\stack[6][27] ), .Z(n16411) );
  NAND U16965 ( .A(n16412), .B(n16411), .Z(n2416) );
  NANDN U16966 ( .A(n2967), .B(\stack[4][27] ), .Z(n16414) );
  NANDN U16967 ( .A(n17472), .B(\stack[6][27] ), .Z(n16413) );
  AND U16968 ( .A(n16414), .B(n16413), .Z(n16416) );
  NANDN U16969 ( .A(n17475), .B(\stack[5][27] ), .Z(n16415) );
  NAND U16970 ( .A(n16416), .B(n16415), .Z(n2417) );
  NANDN U16971 ( .A(n2967), .B(\stack[3][27] ), .Z(n16418) );
  NANDN U16972 ( .A(n17472), .B(\stack[5][27] ), .Z(n16417) );
  AND U16973 ( .A(n16418), .B(n16417), .Z(n16420) );
  NANDN U16974 ( .A(n17475), .B(\stack[4][27] ), .Z(n16419) );
  NAND U16975 ( .A(n16420), .B(n16419), .Z(n2418) );
  NANDN U16976 ( .A(n2967), .B(\stack[2][27] ), .Z(n16422) );
  NANDN U16977 ( .A(n17472), .B(\stack[4][27] ), .Z(n16421) );
  AND U16978 ( .A(n16422), .B(n16421), .Z(n16424) );
  NANDN U16979 ( .A(n17475), .B(\stack[3][27] ), .Z(n16423) );
  NAND U16980 ( .A(n16424), .B(n16423), .Z(n2419) );
  NANDN U16981 ( .A(n2984), .B(n17471), .Z(n16426) );
  NANDN U16982 ( .A(n17472), .B(\stack[3][27] ), .Z(n16425) );
  AND U16983 ( .A(n16426), .B(n16425), .Z(n16428) );
  NANDN U16984 ( .A(n17475), .B(\stack[2][27] ), .Z(n16427) );
  NAND U16985 ( .A(n16428), .B(n16427), .Z(n2420) );
  NANDN U16986 ( .A(n2967), .B(o[27]), .Z(n16430) );
  NANDN U16987 ( .A(n17472), .B(\stack[2][27] ), .Z(n16429) );
  AND U16988 ( .A(n16430), .B(n16429), .Z(n16432) );
  OR U16989 ( .A(n17475), .B(n2984), .Z(n16431) );
  NAND U16990 ( .A(n16432), .B(n16431), .Z(n2421) );
  NANDN U16991 ( .A(n2984), .B(n17461), .Z(n16435) );
  NAND U16992 ( .A(n16433), .B(n17479), .Z(n16434) );
  NAND U16993 ( .A(n16435), .B(n16434), .Z(n16443) );
  NANDN U16994 ( .A(n2967), .B(x[27]), .Z(n16436) );
  XNOR U16995 ( .A(n16438), .B(n16437), .Z(n16439) );
  NAND U16996 ( .A(n16439), .B(n17458), .Z(n16440) );
  NANDN U16997 ( .A(n16441), .B(n16440), .Z(n16442) );
  NOR U16998 ( .A(n16443), .B(n16442), .Z(n16445) );
  NANDN U16999 ( .A(n17481), .B(o[27]), .Z(n16444) );
  NAND U17000 ( .A(n16445), .B(n16444), .Z(n2422) );
  NANDN U17001 ( .A(n2967), .B(\stack[6][26] ), .Z(n16447) );
  NANDN U17002 ( .A(n17471), .B(\stack[7][26] ), .Z(n16446) );
  NAND U17003 ( .A(n16447), .B(n16446), .Z(n2423) );
  NANDN U17004 ( .A(n2967), .B(\stack[5][26] ), .Z(n16449) );
  NANDN U17005 ( .A(n17472), .B(\stack[7][26] ), .Z(n16448) );
  AND U17006 ( .A(n16449), .B(n16448), .Z(n16451) );
  NANDN U17007 ( .A(n17475), .B(\stack[6][26] ), .Z(n16450) );
  NAND U17008 ( .A(n16451), .B(n16450), .Z(n2424) );
  NANDN U17009 ( .A(n2967), .B(\stack[4][26] ), .Z(n16453) );
  NANDN U17010 ( .A(n17472), .B(\stack[6][26] ), .Z(n16452) );
  AND U17011 ( .A(n16453), .B(n16452), .Z(n16455) );
  NANDN U17012 ( .A(n17475), .B(\stack[5][26] ), .Z(n16454) );
  NAND U17013 ( .A(n16455), .B(n16454), .Z(n2425) );
  NANDN U17014 ( .A(n2967), .B(\stack[3][26] ), .Z(n16457) );
  NANDN U17015 ( .A(n17472), .B(\stack[5][26] ), .Z(n16456) );
  AND U17016 ( .A(n16457), .B(n16456), .Z(n16459) );
  NANDN U17017 ( .A(n17475), .B(\stack[4][26] ), .Z(n16458) );
  NAND U17018 ( .A(n16459), .B(n16458), .Z(n2426) );
  NANDN U17019 ( .A(n2967), .B(\stack[2][26] ), .Z(n16461) );
  NANDN U17020 ( .A(n17472), .B(\stack[4][26] ), .Z(n16460) );
  AND U17021 ( .A(n16461), .B(n16460), .Z(n16463) );
  NANDN U17022 ( .A(n17475), .B(\stack[3][26] ), .Z(n16462) );
  NAND U17023 ( .A(n16463), .B(n16462), .Z(n2427) );
  NANDN U17024 ( .A(n2983), .B(n17471), .Z(n16465) );
  NANDN U17025 ( .A(n17472), .B(\stack[3][26] ), .Z(n16464) );
  AND U17026 ( .A(n16465), .B(n16464), .Z(n16467) );
  NANDN U17027 ( .A(n17475), .B(\stack[2][26] ), .Z(n16466) );
  NAND U17028 ( .A(n16467), .B(n16466), .Z(n2428) );
  NANDN U17029 ( .A(n3020), .B(n17471), .Z(n16469) );
  NANDN U17030 ( .A(n17472), .B(\stack[2][26] ), .Z(n16468) );
  AND U17031 ( .A(n16469), .B(n16468), .Z(n16471) );
  OR U17032 ( .A(n17475), .B(n2983), .Z(n16470) );
  NAND U17033 ( .A(n16471), .B(n16470), .Z(n2429) );
  NANDN U17034 ( .A(n2983), .B(n17461), .Z(n16474) );
  NANDN U17035 ( .A(n16472), .B(n17479), .Z(n16473) );
  NAND U17036 ( .A(n16474), .B(n16473), .Z(n16482) );
  XNOR U17037 ( .A(n16476), .B(n16475), .Z(n16477) );
  NAND U17038 ( .A(n16477), .B(n17458), .Z(n16480) );
  NANDN U17039 ( .A(n2967), .B(x[26]), .Z(n16478) );
  NAND U17040 ( .A(n16480), .B(n16479), .Z(n16481) );
  NOR U17041 ( .A(n16482), .B(n16481), .Z(n16484) );
  NANDN U17042 ( .A(n3020), .B(n17467), .Z(n16483) );
  NAND U17043 ( .A(n16484), .B(n16483), .Z(n2430) );
  NANDN U17044 ( .A(n2967), .B(\stack[6][25] ), .Z(n16486) );
  NANDN U17045 ( .A(n17471), .B(\stack[7][25] ), .Z(n16485) );
  NAND U17046 ( .A(n16486), .B(n16485), .Z(n2431) );
  NANDN U17047 ( .A(n2967), .B(\stack[5][25] ), .Z(n16488) );
  NANDN U17048 ( .A(n17472), .B(\stack[7][25] ), .Z(n16487) );
  AND U17049 ( .A(n16488), .B(n16487), .Z(n16490) );
  NANDN U17050 ( .A(n17475), .B(\stack[6][25] ), .Z(n16489) );
  NAND U17051 ( .A(n16490), .B(n16489), .Z(n2432) );
  NANDN U17052 ( .A(n2967), .B(\stack[4][25] ), .Z(n16492) );
  NANDN U17053 ( .A(n17472), .B(\stack[6][25] ), .Z(n16491) );
  AND U17054 ( .A(n16492), .B(n16491), .Z(n16494) );
  NANDN U17055 ( .A(n17475), .B(\stack[5][25] ), .Z(n16493) );
  NAND U17056 ( .A(n16494), .B(n16493), .Z(n2433) );
  NANDN U17057 ( .A(n2967), .B(\stack[3][25] ), .Z(n16496) );
  NANDN U17058 ( .A(n17472), .B(\stack[5][25] ), .Z(n16495) );
  AND U17059 ( .A(n16496), .B(n16495), .Z(n16498) );
  NANDN U17060 ( .A(n17475), .B(\stack[4][25] ), .Z(n16497) );
  NAND U17061 ( .A(n16498), .B(n16497), .Z(n2434) );
  NANDN U17062 ( .A(n2967), .B(\stack[2][25] ), .Z(n16500) );
  NANDN U17063 ( .A(n17472), .B(\stack[4][25] ), .Z(n16499) );
  AND U17064 ( .A(n16500), .B(n16499), .Z(n16502) );
  NANDN U17065 ( .A(n17475), .B(\stack[3][25] ), .Z(n16501) );
  NAND U17066 ( .A(n16502), .B(n16501), .Z(n2435) );
  NANDN U17067 ( .A(n2982), .B(n17471), .Z(n16504) );
  NANDN U17068 ( .A(n17472), .B(\stack[3][25] ), .Z(n16503) );
  AND U17069 ( .A(n16504), .B(n16503), .Z(n16506) );
  NANDN U17070 ( .A(n17475), .B(\stack[2][25] ), .Z(n16505) );
  NAND U17071 ( .A(n16506), .B(n16505), .Z(n2436) );
  NANDN U17072 ( .A(n3019), .B(n17471), .Z(n16508) );
  NANDN U17073 ( .A(n17472), .B(\stack[2][25] ), .Z(n16507) );
  AND U17074 ( .A(n16508), .B(n16507), .Z(n16510) );
  OR U17075 ( .A(n17475), .B(n2982), .Z(n16509) );
  NAND U17076 ( .A(n16510), .B(n16509), .Z(n2437) );
  XNOR U17077 ( .A(n16512), .B(n16511), .Z(n16513) );
  NAND U17078 ( .A(n16513), .B(n17458), .Z(n16518) );
  NANDN U17079 ( .A(n2967), .B(x[25]), .Z(n16516) );
  NAND U17080 ( .A(n16514), .B(n17479), .Z(n16515) );
  NAND U17081 ( .A(n16516), .B(n16515), .Z(n16517) );
  ANDN U17082 ( .B(n16518), .A(n16517), .Z(n16522) );
  NANDN U17083 ( .A(n17483), .B(\stack[1][25] ), .Z(n16519) );
  NANDN U17084 ( .A(o[25]), .B(n16519), .Z(n16520) );
  ANDN U17085 ( .B(n16520), .A(n17481), .Z(n16521) );
  ANDN U17086 ( .B(n16522), .A(n16521), .Z(n16523) );
  NANDN U17087 ( .A(n2967), .B(\stack[6][24] ), .Z(n16525) );
  NANDN U17088 ( .A(n17471), .B(\stack[7][24] ), .Z(n16524) );
  NAND U17089 ( .A(n16525), .B(n16524), .Z(n2439) );
  NANDN U17090 ( .A(n2967), .B(\stack[5][24] ), .Z(n16527) );
  NANDN U17091 ( .A(n17472), .B(\stack[7][24] ), .Z(n16526) );
  AND U17092 ( .A(n16527), .B(n16526), .Z(n16529) );
  NANDN U17093 ( .A(n17475), .B(\stack[6][24] ), .Z(n16528) );
  NAND U17094 ( .A(n16529), .B(n16528), .Z(n2440) );
  NANDN U17095 ( .A(n2967), .B(\stack[4][24] ), .Z(n16531) );
  NANDN U17096 ( .A(n17472), .B(\stack[6][24] ), .Z(n16530) );
  AND U17097 ( .A(n16531), .B(n16530), .Z(n16533) );
  NANDN U17098 ( .A(n17475), .B(\stack[5][24] ), .Z(n16532) );
  NAND U17099 ( .A(n16533), .B(n16532), .Z(n2441) );
  NANDN U17100 ( .A(n2967), .B(\stack[3][24] ), .Z(n16535) );
  NANDN U17101 ( .A(n17472), .B(\stack[5][24] ), .Z(n16534) );
  AND U17102 ( .A(n16535), .B(n16534), .Z(n16537) );
  NANDN U17103 ( .A(n17475), .B(\stack[4][24] ), .Z(n16536) );
  NAND U17104 ( .A(n16537), .B(n16536), .Z(n2442) );
  NANDN U17105 ( .A(n2967), .B(\stack[2][24] ), .Z(n16539) );
  NANDN U17106 ( .A(n17472), .B(\stack[4][24] ), .Z(n16538) );
  AND U17107 ( .A(n16539), .B(n16538), .Z(n16541) );
  NANDN U17108 ( .A(n17475), .B(\stack[3][24] ), .Z(n16540) );
  NAND U17109 ( .A(n16541), .B(n16540), .Z(n2443) );
  NANDN U17110 ( .A(n2981), .B(n17471), .Z(n16543) );
  NANDN U17111 ( .A(n17472), .B(\stack[3][24] ), .Z(n16542) );
  AND U17112 ( .A(n16543), .B(n16542), .Z(n16545) );
  NANDN U17113 ( .A(n17475), .B(\stack[2][24] ), .Z(n16544) );
  NAND U17114 ( .A(n16545), .B(n16544), .Z(n2444) );
  NANDN U17115 ( .A(n3018), .B(n17471), .Z(n16547) );
  NANDN U17116 ( .A(n17472), .B(\stack[2][24] ), .Z(n16546) );
  AND U17117 ( .A(n16547), .B(n16546), .Z(n16549) );
  OR U17118 ( .A(n17475), .B(n2981), .Z(n16548) );
  NAND U17119 ( .A(n16549), .B(n16548), .Z(n2445) );
  NANDN U17120 ( .A(n2967), .B(x[24]), .Z(n16551) );
  NANDN U17121 ( .A(n17483), .B(\stack[1][24] ), .Z(n16550) );
  NAND U17122 ( .A(n16551), .B(n16550), .Z(n16560) );
  XNOR U17123 ( .A(n16553), .B(n16552), .Z(n16554) );
  NAND U17124 ( .A(n16554), .B(n17458), .Z(n16558) );
  NAND U17125 ( .A(n16555), .B(n17479), .Z(n16556) );
  NAND U17126 ( .A(n16558), .B(n16557), .Z(n16559) );
  NOR U17127 ( .A(n16560), .B(n16559), .Z(n16562) );
  NANDN U17128 ( .A(n3018), .B(n17467), .Z(n16561) );
  NAND U17129 ( .A(n16562), .B(n16561), .Z(n2446) );
  NANDN U17130 ( .A(n2967), .B(\stack[6][23] ), .Z(n16564) );
  NANDN U17131 ( .A(n17471), .B(\stack[7][23] ), .Z(n16563) );
  NAND U17132 ( .A(n16564), .B(n16563), .Z(n2447) );
  NANDN U17133 ( .A(n2967), .B(\stack[5][23] ), .Z(n16566) );
  NANDN U17134 ( .A(n17472), .B(\stack[7][23] ), .Z(n16565) );
  AND U17135 ( .A(n16566), .B(n16565), .Z(n16568) );
  NANDN U17136 ( .A(n17475), .B(\stack[6][23] ), .Z(n16567) );
  NAND U17137 ( .A(n16568), .B(n16567), .Z(n2448) );
  NANDN U17138 ( .A(n2967), .B(\stack[4][23] ), .Z(n16570) );
  NANDN U17139 ( .A(n17472), .B(\stack[6][23] ), .Z(n16569) );
  AND U17140 ( .A(n16570), .B(n16569), .Z(n16572) );
  NANDN U17141 ( .A(n17475), .B(\stack[5][23] ), .Z(n16571) );
  NAND U17142 ( .A(n16572), .B(n16571), .Z(n2449) );
  NANDN U17143 ( .A(n2967), .B(\stack[3][23] ), .Z(n16574) );
  NANDN U17144 ( .A(n17472), .B(\stack[5][23] ), .Z(n16573) );
  AND U17145 ( .A(n16574), .B(n16573), .Z(n16576) );
  NANDN U17146 ( .A(n17475), .B(\stack[4][23] ), .Z(n16575) );
  NAND U17147 ( .A(n16576), .B(n16575), .Z(n2450) );
  NANDN U17148 ( .A(n2967), .B(\stack[2][23] ), .Z(n16578) );
  NANDN U17149 ( .A(n17472), .B(\stack[4][23] ), .Z(n16577) );
  AND U17150 ( .A(n16578), .B(n16577), .Z(n16580) );
  NANDN U17151 ( .A(n17475), .B(\stack[3][23] ), .Z(n16579) );
  NAND U17152 ( .A(n16580), .B(n16579), .Z(n2451) );
  NANDN U17153 ( .A(n2980), .B(n17471), .Z(n16582) );
  NANDN U17154 ( .A(n17472), .B(\stack[3][23] ), .Z(n16581) );
  AND U17155 ( .A(n16582), .B(n16581), .Z(n16584) );
  NANDN U17156 ( .A(n17475), .B(\stack[2][23] ), .Z(n16583) );
  NAND U17157 ( .A(n16584), .B(n16583), .Z(n2452) );
  NANDN U17158 ( .A(n3017), .B(n17471), .Z(n16586) );
  NANDN U17159 ( .A(n17472), .B(\stack[2][23] ), .Z(n16585) );
  AND U17160 ( .A(n16586), .B(n16585), .Z(n16588) );
  OR U17161 ( .A(n17475), .B(n2980), .Z(n16587) );
  NAND U17162 ( .A(n16588), .B(n16587), .Z(n2453) );
  NANDN U17163 ( .A(n2967), .B(x[23]), .Z(n16591) );
  NAND U17164 ( .A(n16589), .B(n17479), .Z(n16590) );
  NAND U17165 ( .A(n16591), .B(n16590), .Z(n16599) );
  XNOR U17166 ( .A(n16593), .B(n16592), .Z(n16594) );
  NAND U17167 ( .A(n16594), .B(n17458), .Z(n16597) );
  NANDN U17168 ( .A(n2980), .B(n17461), .Z(n16595) );
  NAND U17169 ( .A(n16597), .B(n16596), .Z(n16598) );
  NOR U17170 ( .A(n16599), .B(n16598), .Z(n16601) );
  NANDN U17171 ( .A(n3017), .B(n17467), .Z(n16600) );
  NAND U17172 ( .A(n16601), .B(n16600), .Z(n2454) );
  NANDN U17173 ( .A(n2967), .B(\stack[6][22] ), .Z(n16603) );
  NANDN U17174 ( .A(n17471), .B(\stack[7][22] ), .Z(n16602) );
  NAND U17175 ( .A(n16603), .B(n16602), .Z(n2455) );
  NANDN U17176 ( .A(n2967), .B(\stack[5][22] ), .Z(n16605) );
  NANDN U17177 ( .A(n17472), .B(\stack[7][22] ), .Z(n16604) );
  AND U17178 ( .A(n16605), .B(n16604), .Z(n16607) );
  NANDN U17179 ( .A(n17475), .B(\stack[6][22] ), .Z(n16606) );
  NAND U17180 ( .A(n16607), .B(n16606), .Z(n2456) );
  NANDN U17181 ( .A(n2967), .B(\stack[4][22] ), .Z(n16609) );
  NANDN U17182 ( .A(n17472), .B(\stack[6][22] ), .Z(n16608) );
  AND U17183 ( .A(n16609), .B(n16608), .Z(n16611) );
  NANDN U17184 ( .A(n17475), .B(\stack[5][22] ), .Z(n16610) );
  NAND U17185 ( .A(n16611), .B(n16610), .Z(n2457) );
  NANDN U17186 ( .A(n2967), .B(\stack[3][22] ), .Z(n16613) );
  NANDN U17187 ( .A(n17472), .B(\stack[5][22] ), .Z(n16612) );
  AND U17188 ( .A(n16613), .B(n16612), .Z(n16615) );
  NANDN U17189 ( .A(n17475), .B(\stack[4][22] ), .Z(n16614) );
  NAND U17190 ( .A(n16615), .B(n16614), .Z(n2458) );
  NANDN U17191 ( .A(n2967), .B(\stack[2][22] ), .Z(n16617) );
  NANDN U17192 ( .A(n17472), .B(\stack[4][22] ), .Z(n16616) );
  AND U17193 ( .A(n16617), .B(n16616), .Z(n16619) );
  NANDN U17194 ( .A(n17475), .B(\stack[3][22] ), .Z(n16618) );
  NAND U17195 ( .A(n16619), .B(n16618), .Z(n2459) );
  NANDN U17196 ( .A(n2979), .B(n17471), .Z(n16621) );
  NANDN U17197 ( .A(n17472), .B(\stack[3][22] ), .Z(n16620) );
  AND U17198 ( .A(n16621), .B(n16620), .Z(n16623) );
  NANDN U17199 ( .A(n17475), .B(\stack[2][22] ), .Z(n16622) );
  NAND U17200 ( .A(n16623), .B(n16622), .Z(n2460) );
  NANDN U17201 ( .A(n3016), .B(n17471), .Z(n16625) );
  NANDN U17202 ( .A(n17472), .B(\stack[2][22] ), .Z(n16624) );
  AND U17203 ( .A(n16625), .B(n16624), .Z(n16627) );
  OR U17204 ( .A(n17475), .B(n2979), .Z(n16626) );
  NAND U17205 ( .A(n16627), .B(n16626), .Z(n2461) );
  NANDN U17206 ( .A(n2967), .B(x[22]), .Z(n16629) );
  NANDN U17207 ( .A(n17483), .B(\stack[1][22] ), .Z(n16628) );
  NAND U17208 ( .A(n16629), .B(n16628), .Z(n16638) );
  XNOR U17209 ( .A(n16631), .B(n16630), .Z(n16632) );
  NAND U17210 ( .A(n16632), .B(n17458), .Z(n16636) );
  NANDN U17211 ( .A(n16633), .B(n17479), .Z(n16634) );
  NAND U17212 ( .A(n16636), .B(n16635), .Z(n16637) );
  NOR U17213 ( .A(n16638), .B(n16637), .Z(n16640) );
  NANDN U17214 ( .A(n3016), .B(n17467), .Z(n16639) );
  NAND U17215 ( .A(n16640), .B(n16639), .Z(n2462) );
  NANDN U17216 ( .A(n2967), .B(\stack[6][21] ), .Z(n16642) );
  NANDN U17217 ( .A(n17471), .B(\stack[7][21] ), .Z(n16641) );
  NAND U17218 ( .A(n16642), .B(n16641), .Z(n2463) );
  NANDN U17219 ( .A(n2967), .B(\stack[5][21] ), .Z(n16644) );
  NANDN U17220 ( .A(n17472), .B(\stack[7][21] ), .Z(n16643) );
  AND U17221 ( .A(n16644), .B(n16643), .Z(n16646) );
  NANDN U17222 ( .A(n17475), .B(\stack[6][21] ), .Z(n16645) );
  NAND U17223 ( .A(n16646), .B(n16645), .Z(n2464) );
  NANDN U17224 ( .A(n2967), .B(\stack[4][21] ), .Z(n16648) );
  NANDN U17225 ( .A(n17472), .B(\stack[6][21] ), .Z(n16647) );
  AND U17226 ( .A(n16648), .B(n16647), .Z(n16650) );
  NANDN U17227 ( .A(n17475), .B(\stack[5][21] ), .Z(n16649) );
  NAND U17228 ( .A(n16650), .B(n16649), .Z(n2465) );
  NANDN U17229 ( .A(n2967), .B(\stack[3][21] ), .Z(n16652) );
  NANDN U17230 ( .A(n17472), .B(\stack[5][21] ), .Z(n16651) );
  AND U17231 ( .A(n16652), .B(n16651), .Z(n16654) );
  NANDN U17232 ( .A(n17475), .B(\stack[4][21] ), .Z(n16653) );
  NAND U17233 ( .A(n16654), .B(n16653), .Z(n2466) );
  NANDN U17234 ( .A(n2967), .B(\stack[2][21] ), .Z(n16656) );
  NANDN U17235 ( .A(n17472), .B(\stack[4][21] ), .Z(n16655) );
  AND U17236 ( .A(n16656), .B(n16655), .Z(n16658) );
  NANDN U17237 ( .A(n17475), .B(\stack[3][21] ), .Z(n16657) );
  NAND U17238 ( .A(n16658), .B(n16657), .Z(n2467) );
  NANDN U17239 ( .A(n2978), .B(n17471), .Z(n16660) );
  NANDN U17240 ( .A(n17472), .B(\stack[3][21] ), .Z(n16659) );
  AND U17241 ( .A(n16660), .B(n16659), .Z(n16662) );
  NANDN U17242 ( .A(n17475), .B(\stack[2][21] ), .Z(n16661) );
  NAND U17243 ( .A(n16662), .B(n16661), .Z(n2468) );
  NANDN U17244 ( .A(n3015), .B(n17471), .Z(n16664) );
  NANDN U17245 ( .A(n17472), .B(\stack[2][21] ), .Z(n16663) );
  AND U17246 ( .A(n16664), .B(n16663), .Z(n16666) );
  OR U17247 ( .A(n17475), .B(n2978), .Z(n16665) );
  NAND U17248 ( .A(n16666), .B(n16665), .Z(n2469) );
  NANDN U17249 ( .A(n2967), .B(x[21]), .Z(n16668) );
  NANDN U17250 ( .A(n17483), .B(\stack[1][21] ), .Z(n16667) );
  NAND U17251 ( .A(n16668), .B(n16667), .Z(n16677) );
  XNOR U17252 ( .A(n16670), .B(n16669), .Z(n16671) );
  NAND U17253 ( .A(n16671), .B(n17458), .Z(n16675) );
  NAND U17254 ( .A(n16672), .B(n17479), .Z(n16673) );
  NAND U17255 ( .A(n16675), .B(n16674), .Z(n16676) );
  NOR U17256 ( .A(n16677), .B(n16676), .Z(n16679) );
  NANDN U17257 ( .A(n3015), .B(n17467), .Z(n16678) );
  NAND U17258 ( .A(n16679), .B(n16678), .Z(n2470) );
  NANDN U17259 ( .A(n2967), .B(\stack[6][20] ), .Z(n16681) );
  NANDN U17260 ( .A(n17471), .B(\stack[7][20] ), .Z(n16680) );
  NAND U17261 ( .A(n16681), .B(n16680), .Z(n2471) );
  NANDN U17262 ( .A(n2967), .B(\stack[5][20] ), .Z(n16683) );
  NANDN U17263 ( .A(n17472), .B(\stack[7][20] ), .Z(n16682) );
  AND U17264 ( .A(n16683), .B(n16682), .Z(n16685) );
  NANDN U17265 ( .A(n17475), .B(\stack[6][20] ), .Z(n16684) );
  NAND U17266 ( .A(n16685), .B(n16684), .Z(n2472) );
  NANDN U17267 ( .A(n2967), .B(\stack[4][20] ), .Z(n16687) );
  NANDN U17268 ( .A(n17472), .B(\stack[6][20] ), .Z(n16686) );
  AND U17269 ( .A(n16687), .B(n16686), .Z(n16689) );
  NANDN U17270 ( .A(n17475), .B(\stack[5][20] ), .Z(n16688) );
  NAND U17271 ( .A(n16689), .B(n16688), .Z(n2473) );
  NANDN U17272 ( .A(n2967), .B(\stack[3][20] ), .Z(n16691) );
  NANDN U17273 ( .A(n17472), .B(\stack[5][20] ), .Z(n16690) );
  AND U17274 ( .A(n16691), .B(n16690), .Z(n16693) );
  NANDN U17275 ( .A(n17475), .B(\stack[4][20] ), .Z(n16692) );
  NAND U17276 ( .A(n16693), .B(n16692), .Z(n2474) );
  NANDN U17277 ( .A(n2967), .B(\stack[2][20] ), .Z(n16695) );
  NANDN U17278 ( .A(n17472), .B(\stack[4][20] ), .Z(n16694) );
  AND U17279 ( .A(n16695), .B(n16694), .Z(n16697) );
  NANDN U17280 ( .A(n17475), .B(\stack[3][20] ), .Z(n16696) );
  NAND U17281 ( .A(n16697), .B(n16696), .Z(n2475) );
  NANDN U17282 ( .A(n16712), .B(n17471), .Z(n16699) );
  NANDN U17283 ( .A(n17472), .B(\stack[3][20] ), .Z(n16698) );
  AND U17284 ( .A(n16699), .B(n16698), .Z(n16701) );
  NANDN U17285 ( .A(n17475), .B(\stack[2][20] ), .Z(n16700) );
  NAND U17286 ( .A(n16701), .B(n16700), .Z(n2476) );
  NANDN U17287 ( .A(n3014), .B(n17471), .Z(n16703) );
  NANDN U17288 ( .A(n17472), .B(\stack[2][20] ), .Z(n16702) );
  AND U17289 ( .A(n16703), .B(n16702), .Z(n16705) );
  OR U17290 ( .A(n17475), .B(n16712), .Z(n16704) );
  NAND U17291 ( .A(n16705), .B(n16704), .Z(n2477) );
  NANDN U17292 ( .A(n2967), .B(x[20]), .Z(n16708) );
  NANDN U17293 ( .A(n16706), .B(n17479), .Z(n16707) );
  NAND U17294 ( .A(n16708), .B(n16707), .Z(n16717) );
  XNOR U17295 ( .A(n16710), .B(n16709), .Z(n16711) );
  NAND U17296 ( .A(n16711), .B(n17458), .Z(n16715) );
  NANDN U17297 ( .A(n16712), .B(n17461), .Z(n16713) );
  NAND U17298 ( .A(n16715), .B(n16714), .Z(n16716) );
  NOR U17299 ( .A(n16717), .B(n16716), .Z(n16719) );
  NANDN U17300 ( .A(n3014), .B(n17467), .Z(n16718) );
  NAND U17301 ( .A(n16719), .B(n16718), .Z(n2478) );
  NANDN U17302 ( .A(n2967), .B(\stack[6][19] ), .Z(n16721) );
  NANDN U17303 ( .A(n17471), .B(\stack[7][19] ), .Z(n16720) );
  NAND U17304 ( .A(n16721), .B(n16720), .Z(n2479) );
  NANDN U17305 ( .A(n2967), .B(\stack[5][19] ), .Z(n16723) );
  NANDN U17306 ( .A(n17472), .B(\stack[7][19] ), .Z(n16722) );
  AND U17307 ( .A(n16723), .B(n16722), .Z(n16725) );
  NANDN U17308 ( .A(n17475), .B(\stack[6][19] ), .Z(n16724) );
  NAND U17309 ( .A(n16725), .B(n16724), .Z(n2480) );
  NANDN U17310 ( .A(n2967), .B(\stack[4][19] ), .Z(n16727) );
  NANDN U17311 ( .A(n17472), .B(\stack[6][19] ), .Z(n16726) );
  AND U17312 ( .A(n16727), .B(n16726), .Z(n16729) );
  NANDN U17313 ( .A(n17475), .B(\stack[5][19] ), .Z(n16728) );
  NAND U17314 ( .A(n16729), .B(n16728), .Z(n2481) );
  NANDN U17315 ( .A(n2967), .B(\stack[3][19] ), .Z(n16731) );
  NANDN U17316 ( .A(n17472), .B(\stack[5][19] ), .Z(n16730) );
  AND U17317 ( .A(n16731), .B(n16730), .Z(n16733) );
  NANDN U17318 ( .A(n17475), .B(\stack[4][19] ), .Z(n16732) );
  NAND U17319 ( .A(n16733), .B(n16732), .Z(n2482) );
  NANDN U17320 ( .A(n2967), .B(\stack[2][19] ), .Z(n16735) );
  NANDN U17321 ( .A(n17472), .B(\stack[4][19] ), .Z(n16734) );
  AND U17322 ( .A(n16735), .B(n16734), .Z(n16737) );
  NANDN U17323 ( .A(n17475), .B(\stack[3][19] ), .Z(n16736) );
  NAND U17324 ( .A(n16737), .B(n16736), .Z(n2483) );
  NANDN U17325 ( .A(n16746), .B(n17471), .Z(n16739) );
  NANDN U17326 ( .A(n17472), .B(\stack[3][19] ), .Z(n16738) );
  AND U17327 ( .A(n16739), .B(n16738), .Z(n16741) );
  NANDN U17328 ( .A(n17475), .B(\stack[2][19] ), .Z(n16740) );
  NAND U17329 ( .A(n16741), .B(n16740), .Z(n2484) );
  NANDN U17330 ( .A(n3013), .B(n17471), .Z(n16743) );
  NANDN U17331 ( .A(n17472), .B(\stack[2][19] ), .Z(n16742) );
  AND U17332 ( .A(n16743), .B(n16742), .Z(n16745) );
  OR U17333 ( .A(n17475), .B(n16746), .Z(n16744) );
  NAND U17334 ( .A(n16745), .B(n16744), .Z(n2485) );
  NANDN U17335 ( .A(n16746), .B(n17461), .Z(n16749) );
  NAND U17336 ( .A(n16747), .B(n17479), .Z(n16748) );
  NAND U17337 ( .A(n16749), .B(n16748), .Z(n16757) );
  XNOR U17338 ( .A(n16751), .B(n16750), .Z(n16752) );
  NAND U17339 ( .A(n16752), .B(n17458), .Z(n16755) );
  NANDN U17340 ( .A(n2967), .B(x[19]), .Z(n16753) );
  NAND U17341 ( .A(n16755), .B(n16754), .Z(n16756) );
  NOR U17342 ( .A(n16757), .B(n16756), .Z(n16759) );
  NANDN U17343 ( .A(n3013), .B(n17467), .Z(n16758) );
  NAND U17344 ( .A(n16759), .B(n16758), .Z(n2486) );
  NANDN U17345 ( .A(n2967), .B(\stack[6][18] ), .Z(n16761) );
  NANDN U17346 ( .A(n17471), .B(\stack[7][18] ), .Z(n16760) );
  NAND U17347 ( .A(n16761), .B(n16760), .Z(n2487) );
  NANDN U17348 ( .A(n2967), .B(\stack[5][18] ), .Z(n16763) );
  NANDN U17349 ( .A(n17472), .B(\stack[7][18] ), .Z(n16762) );
  AND U17350 ( .A(n16763), .B(n16762), .Z(n16765) );
  NANDN U17351 ( .A(n17475), .B(\stack[6][18] ), .Z(n16764) );
  NAND U17352 ( .A(n16765), .B(n16764), .Z(n2488) );
  NANDN U17353 ( .A(n2967), .B(\stack[4][18] ), .Z(n16767) );
  NANDN U17354 ( .A(n17472), .B(\stack[6][18] ), .Z(n16766) );
  AND U17355 ( .A(n16767), .B(n16766), .Z(n16769) );
  NANDN U17356 ( .A(n17475), .B(\stack[5][18] ), .Z(n16768) );
  NAND U17357 ( .A(n16769), .B(n16768), .Z(n2489) );
  NANDN U17358 ( .A(n2967), .B(\stack[3][18] ), .Z(n16771) );
  NANDN U17359 ( .A(n17472), .B(\stack[5][18] ), .Z(n16770) );
  AND U17360 ( .A(n16771), .B(n16770), .Z(n16773) );
  NANDN U17361 ( .A(n17475), .B(\stack[4][18] ), .Z(n16772) );
  NAND U17362 ( .A(n16773), .B(n16772), .Z(n2490) );
  NANDN U17363 ( .A(n2967), .B(\stack[2][18] ), .Z(n16775) );
  NANDN U17364 ( .A(n17472), .B(\stack[4][18] ), .Z(n16774) );
  AND U17365 ( .A(n16775), .B(n16774), .Z(n16777) );
  NANDN U17366 ( .A(n17475), .B(\stack[3][18] ), .Z(n16776) );
  NAND U17367 ( .A(n16777), .B(n16776), .Z(n2491) );
  NANDN U17368 ( .A(n16786), .B(n17471), .Z(n16779) );
  NANDN U17369 ( .A(n17472), .B(\stack[3][18] ), .Z(n16778) );
  AND U17370 ( .A(n16779), .B(n16778), .Z(n16781) );
  NANDN U17371 ( .A(n17475), .B(\stack[2][18] ), .Z(n16780) );
  NAND U17372 ( .A(n16781), .B(n16780), .Z(n2492) );
  NANDN U17373 ( .A(n3012), .B(n17471), .Z(n16783) );
  NANDN U17374 ( .A(n17472), .B(\stack[2][18] ), .Z(n16782) );
  AND U17375 ( .A(n16783), .B(n16782), .Z(n16785) );
  OR U17376 ( .A(n17475), .B(n16786), .Z(n16784) );
  NAND U17377 ( .A(n16785), .B(n16784), .Z(n2493) );
  NANDN U17378 ( .A(n16786), .B(n17461), .Z(n16789) );
  NANDN U17379 ( .A(n16787), .B(n17479), .Z(n16788) );
  NAND U17380 ( .A(n16789), .B(n16788), .Z(n16797) );
  XNOR U17381 ( .A(n16791), .B(n16790), .Z(n16792) );
  NAND U17382 ( .A(n16792), .B(n17458), .Z(n16795) );
  NANDN U17383 ( .A(n2967), .B(x[18]), .Z(n16793) );
  NAND U17384 ( .A(n16795), .B(n16794), .Z(n16796) );
  NOR U17385 ( .A(n16797), .B(n16796), .Z(n16799) );
  NANDN U17386 ( .A(n3012), .B(n17467), .Z(n16798) );
  NAND U17387 ( .A(n16799), .B(n16798), .Z(n2494) );
  NANDN U17388 ( .A(n2967), .B(\stack[6][17] ), .Z(n16801) );
  NANDN U17389 ( .A(n17471), .B(\stack[7][17] ), .Z(n16800) );
  NAND U17390 ( .A(n16801), .B(n16800), .Z(n2495) );
  NANDN U17391 ( .A(n2967), .B(\stack[5][17] ), .Z(n16803) );
  NANDN U17392 ( .A(n17472), .B(\stack[7][17] ), .Z(n16802) );
  AND U17393 ( .A(n16803), .B(n16802), .Z(n16805) );
  NANDN U17394 ( .A(n17475), .B(\stack[6][17] ), .Z(n16804) );
  NAND U17395 ( .A(n16805), .B(n16804), .Z(n2496) );
  NANDN U17396 ( .A(n2967), .B(\stack[4][17] ), .Z(n16807) );
  NANDN U17397 ( .A(n17472), .B(\stack[6][17] ), .Z(n16806) );
  AND U17398 ( .A(n16807), .B(n16806), .Z(n16809) );
  NANDN U17399 ( .A(n17475), .B(\stack[5][17] ), .Z(n16808) );
  NAND U17400 ( .A(n16809), .B(n16808), .Z(n2497) );
  NANDN U17401 ( .A(n2967), .B(\stack[3][17] ), .Z(n16811) );
  NANDN U17402 ( .A(n17472), .B(\stack[5][17] ), .Z(n16810) );
  AND U17403 ( .A(n16811), .B(n16810), .Z(n16813) );
  NANDN U17404 ( .A(n17475), .B(\stack[4][17] ), .Z(n16812) );
  NAND U17405 ( .A(n16813), .B(n16812), .Z(n2498) );
  NANDN U17406 ( .A(n2967), .B(\stack[2][17] ), .Z(n16815) );
  NANDN U17407 ( .A(n17472), .B(\stack[4][17] ), .Z(n16814) );
  AND U17408 ( .A(n16815), .B(n16814), .Z(n16817) );
  NANDN U17409 ( .A(n17475), .B(\stack[3][17] ), .Z(n16816) );
  NAND U17410 ( .A(n16817), .B(n16816), .Z(n2499) );
  NANDN U17411 ( .A(n16826), .B(n17471), .Z(n16819) );
  NANDN U17412 ( .A(n17472), .B(\stack[3][17] ), .Z(n16818) );
  AND U17413 ( .A(n16819), .B(n16818), .Z(n16821) );
  NANDN U17414 ( .A(n17475), .B(\stack[2][17] ), .Z(n16820) );
  NAND U17415 ( .A(n16821), .B(n16820), .Z(n2500) );
  NANDN U17416 ( .A(n3011), .B(n17471), .Z(n16823) );
  NANDN U17417 ( .A(n17472), .B(\stack[2][17] ), .Z(n16822) );
  AND U17418 ( .A(n16823), .B(n16822), .Z(n16825) );
  OR U17419 ( .A(n17475), .B(n16826), .Z(n16824) );
  NAND U17420 ( .A(n16825), .B(n16824), .Z(n2501) );
  NANDN U17421 ( .A(n16826), .B(n17461), .Z(n16829) );
  NAND U17422 ( .A(n16827), .B(n17479), .Z(n16828) );
  NAND U17423 ( .A(n16829), .B(n16828), .Z(n16837) );
  XNOR U17424 ( .A(n16831), .B(n16830), .Z(n16832) );
  NAND U17425 ( .A(n16832), .B(n17458), .Z(n16835) );
  NANDN U17426 ( .A(n2967), .B(x[17]), .Z(n16833) );
  NAND U17427 ( .A(n16835), .B(n16834), .Z(n16836) );
  NOR U17428 ( .A(n16837), .B(n16836), .Z(n16839) );
  NANDN U17429 ( .A(n3011), .B(n17467), .Z(n16838) );
  NAND U17430 ( .A(n16839), .B(n16838), .Z(n2502) );
  NANDN U17431 ( .A(n2967), .B(\stack[6][16] ), .Z(n16841) );
  NANDN U17432 ( .A(n17471), .B(\stack[7][16] ), .Z(n16840) );
  NAND U17433 ( .A(n16841), .B(n16840), .Z(n2503) );
  NANDN U17434 ( .A(n2967), .B(\stack[5][16] ), .Z(n16843) );
  NANDN U17435 ( .A(n17472), .B(\stack[7][16] ), .Z(n16842) );
  AND U17436 ( .A(n16843), .B(n16842), .Z(n16845) );
  NANDN U17437 ( .A(n17475), .B(\stack[6][16] ), .Z(n16844) );
  NAND U17438 ( .A(n16845), .B(n16844), .Z(n2504) );
  NANDN U17439 ( .A(n2967), .B(\stack[4][16] ), .Z(n16847) );
  NANDN U17440 ( .A(n17472), .B(\stack[6][16] ), .Z(n16846) );
  AND U17441 ( .A(n16847), .B(n16846), .Z(n16849) );
  NANDN U17442 ( .A(n17475), .B(\stack[5][16] ), .Z(n16848) );
  NAND U17443 ( .A(n16849), .B(n16848), .Z(n2505) );
  NANDN U17444 ( .A(n2967), .B(\stack[3][16] ), .Z(n16851) );
  NANDN U17445 ( .A(n17472), .B(\stack[5][16] ), .Z(n16850) );
  AND U17446 ( .A(n16851), .B(n16850), .Z(n16853) );
  NANDN U17447 ( .A(n17475), .B(\stack[4][16] ), .Z(n16852) );
  NAND U17448 ( .A(n16853), .B(n16852), .Z(n2506) );
  NANDN U17449 ( .A(n2967), .B(\stack[2][16] ), .Z(n16855) );
  NANDN U17450 ( .A(n17472), .B(\stack[4][16] ), .Z(n16854) );
  AND U17451 ( .A(n16855), .B(n16854), .Z(n16857) );
  NANDN U17452 ( .A(n17475), .B(\stack[3][16] ), .Z(n16856) );
  NAND U17453 ( .A(n16857), .B(n16856), .Z(n2507) );
  NANDN U17454 ( .A(n2977), .B(n17471), .Z(n16859) );
  NANDN U17455 ( .A(n17472), .B(\stack[3][16] ), .Z(n16858) );
  AND U17456 ( .A(n16859), .B(n16858), .Z(n16861) );
  NANDN U17457 ( .A(n17475), .B(\stack[2][16] ), .Z(n16860) );
  NAND U17458 ( .A(n16861), .B(n16860), .Z(n2508) );
  NANDN U17459 ( .A(n3010), .B(n17471), .Z(n16863) );
  NANDN U17460 ( .A(n17472), .B(\stack[2][16] ), .Z(n16862) );
  AND U17461 ( .A(n16863), .B(n16862), .Z(n16865) );
  OR U17462 ( .A(n17475), .B(n2977), .Z(n16864) );
  NAND U17463 ( .A(n16865), .B(n16864), .Z(n2509) );
  XNOR U17464 ( .A(n16867), .B(n16866), .Z(n16868) );
  NAND U17465 ( .A(n16868), .B(n17458), .Z(n16873) );
  NANDN U17466 ( .A(n2967), .B(x[16]), .Z(n16871) );
  NANDN U17467 ( .A(n16869), .B(n17479), .Z(n16870) );
  NAND U17468 ( .A(n16871), .B(n16870), .Z(n16872) );
  ANDN U17469 ( .B(n16873), .A(n16872), .Z(n16877) );
  NANDN U17470 ( .A(n17483), .B(\stack[1][16] ), .Z(n16874) );
  NANDN U17471 ( .A(o[16]), .B(n16874), .Z(n16875) );
  ANDN U17472 ( .B(n16875), .A(n17481), .Z(n16876) );
  ANDN U17473 ( .B(n16877), .A(n16876), .Z(n16878) );
  NANDN U17474 ( .A(n2967), .B(\stack[6][15] ), .Z(n16880) );
  NANDN U17475 ( .A(n17471), .B(\stack[7][15] ), .Z(n16879) );
  NAND U17476 ( .A(n16880), .B(n16879), .Z(n2511) );
  NANDN U17477 ( .A(n2967), .B(\stack[5][15] ), .Z(n16882) );
  NANDN U17478 ( .A(n17472), .B(\stack[7][15] ), .Z(n16881) );
  AND U17479 ( .A(n16882), .B(n16881), .Z(n16884) );
  NANDN U17480 ( .A(n17475), .B(\stack[6][15] ), .Z(n16883) );
  NAND U17481 ( .A(n16884), .B(n16883), .Z(n2512) );
  NANDN U17482 ( .A(n2967), .B(\stack[4][15] ), .Z(n16886) );
  NANDN U17483 ( .A(n17472), .B(\stack[6][15] ), .Z(n16885) );
  AND U17484 ( .A(n16886), .B(n16885), .Z(n16888) );
  NANDN U17485 ( .A(n17475), .B(\stack[5][15] ), .Z(n16887) );
  NAND U17486 ( .A(n16888), .B(n16887), .Z(n2513) );
  NANDN U17487 ( .A(n2967), .B(\stack[3][15] ), .Z(n16890) );
  NANDN U17488 ( .A(n17472), .B(\stack[5][15] ), .Z(n16889) );
  AND U17489 ( .A(n16890), .B(n16889), .Z(n16892) );
  NANDN U17490 ( .A(n17475), .B(\stack[4][15] ), .Z(n16891) );
  NAND U17491 ( .A(n16892), .B(n16891), .Z(n2514) );
  NANDN U17492 ( .A(n2967), .B(\stack[2][15] ), .Z(n16894) );
  NANDN U17493 ( .A(n17472), .B(\stack[4][15] ), .Z(n16893) );
  AND U17494 ( .A(n16894), .B(n16893), .Z(n16896) );
  NANDN U17495 ( .A(n17475), .B(\stack[3][15] ), .Z(n16895) );
  NAND U17496 ( .A(n16896), .B(n16895), .Z(n2515) );
  NANDN U17497 ( .A(n2976), .B(n17471), .Z(n16898) );
  NANDN U17498 ( .A(n17472), .B(\stack[3][15] ), .Z(n16897) );
  AND U17499 ( .A(n16898), .B(n16897), .Z(n16900) );
  NANDN U17500 ( .A(n17475), .B(\stack[2][15] ), .Z(n16899) );
  NAND U17501 ( .A(n16900), .B(n16899), .Z(n2516) );
  NANDN U17502 ( .A(n3009), .B(n17471), .Z(n16902) );
  NANDN U17503 ( .A(n17472), .B(\stack[2][15] ), .Z(n16901) );
  AND U17504 ( .A(n16902), .B(n16901), .Z(n16904) );
  OR U17505 ( .A(n17475), .B(n2976), .Z(n16903) );
  NAND U17506 ( .A(n16904), .B(n16903), .Z(n2517) );
  NANDN U17507 ( .A(n2976), .B(n17461), .Z(n16907) );
  NAND U17508 ( .A(n16905), .B(n17479), .Z(n16906) );
  NAND U17509 ( .A(n16907), .B(n16906), .Z(n16915) );
  XNOR U17510 ( .A(n16909), .B(n16908), .Z(n16910) );
  NAND U17511 ( .A(n16910), .B(n17458), .Z(n16913) );
  NANDN U17512 ( .A(n2967), .B(x[15]), .Z(n16911) );
  NAND U17513 ( .A(n16913), .B(n16912), .Z(n16914) );
  NOR U17514 ( .A(n16915), .B(n16914), .Z(n16917) );
  NANDN U17515 ( .A(n3009), .B(n17467), .Z(n16916) );
  NAND U17516 ( .A(n16917), .B(n16916), .Z(n2518) );
  NANDN U17517 ( .A(n2967), .B(\stack[6][14] ), .Z(n16919) );
  NANDN U17518 ( .A(n17471), .B(\stack[7][14] ), .Z(n16918) );
  NAND U17519 ( .A(n16919), .B(n16918), .Z(n2519) );
  NANDN U17520 ( .A(n2967), .B(\stack[5][14] ), .Z(n16921) );
  NANDN U17521 ( .A(n17472), .B(\stack[7][14] ), .Z(n16920) );
  AND U17522 ( .A(n16921), .B(n16920), .Z(n16923) );
  NANDN U17523 ( .A(n17475), .B(\stack[6][14] ), .Z(n16922) );
  NAND U17524 ( .A(n16923), .B(n16922), .Z(n2520) );
  NANDN U17525 ( .A(n2967), .B(\stack[4][14] ), .Z(n16925) );
  NANDN U17526 ( .A(n17472), .B(\stack[6][14] ), .Z(n16924) );
  AND U17527 ( .A(n16925), .B(n16924), .Z(n16927) );
  NANDN U17528 ( .A(n17475), .B(\stack[5][14] ), .Z(n16926) );
  NAND U17529 ( .A(n16927), .B(n16926), .Z(n2521) );
  NANDN U17530 ( .A(n2967), .B(\stack[3][14] ), .Z(n16929) );
  NANDN U17531 ( .A(n17472), .B(\stack[5][14] ), .Z(n16928) );
  AND U17532 ( .A(n16929), .B(n16928), .Z(n16931) );
  NANDN U17533 ( .A(n17475), .B(\stack[4][14] ), .Z(n16930) );
  NAND U17534 ( .A(n16931), .B(n16930), .Z(n2522) );
  NANDN U17535 ( .A(n2967), .B(\stack[2][14] ), .Z(n16933) );
  NANDN U17536 ( .A(n17472), .B(\stack[4][14] ), .Z(n16932) );
  AND U17537 ( .A(n16933), .B(n16932), .Z(n16935) );
  NANDN U17538 ( .A(n17475), .B(\stack[3][14] ), .Z(n16934) );
  NAND U17539 ( .A(n16935), .B(n16934), .Z(n2523) );
  NANDN U17540 ( .A(n2975), .B(n17471), .Z(n16937) );
  NANDN U17541 ( .A(n17472), .B(\stack[3][14] ), .Z(n16936) );
  AND U17542 ( .A(n16937), .B(n16936), .Z(n16939) );
  NANDN U17543 ( .A(n17475), .B(\stack[2][14] ), .Z(n16938) );
  NAND U17544 ( .A(n16939), .B(n16938), .Z(n2524) );
  NANDN U17545 ( .A(n3008), .B(n17471), .Z(n16941) );
  NANDN U17546 ( .A(n17472), .B(\stack[2][14] ), .Z(n16940) );
  AND U17547 ( .A(n16941), .B(n16940), .Z(n16943) );
  OR U17548 ( .A(n17475), .B(n2975), .Z(n16942) );
  NAND U17549 ( .A(n16943), .B(n16942), .Z(n2525) );
  NANDN U17550 ( .A(n2967), .B(x[14]), .Z(n16946) );
  NANDN U17551 ( .A(n16944), .B(n17479), .Z(n16945) );
  NAND U17552 ( .A(n16946), .B(n16945), .Z(n16954) );
  XNOR U17553 ( .A(n16948), .B(n16947), .Z(n16949) );
  NAND U17554 ( .A(n16949), .B(n17458), .Z(n16952) );
  NANDN U17555 ( .A(n2975), .B(n17461), .Z(n16950) );
  NAND U17556 ( .A(n16952), .B(n16951), .Z(n16953) );
  NOR U17557 ( .A(n16954), .B(n16953), .Z(n16956) );
  NANDN U17558 ( .A(n3008), .B(n17467), .Z(n16955) );
  NAND U17559 ( .A(n16956), .B(n16955), .Z(n2526) );
  NANDN U17560 ( .A(n2967), .B(\stack[6][13] ), .Z(n16958) );
  NANDN U17561 ( .A(n17471), .B(\stack[7][13] ), .Z(n16957) );
  NAND U17562 ( .A(n16958), .B(n16957), .Z(n2527) );
  NANDN U17563 ( .A(n2967), .B(\stack[5][13] ), .Z(n16960) );
  NANDN U17564 ( .A(n17472), .B(\stack[7][13] ), .Z(n16959) );
  AND U17565 ( .A(n16960), .B(n16959), .Z(n16962) );
  NANDN U17566 ( .A(n17475), .B(\stack[6][13] ), .Z(n16961) );
  NAND U17567 ( .A(n16962), .B(n16961), .Z(n2528) );
  NANDN U17568 ( .A(n2967), .B(\stack[4][13] ), .Z(n16964) );
  NANDN U17569 ( .A(n17472), .B(\stack[6][13] ), .Z(n16963) );
  AND U17570 ( .A(n16964), .B(n16963), .Z(n16966) );
  NANDN U17571 ( .A(n17475), .B(\stack[5][13] ), .Z(n16965) );
  NAND U17572 ( .A(n16966), .B(n16965), .Z(n2529) );
  NANDN U17573 ( .A(n2967), .B(\stack[3][13] ), .Z(n16968) );
  NANDN U17574 ( .A(n17472), .B(\stack[5][13] ), .Z(n16967) );
  AND U17575 ( .A(n16968), .B(n16967), .Z(n16970) );
  NANDN U17576 ( .A(n17475), .B(\stack[4][13] ), .Z(n16969) );
  NAND U17577 ( .A(n16970), .B(n16969), .Z(n2530) );
  NANDN U17578 ( .A(n2967), .B(\stack[2][13] ), .Z(n16972) );
  NANDN U17579 ( .A(n17472), .B(\stack[4][13] ), .Z(n16971) );
  AND U17580 ( .A(n16972), .B(n16971), .Z(n16974) );
  NANDN U17581 ( .A(n17475), .B(\stack[3][13] ), .Z(n16973) );
  NAND U17582 ( .A(n16974), .B(n16973), .Z(n2531) );
  NANDN U17583 ( .A(n2974), .B(n17471), .Z(n16976) );
  NANDN U17584 ( .A(n17472), .B(\stack[3][13] ), .Z(n16975) );
  AND U17585 ( .A(n16976), .B(n16975), .Z(n16978) );
  NANDN U17586 ( .A(n17475), .B(\stack[2][13] ), .Z(n16977) );
  NAND U17587 ( .A(n16978), .B(n16977), .Z(n2532) );
  NANDN U17588 ( .A(n3007), .B(n17471), .Z(n16980) );
  NANDN U17589 ( .A(n17472), .B(\stack[2][13] ), .Z(n16979) );
  AND U17590 ( .A(n16980), .B(n16979), .Z(n16982) );
  OR U17591 ( .A(n17475), .B(n2974), .Z(n16981) );
  NAND U17592 ( .A(n16982), .B(n16981), .Z(n2533) );
  NANDN U17593 ( .A(n2974), .B(n17461), .Z(n16985) );
  NAND U17594 ( .A(n16983), .B(n17479), .Z(n16984) );
  NAND U17595 ( .A(n16985), .B(n16984), .Z(n16993) );
  XNOR U17596 ( .A(n16987), .B(n16986), .Z(n16988) );
  NAND U17597 ( .A(n16988), .B(n17458), .Z(n16991) );
  NANDN U17598 ( .A(n2967), .B(x[13]), .Z(n16989) );
  NAND U17599 ( .A(n16991), .B(n16990), .Z(n16992) );
  NOR U17600 ( .A(n16993), .B(n16992), .Z(n16995) );
  NANDN U17601 ( .A(n3007), .B(n17467), .Z(n16994) );
  NAND U17602 ( .A(n16995), .B(n16994), .Z(n2534) );
  NANDN U17603 ( .A(n2967), .B(\stack[6][12] ), .Z(n16997) );
  NANDN U17604 ( .A(n17471), .B(\stack[7][12] ), .Z(n16996) );
  NAND U17605 ( .A(n16997), .B(n16996), .Z(n2535) );
  NANDN U17606 ( .A(n2967), .B(\stack[5][12] ), .Z(n16999) );
  NANDN U17607 ( .A(n17472), .B(\stack[7][12] ), .Z(n16998) );
  AND U17608 ( .A(n16999), .B(n16998), .Z(n17001) );
  NANDN U17609 ( .A(n17475), .B(\stack[6][12] ), .Z(n17000) );
  NAND U17610 ( .A(n17001), .B(n17000), .Z(n2536) );
  NANDN U17611 ( .A(n2967), .B(\stack[4][12] ), .Z(n17003) );
  NANDN U17612 ( .A(n17472), .B(\stack[6][12] ), .Z(n17002) );
  AND U17613 ( .A(n17003), .B(n17002), .Z(n17005) );
  NANDN U17614 ( .A(n17475), .B(\stack[5][12] ), .Z(n17004) );
  NAND U17615 ( .A(n17005), .B(n17004), .Z(n2537) );
  NANDN U17616 ( .A(n2967), .B(\stack[3][12] ), .Z(n17007) );
  NANDN U17617 ( .A(n17472), .B(\stack[5][12] ), .Z(n17006) );
  AND U17618 ( .A(n17007), .B(n17006), .Z(n17009) );
  NANDN U17619 ( .A(n17475), .B(\stack[4][12] ), .Z(n17008) );
  NAND U17620 ( .A(n17009), .B(n17008), .Z(n2538) );
  NANDN U17621 ( .A(n2967), .B(\stack[2][12] ), .Z(n17011) );
  NANDN U17622 ( .A(n17472), .B(\stack[4][12] ), .Z(n17010) );
  AND U17623 ( .A(n17011), .B(n17010), .Z(n17013) );
  NANDN U17624 ( .A(n17475), .B(\stack[3][12] ), .Z(n17012) );
  NAND U17625 ( .A(n17013), .B(n17012), .Z(n2539) );
  NANDN U17626 ( .A(n2973), .B(n17471), .Z(n17015) );
  NANDN U17627 ( .A(n17472), .B(\stack[3][12] ), .Z(n17014) );
  AND U17628 ( .A(n17015), .B(n17014), .Z(n17017) );
  NANDN U17629 ( .A(n17475), .B(\stack[2][12] ), .Z(n17016) );
  NAND U17630 ( .A(n17017), .B(n17016), .Z(n2540) );
  NANDN U17631 ( .A(n3006), .B(n17471), .Z(n17019) );
  NANDN U17632 ( .A(n17472), .B(\stack[2][12] ), .Z(n17018) );
  AND U17633 ( .A(n17019), .B(n17018), .Z(n17021) );
  OR U17634 ( .A(n17475), .B(n2973), .Z(n17020) );
  NAND U17635 ( .A(n17021), .B(n17020), .Z(n2541) );
  NANDN U17636 ( .A(n2967), .B(x[12]), .Z(n17023) );
  NANDN U17637 ( .A(n17483), .B(\stack[1][12] ), .Z(n17022) );
  NAND U17638 ( .A(n17023), .B(n17022), .Z(n17032) );
  XNOR U17639 ( .A(n17025), .B(n17024), .Z(n17026) );
  NAND U17640 ( .A(n17026), .B(n17458), .Z(n17030) );
  NAND U17641 ( .A(n17027), .B(n17479), .Z(n17028) );
  NAND U17642 ( .A(n17030), .B(n17029), .Z(n17031) );
  NOR U17643 ( .A(n17032), .B(n17031), .Z(n17034) );
  NANDN U17644 ( .A(n3006), .B(n17467), .Z(n17033) );
  NAND U17645 ( .A(n17034), .B(n17033), .Z(n2542) );
  NANDN U17646 ( .A(n2967), .B(\stack[6][11] ), .Z(n17036) );
  NANDN U17647 ( .A(n17471), .B(\stack[7][11] ), .Z(n17035) );
  NAND U17648 ( .A(n17036), .B(n17035), .Z(n2543) );
  NANDN U17649 ( .A(n2967), .B(\stack[5][11] ), .Z(n17038) );
  NANDN U17650 ( .A(n17472), .B(\stack[7][11] ), .Z(n17037) );
  AND U17651 ( .A(n17038), .B(n17037), .Z(n17040) );
  NANDN U17652 ( .A(n17475), .B(\stack[6][11] ), .Z(n17039) );
  NAND U17653 ( .A(n17040), .B(n17039), .Z(n2544) );
  NANDN U17654 ( .A(n2967), .B(\stack[4][11] ), .Z(n17042) );
  NANDN U17655 ( .A(n17472), .B(\stack[6][11] ), .Z(n17041) );
  AND U17656 ( .A(n17042), .B(n17041), .Z(n17044) );
  NANDN U17657 ( .A(n17475), .B(\stack[5][11] ), .Z(n17043) );
  NAND U17658 ( .A(n17044), .B(n17043), .Z(n2545) );
  NANDN U17659 ( .A(n2967), .B(\stack[3][11] ), .Z(n17046) );
  NANDN U17660 ( .A(n17472), .B(\stack[5][11] ), .Z(n17045) );
  AND U17661 ( .A(n17046), .B(n17045), .Z(n17048) );
  NANDN U17662 ( .A(n17475), .B(\stack[4][11] ), .Z(n17047) );
  NAND U17663 ( .A(n17048), .B(n17047), .Z(n2546) );
  NANDN U17664 ( .A(n2967), .B(\stack[2][11] ), .Z(n17050) );
  NANDN U17665 ( .A(n17472), .B(\stack[4][11] ), .Z(n17049) );
  AND U17666 ( .A(n17050), .B(n17049), .Z(n17052) );
  NANDN U17667 ( .A(n17475), .B(\stack[3][11] ), .Z(n17051) );
  NAND U17668 ( .A(n17052), .B(n17051), .Z(n2547) );
  NANDN U17669 ( .A(n2972), .B(n17471), .Z(n17054) );
  NANDN U17670 ( .A(n17472), .B(\stack[3][11] ), .Z(n17053) );
  AND U17671 ( .A(n17054), .B(n17053), .Z(n17056) );
  NANDN U17672 ( .A(n17475), .B(\stack[2][11] ), .Z(n17055) );
  NAND U17673 ( .A(n17056), .B(n17055), .Z(n2548) );
  NANDN U17674 ( .A(n3005), .B(n17471), .Z(n17058) );
  NANDN U17675 ( .A(n17472), .B(\stack[2][11] ), .Z(n17057) );
  AND U17676 ( .A(n17058), .B(n17057), .Z(n17060) );
  OR U17677 ( .A(n17475), .B(n2972), .Z(n17059) );
  NAND U17678 ( .A(n17060), .B(n17059), .Z(n2549) );
  NANDN U17679 ( .A(n2967), .B(x[11]), .Z(n17063) );
  NAND U17680 ( .A(n17061), .B(n17479), .Z(n17062) );
  NAND U17681 ( .A(n17063), .B(n17062), .Z(n17071) );
  XNOR U17682 ( .A(n17065), .B(n17064), .Z(n17066) );
  NAND U17683 ( .A(n17066), .B(n17458), .Z(n17069) );
  NANDN U17684 ( .A(n2972), .B(n17461), .Z(n17067) );
  NAND U17685 ( .A(n17069), .B(n17068), .Z(n17070) );
  NOR U17686 ( .A(n17071), .B(n17070), .Z(n17073) );
  NANDN U17687 ( .A(n3005), .B(n17467), .Z(n17072) );
  NAND U17688 ( .A(n17073), .B(n17072), .Z(n2550) );
  NANDN U17689 ( .A(n2967), .B(\stack[6][10] ), .Z(n17075) );
  NANDN U17690 ( .A(n17471), .B(\stack[7][10] ), .Z(n17074) );
  NAND U17691 ( .A(n17075), .B(n17074), .Z(n2551) );
  NANDN U17692 ( .A(n2967), .B(\stack[5][10] ), .Z(n17077) );
  NANDN U17693 ( .A(n17472), .B(\stack[7][10] ), .Z(n17076) );
  AND U17694 ( .A(n17077), .B(n17076), .Z(n17079) );
  NANDN U17695 ( .A(n17475), .B(\stack[6][10] ), .Z(n17078) );
  NAND U17696 ( .A(n17079), .B(n17078), .Z(n2552) );
  NANDN U17697 ( .A(n2967), .B(\stack[4][10] ), .Z(n17081) );
  NANDN U17698 ( .A(n17472), .B(\stack[6][10] ), .Z(n17080) );
  AND U17699 ( .A(n17081), .B(n17080), .Z(n17083) );
  NANDN U17700 ( .A(n17475), .B(\stack[5][10] ), .Z(n17082) );
  NAND U17701 ( .A(n17083), .B(n17082), .Z(n2553) );
  NANDN U17702 ( .A(n2967), .B(\stack[3][10] ), .Z(n17085) );
  NANDN U17703 ( .A(n17472), .B(\stack[5][10] ), .Z(n17084) );
  AND U17704 ( .A(n17085), .B(n17084), .Z(n17087) );
  NANDN U17705 ( .A(n17475), .B(\stack[4][10] ), .Z(n17086) );
  NAND U17706 ( .A(n17087), .B(n17086), .Z(n2554) );
  NANDN U17707 ( .A(n2967), .B(\stack[2][10] ), .Z(n17089) );
  NANDN U17708 ( .A(n17472), .B(\stack[4][10] ), .Z(n17088) );
  AND U17709 ( .A(n17089), .B(n17088), .Z(n17091) );
  NANDN U17710 ( .A(n17475), .B(\stack[3][10] ), .Z(n17090) );
  NAND U17711 ( .A(n17091), .B(n17090), .Z(n2555) );
  NANDN U17712 ( .A(n17101), .B(n17471), .Z(n17093) );
  NANDN U17713 ( .A(n17472), .B(\stack[3][10] ), .Z(n17092) );
  AND U17714 ( .A(n17093), .B(n17092), .Z(n17095) );
  NANDN U17715 ( .A(n17475), .B(\stack[2][10] ), .Z(n17094) );
  NAND U17716 ( .A(n17095), .B(n17094), .Z(n2556) );
  NANDN U17717 ( .A(n3004), .B(n17471), .Z(n17097) );
  NANDN U17718 ( .A(n17472), .B(\stack[2][10] ), .Z(n17096) );
  AND U17719 ( .A(n17097), .B(n17096), .Z(n17099) );
  OR U17720 ( .A(n17475), .B(n17101), .Z(n17098) );
  NAND U17721 ( .A(n17099), .B(n17098), .Z(n2557) );
  NANDN U17722 ( .A(n3004), .B(n17479), .Z(n17100) );
  NANDN U17723 ( .A(n17461), .B(n17100), .Z(n17102) );
  ANDN U17724 ( .B(n17102), .A(n17101), .Z(n17110) );
  XNOR U17725 ( .A(n17104), .B(n17103), .Z(n17105) );
  NAND U17726 ( .A(n17105), .B(n17458), .Z(n17108) );
  NANDN U17727 ( .A(n2967), .B(x[10]), .Z(n17106) );
  NAND U17728 ( .A(n17108), .B(n17107), .Z(n17109) );
  NOR U17729 ( .A(n17110), .B(n17109), .Z(n17112) );
  NANDN U17730 ( .A(n3004), .B(n17467), .Z(n17111) );
  NAND U17731 ( .A(n17112), .B(n17111), .Z(n2558) );
  NANDN U17732 ( .A(n2967), .B(\stack[6][9] ), .Z(n17114) );
  NANDN U17733 ( .A(n17471), .B(\stack[7][9] ), .Z(n17113) );
  NAND U17734 ( .A(n17114), .B(n17113), .Z(n2559) );
  NANDN U17735 ( .A(n2967), .B(\stack[5][9] ), .Z(n17116) );
  NANDN U17736 ( .A(n17472), .B(\stack[7][9] ), .Z(n17115) );
  AND U17737 ( .A(n17116), .B(n17115), .Z(n17118) );
  NANDN U17738 ( .A(n17475), .B(\stack[6][9] ), .Z(n17117) );
  NAND U17739 ( .A(n17118), .B(n17117), .Z(n2560) );
  NANDN U17740 ( .A(n2967), .B(\stack[4][9] ), .Z(n17120) );
  NANDN U17741 ( .A(n17472), .B(\stack[6][9] ), .Z(n17119) );
  AND U17742 ( .A(n17120), .B(n17119), .Z(n17122) );
  NANDN U17743 ( .A(n17475), .B(\stack[5][9] ), .Z(n17121) );
  NAND U17744 ( .A(n17122), .B(n17121), .Z(n2561) );
  NANDN U17745 ( .A(n2967), .B(\stack[3][9] ), .Z(n17124) );
  NANDN U17746 ( .A(n17472), .B(\stack[5][9] ), .Z(n17123) );
  AND U17747 ( .A(n17124), .B(n17123), .Z(n17126) );
  NANDN U17748 ( .A(n17475), .B(\stack[4][9] ), .Z(n17125) );
  NAND U17749 ( .A(n17126), .B(n17125), .Z(n2562) );
  NANDN U17750 ( .A(n2967), .B(\stack[2][9] ), .Z(n17128) );
  NANDN U17751 ( .A(n17472), .B(\stack[4][9] ), .Z(n17127) );
  AND U17752 ( .A(n17128), .B(n17127), .Z(n17130) );
  NANDN U17753 ( .A(n17475), .B(\stack[3][9] ), .Z(n17129) );
  NAND U17754 ( .A(n17130), .B(n17129), .Z(n2563) );
  NANDN U17755 ( .A(n17145), .B(n17471), .Z(n17132) );
  NANDN U17756 ( .A(n17472), .B(\stack[3][9] ), .Z(n17131) );
  AND U17757 ( .A(n17132), .B(n17131), .Z(n17134) );
  NANDN U17758 ( .A(n17475), .B(\stack[2][9] ), .Z(n17133) );
  NAND U17759 ( .A(n17134), .B(n17133), .Z(n2564) );
  NANDN U17760 ( .A(n3003), .B(n17471), .Z(n17136) );
  NANDN U17761 ( .A(n17472), .B(\stack[2][9] ), .Z(n17135) );
  AND U17762 ( .A(n17136), .B(n17135), .Z(n17138) );
  OR U17763 ( .A(n17475), .B(n17145), .Z(n17137) );
  NAND U17764 ( .A(n17138), .B(n17137), .Z(n2565) );
  NAND U17765 ( .A(n17479), .B(n17139), .Z(n17141) );
  NANDN U17766 ( .A(n2967), .B(x[9]), .Z(n17140) );
  NAND U17767 ( .A(n17141), .B(n17140), .Z(n17150) );
  XNOR U17768 ( .A(n17143), .B(n17142), .Z(n17144) );
  NAND U17769 ( .A(n17144), .B(n17458), .Z(n17148) );
  NANDN U17770 ( .A(n17145), .B(n17461), .Z(n17146) );
  NAND U17771 ( .A(n17148), .B(n17147), .Z(n17149) );
  NOR U17772 ( .A(n17150), .B(n17149), .Z(n17152) );
  NANDN U17773 ( .A(n3003), .B(n17467), .Z(n17151) );
  NAND U17774 ( .A(n17152), .B(n17151), .Z(n2566) );
  NANDN U17775 ( .A(n2967), .B(\stack[6][8] ), .Z(n17154) );
  NANDN U17776 ( .A(n17471), .B(\stack[7][8] ), .Z(n17153) );
  NAND U17777 ( .A(n17154), .B(n17153), .Z(n2567) );
  NANDN U17778 ( .A(n2967), .B(\stack[5][8] ), .Z(n17156) );
  NANDN U17779 ( .A(n17472), .B(\stack[7][8] ), .Z(n17155) );
  AND U17780 ( .A(n17156), .B(n17155), .Z(n17158) );
  NANDN U17781 ( .A(n17475), .B(\stack[6][8] ), .Z(n17157) );
  NAND U17782 ( .A(n17158), .B(n17157), .Z(n2568) );
  NANDN U17783 ( .A(n2967), .B(\stack[4][8] ), .Z(n17160) );
  NANDN U17784 ( .A(n17472), .B(\stack[6][8] ), .Z(n17159) );
  AND U17785 ( .A(n17160), .B(n17159), .Z(n17162) );
  NANDN U17786 ( .A(n17475), .B(\stack[5][8] ), .Z(n17161) );
  NAND U17787 ( .A(n17162), .B(n17161), .Z(n2569) );
  NANDN U17788 ( .A(n2967), .B(\stack[3][8] ), .Z(n17164) );
  NANDN U17789 ( .A(n17472), .B(\stack[5][8] ), .Z(n17163) );
  AND U17790 ( .A(n17164), .B(n17163), .Z(n17166) );
  NANDN U17791 ( .A(n17475), .B(\stack[4][8] ), .Z(n17165) );
  NAND U17792 ( .A(n17166), .B(n17165), .Z(n2570) );
  NANDN U17793 ( .A(n2967), .B(\stack[2][8] ), .Z(n17168) );
  NANDN U17794 ( .A(n17472), .B(\stack[4][8] ), .Z(n17167) );
  AND U17795 ( .A(n17168), .B(n17167), .Z(n17170) );
  NANDN U17796 ( .A(n17475), .B(\stack[3][8] ), .Z(n17169) );
  NAND U17797 ( .A(n17170), .B(n17169), .Z(n2571) );
  NANDN U17798 ( .A(n17179), .B(n17471), .Z(n17172) );
  NANDN U17799 ( .A(n17472), .B(\stack[3][8] ), .Z(n17171) );
  AND U17800 ( .A(n17172), .B(n17171), .Z(n17174) );
  NANDN U17801 ( .A(n17475), .B(\stack[2][8] ), .Z(n17173) );
  NAND U17802 ( .A(n17174), .B(n17173), .Z(n2572) );
  NANDN U17803 ( .A(n3002), .B(n17471), .Z(n17176) );
  NANDN U17804 ( .A(n17472), .B(\stack[2][8] ), .Z(n17175) );
  AND U17805 ( .A(n17176), .B(n17175), .Z(n17178) );
  OR U17806 ( .A(n17475), .B(n17179), .Z(n17177) );
  NAND U17807 ( .A(n17178), .B(n17177), .Z(n2573) );
  NANDN U17808 ( .A(n17179), .B(n17461), .Z(n17182) );
  NAND U17809 ( .A(n17180), .B(n17479), .Z(n17181) );
  NAND U17810 ( .A(n17182), .B(n17181), .Z(n17190) );
  XNOR U17811 ( .A(n17184), .B(n17183), .Z(n17185) );
  NAND U17812 ( .A(n17185), .B(n17458), .Z(n17188) );
  NANDN U17813 ( .A(n2967), .B(x[8]), .Z(n17186) );
  NAND U17814 ( .A(n17188), .B(n17187), .Z(n17189) );
  NOR U17815 ( .A(n17190), .B(n17189), .Z(n17192) );
  NANDN U17816 ( .A(n3002), .B(n17467), .Z(n17191) );
  NAND U17817 ( .A(n17192), .B(n17191), .Z(n2574) );
  NANDN U17818 ( .A(n2967), .B(\stack[6][7] ), .Z(n17194) );
  NANDN U17819 ( .A(n17471), .B(\stack[7][7] ), .Z(n17193) );
  NAND U17820 ( .A(n17194), .B(n17193), .Z(n2575) );
  NANDN U17821 ( .A(n2967), .B(\stack[5][7] ), .Z(n17196) );
  NANDN U17822 ( .A(n17472), .B(\stack[7][7] ), .Z(n17195) );
  AND U17823 ( .A(n17196), .B(n17195), .Z(n17198) );
  NANDN U17824 ( .A(n17475), .B(\stack[6][7] ), .Z(n17197) );
  NAND U17825 ( .A(n17198), .B(n17197), .Z(n2576) );
  NANDN U17826 ( .A(n2967), .B(\stack[4][7] ), .Z(n17200) );
  NANDN U17827 ( .A(n17472), .B(\stack[6][7] ), .Z(n17199) );
  AND U17828 ( .A(n17200), .B(n17199), .Z(n17202) );
  NANDN U17829 ( .A(n17475), .B(\stack[5][7] ), .Z(n17201) );
  NAND U17830 ( .A(n17202), .B(n17201), .Z(n2577) );
  NANDN U17831 ( .A(n2967), .B(\stack[3][7] ), .Z(n17204) );
  NANDN U17832 ( .A(n17472), .B(\stack[5][7] ), .Z(n17203) );
  AND U17833 ( .A(n17204), .B(n17203), .Z(n17206) );
  NANDN U17834 ( .A(n17475), .B(\stack[4][7] ), .Z(n17205) );
  NAND U17835 ( .A(n17206), .B(n17205), .Z(n2578) );
  NANDN U17836 ( .A(n2967), .B(\stack[2][7] ), .Z(n17208) );
  NANDN U17837 ( .A(n17472), .B(\stack[4][7] ), .Z(n17207) );
  AND U17838 ( .A(n17208), .B(n17207), .Z(n17210) );
  NANDN U17839 ( .A(n17475), .B(\stack[3][7] ), .Z(n17209) );
  NAND U17840 ( .A(n17210), .B(n17209), .Z(n2579) );
  NANDN U17841 ( .A(n17219), .B(n17471), .Z(n17212) );
  NANDN U17842 ( .A(n17472), .B(\stack[3][7] ), .Z(n17211) );
  AND U17843 ( .A(n17212), .B(n17211), .Z(n17214) );
  NANDN U17844 ( .A(n17475), .B(\stack[2][7] ), .Z(n17213) );
  NAND U17845 ( .A(n17214), .B(n17213), .Z(n2580) );
  NANDN U17846 ( .A(n3001), .B(n17471), .Z(n17216) );
  NANDN U17847 ( .A(n17472), .B(\stack[2][7] ), .Z(n17215) );
  AND U17848 ( .A(n17216), .B(n17215), .Z(n17218) );
  OR U17849 ( .A(n17475), .B(n17219), .Z(n17217) );
  NAND U17850 ( .A(n17218), .B(n17217), .Z(n2581) );
  NANDN U17851 ( .A(n17219), .B(n17479), .Z(n17220) );
  NANDN U17852 ( .A(n17467), .B(n17220), .Z(n17221) );
  ANDN U17853 ( .B(n17221), .A(n3001), .Z(n17230) );
  XNOR U17854 ( .A(n17223), .B(n17222), .Z(n17224) );
  NAND U17855 ( .A(n17224), .B(n17458), .Z(n17228) );
  NANDN U17856 ( .A(n2967), .B(x[7]), .Z(n17226) );
  NANDN U17857 ( .A(n17483), .B(\stack[1][7] ), .Z(n17225) );
  AND U17858 ( .A(n17226), .B(n17225), .Z(n17227) );
  NAND U17859 ( .A(n17228), .B(n17227), .Z(n17229) );
  NOR U17860 ( .A(n17230), .B(n17229), .Z(n17231) );
  NANDN U17861 ( .A(n2967), .B(\stack[6][6] ), .Z(n17233) );
  NANDN U17862 ( .A(n17471), .B(\stack[7][6] ), .Z(n17232) );
  NAND U17863 ( .A(n17233), .B(n17232), .Z(n2583) );
  NANDN U17864 ( .A(n2967), .B(\stack[5][6] ), .Z(n17235) );
  NANDN U17865 ( .A(n17472), .B(\stack[7][6] ), .Z(n17234) );
  AND U17866 ( .A(n17235), .B(n17234), .Z(n17237) );
  NANDN U17867 ( .A(n17475), .B(\stack[6][6] ), .Z(n17236) );
  NAND U17868 ( .A(n17237), .B(n17236), .Z(n2584) );
  NANDN U17869 ( .A(n2967), .B(\stack[4][6] ), .Z(n17239) );
  NANDN U17870 ( .A(n17472), .B(\stack[6][6] ), .Z(n17238) );
  AND U17871 ( .A(n17239), .B(n17238), .Z(n17241) );
  NANDN U17872 ( .A(n17475), .B(\stack[5][6] ), .Z(n17240) );
  NAND U17873 ( .A(n17241), .B(n17240), .Z(n2585) );
  NANDN U17874 ( .A(n2967), .B(\stack[3][6] ), .Z(n17243) );
  NANDN U17875 ( .A(n17472), .B(\stack[5][6] ), .Z(n17242) );
  AND U17876 ( .A(n17243), .B(n17242), .Z(n17245) );
  NANDN U17877 ( .A(n17475), .B(\stack[4][6] ), .Z(n17244) );
  NAND U17878 ( .A(n17245), .B(n17244), .Z(n2586) );
  NANDN U17879 ( .A(n2967), .B(\stack[2][6] ), .Z(n17247) );
  NANDN U17880 ( .A(n17472), .B(\stack[4][6] ), .Z(n17246) );
  AND U17881 ( .A(n17247), .B(n17246), .Z(n17249) );
  NANDN U17882 ( .A(n17475), .B(\stack[3][6] ), .Z(n17248) );
  NAND U17883 ( .A(n17249), .B(n17248), .Z(n2587) );
  NANDN U17884 ( .A(n17256), .B(n17471), .Z(n17251) );
  NANDN U17885 ( .A(n17472), .B(\stack[3][6] ), .Z(n17250) );
  AND U17886 ( .A(n17251), .B(n17250), .Z(n17253) );
  NANDN U17887 ( .A(n17475), .B(\stack[2][6] ), .Z(n17252) );
  NAND U17888 ( .A(n17253), .B(n17252), .Z(n2588) );
  NANDN U17889 ( .A(n3000), .B(n17471), .Z(n17255) );
  NANDN U17890 ( .A(n17472), .B(\stack[2][6] ), .Z(n17254) );
  AND U17891 ( .A(n17255), .B(n17254), .Z(n17258) );
  OR U17892 ( .A(n17475), .B(n17256), .Z(n17257) );
  NAND U17893 ( .A(n17258), .B(n17257), .Z(n2589) );
  NANDN U17894 ( .A(n2967), .B(x[6]), .Z(n17259) );
  XNOR U17895 ( .A(n17261), .B(n17260), .Z(n17262) );
  NAND U17896 ( .A(n17262), .B(n17458), .Z(n17263) );
  AND U17897 ( .A(n17264), .B(n17263), .Z(n17269) );
  NAND U17898 ( .A(n17265), .B(n17479), .Z(n17267) );
  NANDN U17899 ( .A(n17483), .B(\stack[1][6] ), .Z(n17266) );
  AND U17900 ( .A(n17267), .B(n17266), .Z(n17268) );
  AND U17901 ( .A(n17269), .B(n17268), .Z(n17271) );
  NANDN U17902 ( .A(n3000), .B(n17467), .Z(n17270) );
  NAND U17903 ( .A(n17271), .B(n17270), .Z(n2590) );
  NANDN U17904 ( .A(n2967), .B(\stack[6][5] ), .Z(n17273) );
  NANDN U17905 ( .A(n17471), .B(\stack[7][5] ), .Z(n17272) );
  NAND U17906 ( .A(n17273), .B(n17272), .Z(n2591) );
  NANDN U17907 ( .A(n2967), .B(\stack[5][5] ), .Z(n17275) );
  NANDN U17908 ( .A(n17472), .B(\stack[7][5] ), .Z(n17274) );
  AND U17909 ( .A(n17275), .B(n17274), .Z(n17277) );
  NANDN U17910 ( .A(n17475), .B(\stack[6][5] ), .Z(n17276) );
  NAND U17911 ( .A(n17277), .B(n17276), .Z(n2592) );
  NANDN U17912 ( .A(n2967), .B(\stack[4][5] ), .Z(n17279) );
  NANDN U17913 ( .A(n17472), .B(\stack[6][5] ), .Z(n17278) );
  AND U17914 ( .A(n17279), .B(n17278), .Z(n17281) );
  NANDN U17915 ( .A(n17475), .B(\stack[5][5] ), .Z(n17280) );
  NAND U17916 ( .A(n17281), .B(n17280), .Z(n2593) );
  NANDN U17917 ( .A(n2967), .B(\stack[3][5] ), .Z(n17283) );
  NANDN U17918 ( .A(n17472), .B(\stack[5][5] ), .Z(n17282) );
  AND U17919 ( .A(n17283), .B(n17282), .Z(n17285) );
  NANDN U17920 ( .A(n17475), .B(\stack[4][5] ), .Z(n17284) );
  NAND U17921 ( .A(n17285), .B(n17284), .Z(n2594) );
  NANDN U17922 ( .A(n2967), .B(\stack[2][5] ), .Z(n17287) );
  NANDN U17923 ( .A(n17472), .B(\stack[4][5] ), .Z(n17286) );
  AND U17924 ( .A(n17287), .B(n17286), .Z(n17289) );
  NANDN U17925 ( .A(n17475), .B(\stack[3][5] ), .Z(n17288) );
  NAND U17926 ( .A(n17289), .B(n17288), .Z(n2595) );
  NANDN U17927 ( .A(n17296), .B(n17471), .Z(n17291) );
  NANDN U17928 ( .A(n17472), .B(\stack[3][5] ), .Z(n17290) );
  AND U17929 ( .A(n17291), .B(n17290), .Z(n17293) );
  NANDN U17930 ( .A(n17475), .B(\stack[2][5] ), .Z(n17292) );
  NAND U17931 ( .A(n17293), .B(n17292), .Z(n2596) );
  NANDN U17932 ( .A(n2999), .B(n17471), .Z(n17295) );
  NANDN U17933 ( .A(n17472), .B(\stack[2][5] ), .Z(n17294) );
  AND U17934 ( .A(n17295), .B(n17294), .Z(n17298) );
  OR U17935 ( .A(n17475), .B(n17296), .Z(n17297) );
  NAND U17936 ( .A(n17298), .B(n17297), .Z(n2597) );
  XNOR U17937 ( .A(n17300), .B(n17299), .Z(n17301) );
  NAND U17938 ( .A(n17301), .B(n17458), .Z(n17305) );
  NAND U17939 ( .A(n17302), .B(n17479), .Z(n17303) );
  ANDN U17940 ( .B(n17305), .A(n17304), .Z(n17309) );
  NANDN U17941 ( .A(n2967), .B(x[5]), .Z(n17307) );
  NANDN U17942 ( .A(n17483), .B(\stack[1][5] ), .Z(n17306) );
  NAND U17943 ( .A(n17307), .B(n17306), .Z(n17308) );
  ANDN U17944 ( .B(n17309), .A(n17308), .Z(n17311) );
  NANDN U17945 ( .A(n2999), .B(n17467), .Z(n17310) );
  NAND U17946 ( .A(n17311), .B(n17310), .Z(n2598) );
  NANDN U17947 ( .A(n2967), .B(\stack[6][4] ), .Z(n17313) );
  NANDN U17948 ( .A(n17471), .B(\stack[7][4] ), .Z(n17312) );
  NAND U17949 ( .A(n17313), .B(n17312), .Z(n2599) );
  NANDN U17950 ( .A(n2967), .B(\stack[5][4] ), .Z(n17315) );
  NANDN U17951 ( .A(n17472), .B(\stack[7][4] ), .Z(n17314) );
  AND U17952 ( .A(n17315), .B(n17314), .Z(n17317) );
  NANDN U17953 ( .A(n17475), .B(\stack[6][4] ), .Z(n17316) );
  NAND U17954 ( .A(n17317), .B(n17316), .Z(n2600) );
  NANDN U17955 ( .A(n2967), .B(\stack[4][4] ), .Z(n17319) );
  NANDN U17956 ( .A(n17472), .B(\stack[6][4] ), .Z(n17318) );
  AND U17957 ( .A(n17319), .B(n17318), .Z(n17321) );
  NANDN U17958 ( .A(n17475), .B(\stack[5][4] ), .Z(n17320) );
  NAND U17959 ( .A(n17321), .B(n17320), .Z(n2601) );
  NANDN U17960 ( .A(n2967), .B(\stack[3][4] ), .Z(n17323) );
  NANDN U17961 ( .A(n17472), .B(\stack[5][4] ), .Z(n17322) );
  AND U17962 ( .A(n17323), .B(n17322), .Z(n17325) );
  NANDN U17963 ( .A(n17475), .B(\stack[4][4] ), .Z(n17324) );
  NAND U17964 ( .A(n17325), .B(n17324), .Z(n2602) );
  NANDN U17965 ( .A(n2967), .B(\stack[2][4] ), .Z(n17327) );
  NANDN U17966 ( .A(n17472), .B(\stack[4][4] ), .Z(n17326) );
  AND U17967 ( .A(n17327), .B(n17326), .Z(n17329) );
  NANDN U17968 ( .A(n17475), .B(\stack[3][4] ), .Z(n17328) );
  NAND U17969 ( .A(n17329), .B(n17328), .Z(n2603) );
  NANDN U17970 ( .A(n2971), .B(n17471), .Z(n17331) );
  NANDN U17971 ( .A(n17472), .B(\stack[3][4] ), .Z(n17330) );
  AND U17972 ( .A(n17331), .B(n17330), .Z(n17333) );
  NANDN U17973 ( .A(n17475), .B(\stack[2][4] ), .Z(n17332) );
  NAND U17974 ( .A(n17333), .B(n17332), .Z(n2604) );
  NANDN U17975 ( .A(n2998), .B(n17471), .Z(n17335) );
  NANDN U17976 ( .A(n17472), .B(\stack[2][4] ), .Z(n17334) );
  AND U17977 ( .A(n17335), .B(n17334), .Z(n17337) );
  OR U17978 ( .A(n17475), .B(n2971), .Z(n17336) );
  NAND U17979 ( .A(n17337), .B(n17336), .Z(n2605) );
  NANDN U17980 ( .A(n2971), .B(n17461), .Z(n17340) );
  NAND U17981 ( .A(n17338), .B(n17479), .Z(n17339) );
  NAND U17982 ( .A(n17340), .B(n17339), .Z(n17348) );
  XNOR U17983 ( .A(n17342), .B(n17341), .Z(n17343) );
  NAND U17984 ( .A(n17343), .B(n17458), .Z(n17346) );
  NANDN U17985 ( .A(n2967), .B(x[4]), .Z(n17344) );
  NAND U17986 ( .A(n17346), .B(n17345), .Z(n17347) );
  NOR U17987 ( .A(n17348), .B(n17347), .Z(n17350) );
  NANDN U17988 ( .A(n2998), .B(n17467), .Z(n17349) );
  NAND U17989 ( .A(n17350), .B(n17349), .Z(n2606) );
  NANDN U17990 ( .A(n2967), .B(\stack[6][3] ), .Z(n17352) );
  NANDN U17991 ( .A(n17471), .B(\stack[7][3] ), .Z(n17351) );
  NAND U17992 ( .A(n17352), .B(n17351), .Z(n2607) );
  NANDN U17993 ( .A(n2967), .B(\stack[5][3] ), .Z(n17354) );
  NANDN U17994 ( .A(n17472), .B(\stack[7][3] ), .Z(n17353) );
  AND U17995 ( .A(n17354), .B(n17353), .Z(n17356) );
  NANDN U17996 ( .A(n17475), .B(\stack[6][3] ), .Z(n17355) );
  NAND U17997 ( .A(n17356), .B(n17355), .Z(n2608) );
  NANDN U17998 ( .A(n2967), .B(\stack[4][3] ), .Z(n17358) );
  NANDN U17999 ( .A(n17472), .B(\stack[6][3] ), .Z(n17357) );
  AND U18000 ( .A(n17358), .B(n17357), .Z(n17360) );
  NANDN U18001 ( .A(n17475), .B(\stack[5][3] ), .Z(n17359) );
  NAND U18002 ( .A(n17360), .B(n17359), .Z(n2609) );
  NANDN U18003 ( .A(n2967), .B(\stack[3][3] ), .Z(n17362) );
  NANDN U18004 ( .A(n17472), .B(\stack[5][3] ), .Z(n17361) );
  AND U18005 ( .A(n17362), .B(n17361), .Z(n17364) );
  NANDN U18006 ( .A(n17475), .B(\stack[4][3] ), .Z(n17363) );
  NAND U18007 ( .A(n17364), .B(n17363), .Z(n2610) );
  NANDN U18008 ( .A(n2967), .B(\stack[2][3] ), .Z(n17366) );
  NANDN U18009 ( .A(n17472), .B(\stack[4][3] ), .Z(n17365) );
  AND U18010 ( .A(n17366), .B(n17365), .Z(n17368) );
  NANDN U18011 ( .A(n17475), .B(\stack[3][3] ), .Z(n17367) );
  NAND U18012 ( .A(n17368), .B(n17367), .Z(n2611) );
  NANDN U18013 ( .A(n17375), .B(n17471), .Z(n17370) );
  NANDN U18014 ( .A(n17472), .B(\stack[3][3] ), .Z(n17369) );
  AND U18015 ( .A(n17370), .B(n17369), .Z(n17372) );
  NANDN U18016 ( .A(n17475), .B(\stack[2][3] ), .Z(n17371) );
  NAND U18017 ( .A(n17372), .B(n17371), .Z(n2612) );
  NANDN U18018 ( .A(n2997), .B(n17471), .Z(n17374) );
  NANDN U18019 ( .A(n17472), .B(\stack[2][3] ), .Z(n17373) );
  AND U18020 ( .A(n17374), .B(n17373), .Z(n17377) );
  OR U18021 ( .A(n17475), .B(n17375), .Z(n17376) );
  NAND U18022 ( .A(n17377), .B(n17376), .Z(n2613) );
  NANDN U18023 ( .A(n2967), .B(x[3]), .Z(n17378) );
  XNOR U18024 ( .A(n17380), .B(n17379), .Z(n17381) );
  NAND U18025 ( .A(n17381), .B(n17458), .Z(n17382) );
  AND U18026 ( .A(n17383), .B(n17382), .Z(n17388) );
  NAND U18027 ( .A(n17384), .B(n17479), .Z(n17386) );
  NANDN U18028 ( .A(n17483), .B(\stack[1][3] ), .Z(n17385) );
  AND U18029 ( .A(n17386), .B(n17385), .Z(n17387) );
  AND U18030 ( .A(n17388), .B(n17387), .Z(n17390) );
  NANDN U18031 ( .A(n2997), .B(n17467), .Z(n17389) );
  NAND U18032 ( .A(n17390), .B(n17389), .Z(n2614) );
  NANDN U18033 ( .A(n2967), .B(\stack[6][2] ), .Z(n17392) );
  NANDN U18034 ( .A(n17471), .B(\stack[7][2] ), .Z(n17391) );
  NAND U18035 ( .A(n17392), .B(n17391), .Z(n2615) );
  NANDN U18036 ( .A(n2967), .B(\stack[5][2] ), .Z(n17394) );
  NANDN U18037 ( .A(n17472), .B(\stack[7][2] ), .Z(n17393) );
  AND U18038 ( .A(n17394), .B(n17393), .Z(n17396) );
  NANDN U18039 ( .A(n17475), .B(\stack[6][2] ), .Z(n17395) );
  NAND U18040 ( .A(n17396), .B(n17395), .Z(n2616) );
  NANDN U18041 ( .A(n2967), .B(\stack[4][2] ), .Z(n17398) );
  NANDN U18042 ( .A(n17472), .B(\stack[6][2] ), .Z(n17397) );
  AND U18043 ( .A(n17398), .B(n17397), .Z(n17400) );
  NANDN U18044 ( .A(n17475), .B(\stack[5][2] ), .Z(n17399) );
  NAND U18045 ( .A(n17400), .B(n17399), .Z(n2617) );
  NANDN U18046 ( .A(n2967), .B(\stack[3][2] ), .Z(n17402) );
  NANDN U18047 ( .A(n17472), .B(\stack[5][2] ), .Z(n17401) );
  AND U18048 ( .A(n17402), .B(n17401), .Z(n17404) );
  NANDN U18049 ( .A(n17475), .B(\stack[4][2] ), .Z(n17403) );
  NAND U18050 ( .A(n17404), .B(n17403), .Z(n2618) );
  NANDN U18051 ( .A(n2967), .B(\stack[2][2] ), .Z(n17406) );
  NANDN U18052 ( .A(n17472), .B(\stack[4][2] ), .Z(n17405) );
  AND U18053 ( .A(n17406), .B(n17405), .Z(n17408) );
  NANDN U18054 ( .A(n17475), .B(\stack[3][2] ), .Z(n17407) );
  NAND U18055 ( .A(n17408), .B(n17407), .Z(n2619) );
  NANDN U18056 ( .A(n2970), .B(n17471), .Z(n17410) );
  NANDN U18057 ( .A(n17472), .B(\stack[3][2] ), .Z(n17409) );
  AND U18058 ( .A(n17410), .B(n17409), .Z(n17412) );
  NANDN U18059 ( .A(n17475), .B(\stack[2][2] ), .Z(n17411) );
  NAND U18060 ( .A(n17412), .B(n17411), .Z(n2620) );
  NANDN U18061 ( .A(n2996), .B(n17471), .Z(n17414) );
  NANDN U18062 ( .A(n17472), .B(\stack[2][2] ), .Z(n17413) );
  AND U18063 ( .A(n17414), .B(n17413), .Z(n17416) );
  OR U18064 ( .A(n17475), .B(n2970), .Z(n17415) );
  NAND U18065 ( .A(n17416), .B(n17415), .Z(n2621) );
  XNOR U18066 ( .A(n17418), .B(n17417), .Z(n17419) );
  NAND U18067 ( .A(n17419), .B(n17458), .Z(n17429) );
  NANDN U18068 ( .A(n17420), .B(n17479), .Z(n17421) );
  NANDN U18069 ( .A(n2967), .B(x[2]), .Z(n17423) );
  NANDN U18070 ( .A(n17483), .B(\stack[1][2] ), .Z(n17422) );
  NAND U18071 ( .A(n17423), .B(n17422), .Z(n17424) );
  NOR U18072 ( .A(n17425), .B(n17424), .Z(n17427) );
  NANDN U18073 ( .A(n2996), .B(n17467), .Z(n17426) );
  AND U18074 ( .A(n17427), .B(n17426), .Z(n17428) );
  NAND U18075 ( .A(n17429), .B(n17428), .Z(n2622) );
  NANDN U18076 ( .A(n2967), .B(\stack[6][1] ), .Z(n17431) );
  NANDN U18077 ( .A(n17471), .B(\stack[7][1] ), .Z(n17430) );
  NAND U18078 ( .A(n17431), .B(n17430), .Z(n2623) );
  NANDN U18079 ( .A(n2967), .B(\stack[5][1] ), .Z(n17433) );
  NANDN U18080 ( .A(n17472), .B(\stack[7][1] ), .Z(n17432) );
  AND U18081 ( .A(n17433), .B(n17432), .Z(n17435) );
  NANDN U18082 ( .A(n17475), .B(\stack[6][1] ), .Z(n17434) );
  NAND U18083 ( .A(n17435), .B(n17434), .Z(n2624) );
  NANDN U18084 ( .A(n2967), .B(\stack[4][1] ), .Z(n17437) );
  NANDN U18085 ( .A(n17472), .B(\stack[6][1] ), .Z(n17436) );
  AND U18086 ( .A(n17437), .B(n17436), .Z(n17439) );
  NANDN U18087 ( .A(n17475), .B(\stack[5][1] ), .Z(n17438) );
  NAND U18088 ( .A(n17439), .B(n17438), .Z(n2625) );
  NANDN U18089 ( .A(n2967), .B(\stack[3][1] ), .Z(n17441) );
  NANDN U18090 ( .A(n17472), .B(\stack[5][1] ), .Z(n17440) );
  AND U18091 ( .A(n17441), .B(n17440), .Z(n17443) );
  NANDN U18092 ( .A(n17475), .B(\stack[4][1] ), .Z(n17442) );
  NAND U18093 ( .A(n17443), .B(n17442), .Z(n2626) );
  NANDN U18094 ( .A(n2967), .B(\stack[2][1] ), .Z(n17445) );
  NANDN U18095 ( .A(n17472), .B(\stack[4][1] ), .Z(n17444) );
  AND U18096 ( .A(n17445), .B(n17444), .Z(n17447) );
  NANDN U18097 ( .A(n17475), .B(\stack[3][1] ), .Z(n17446) );
  NAND U18098 ( .A(n17447), .B(n17446), .Z(n2627) );
  NANDN U18099 ( .A(n2969), .B(n17471), .Z(n17449) );
  NANDN U18100 ( .A(n17472), .B(\stack[3][1] ), .Z(n17448) );
  AND U18101 ( .A(n17449), .B(n17448), .Z(n17451) );
  NANDN U18102 ( .A(n17475), .B(\stack[2][1] ), .Z(n17450) );
  NAND U18103 ( .A(n17451), .B(n17450), .Z(n2628) );
  NANDN U18104 ( .A(n2995), .B(n17471), .Z(n17453) );
  NANDN U18105 ( .A(n17472), .B(\stack[2][1] ), .Z(n17452) );
  AND U18106 ( .A(n17453), .B(n17452), .Z(n17455) );
  OR U18107 ( .A(n17475), .B(n2969), .Z(n17454) );
  NAND U18108 ( .A(n17455), .B(n17454), .Z(n2629) );
  XNOR U18109 ( .A(n17457), .B(n17456), .Z(n17459) );
  NAND U18110 ( .A(n17459), .B(n17458), .Z(n17464) );
  NANDN U18111 ( .A(n2995), .B(n17479), .Z(n17460) );
  NANDN U18112 ( .A(n17461), .B(n17460), .Z(n17462) );
  NANDN U18113 ( .A(n2969), .B(n17462), .Z(n17463) );
  AND U18114 ( .A(n17464), .B(n17463), .Z(n17466) );
  NANDN U18115 ( .A(n2967), .B(x[1]), .Z(n17465) );
  AND U18116 ( .A(n17466), .B(n17465), .Z(n17470) );
  NANDN U18117 ( .A(n2995), .B(n17467), .Z(n17468) );
  NAND U18118 ( .A(n17470), .B(n17469), .Z(n2630) );
  NANDN U18119 ( .A(n2994), .B(n17471), .Z(n17474) );
  NANDN U18120 ( .A(n17472), .B(\stack[2][0] ), .Z(n17473) );
  AND U18121 ( .A(n17474), .B(n17473), .Z(n17477) );
  OR U18122 ( .A(n17475), .B(n2968), .Z(n17476) );
  NAND U18123 ( .A(n17477), .B(n17476), .Z(n2631) );
  NANDN U18124 ( .A(n17479), .B(n17478), .Z(n17480) );
  ANDN U18125 ( .B(n17480), .A(n2968), .Z(n17482) );
  NANDN U18126 ( .A(n17482), .B(n17481), .Z(n17486) );
  NANDN U18127 ( .A(n17483), .B(n17482), .Z(n17484) );
  NANDN U18128 ( .A(o[0]), .B(n17484), .Z(n17485) );
  NAND U18129 ( .A(n17486), .B(n17485), .Z(n17489) );
  NANDN U18130 ( .A(n2967), .B(x[0]), .Z(n17487) );
  NAND U18131 ( .A(n17489), .B(n17488), .Z(n2632) );
endmodule

