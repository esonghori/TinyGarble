
module mult_N64_CC32 ( clk, rst, a, b, c );
  input [63:0] a;
  input [1:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822;
  wire   [127:0] sreg;

  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U5 ( .A(n797), .B(n796), .Z(n1) );
  XOR U6 ( .A(n796), .B(n797), .Z(n2) );
  NAND U7 ( .A(n2), .B(n795), .Z(n3) );
  NAND U8 ( .A(n1), .B(n3), .Z(n804) );
  NAND U9 ( .A(n405), .B(n403), .Z(n4) );
  XOR U10 ( .A(n403), .B(n405), .Z(n5) );
  NAND U11 ( .A(n5), .B(n404), .Z(n6) );
  NAND U12 ( .A(n4), .B(n6), .Z(n411) );
  NAND U13 ( .A(n426), .B(n425), .Z(n7) );
  XOR U14 ( .A(n425), .B(n426), .Z(n8) );
  NAND U15 ( .A(n8), .B(n424), .Z(n9) );
  NAND U16 ( .A(n7), .B(n9), .Z(n432) );
  NAND U17 ( .A(n447), .B(n446), .Z(n10) );
  XOR U18 ( .A(n446), .B(n447), .Z(n11) );
  NAND U19 ( .A(n11), .B(n445), .Z(n12) );
  NAND U20 ( .A(n10), .B(n12), .Z(n453) );
  NAND U21 ( .A(n468), .B(n467), .Z(n13) );
  XOR U22 ( .A(n467), .B(n468), .Z(n14) );
  NAND U23 ( .A(n14), .B(n466), .Z(n15) );
  NAND U24 ( .A(n13), .B(n15), .Z(n474) );
  NAND U25 ( .A(n489), .B(n487), .Z(n16) );
  XOR U26 ( .A(n487), .B(n489), .Z(n17) );
  NAND U27 ( .A(n17), .B(n488), .Z(n18) );
  NAND U28 ( .A(n16), .B(n18), .Z(n495) );
  NAND U29 ( .A(n510), .B(n509), .Z(n19) );
  XOR U30 ( .A(n509), .B(n510), .Z(n20) );
  NAND U31 ( .A(n20), .B(n508), .Z(n21) );
  NAND U32 ( .A(n19), .B(n21), .Z(n516) );
  NAND U33 ( .A(n531), .B(n530), .Z(n22) );
  XOR U34 ( .A(n530), .B(n531), .Z(n23) );
  NAND U35 ( .A(n23), .B(n529), .Z(n24) );
  NAND U36 ( .A(n22), .B(n24), .Z(n537) );
  NAND U37 ( .A(n552), .B(n551), .Z(n25) );
  XOR U38 ( .A(n551), .B(n552), .Z(n26) );
  NAND U39 ( .A(n26), .B(n550), .Z(n27) );
  NAND U40 ( .A(n25), .B(n27), .Z(n558) );
  NAND U41 ( .A(n573), .B(n572), .Z(n28) );
  XOR U42 ( .A(n572), .B(n573), .Z(n29) );
  NAND U43 ( .A(n29), .B(n571), .Z(n30) );
  NAND U44 ( .A(n28), .B(n30), .Z(n579) );
  NAND U45 ( .A(n594), .B(n593), .Z(n31) );
  XOR U46 ( .A(n593), .B(n594), .Z(n32) );
  NAND U47 ( .A(n32), .B(n592), .Z(n33) );
  NAND U48 ( .A(n31), .B(n33), .Z(n600) );
  NAND U49 ( .A(n615), .B(n614), .Z(n34) );
  XOR U50 ( .A(n614), .B(n615), .Z(n35) );
  NAND U51 ( .A(n35), .B(n613), .Z(n36) );
  NAND U52 ( .A(n34), .B(n36), .Z(n621) );
  NAND U53 ( .A(n636), .B(n635), .Z(n37) );
  XOR U54 ( .A(n635), .B(n636), .Z(n38) );
  NAND U55 ( .A(n38), .B(n634), .Z(n39) );
  NAND U56 ( .A(n37), .B(n39), .Z(n642) );
  NAND U57 ( .A(n657), .B(n656), .Z(n40) );
  XOR U58 ( .A(n656), .B(n657), .Z(n41) );
  NAND U59 ( .A(n41), .B(n655), .Z(n42) );
  NAND U60 ( .A(n40), .B(n42), .Z(n663) );
  NAND U61 ( .A(n678), .B(n677), .Z(n43) );
  XOR U62 ( .A(n677), .B(n678), .Z(n44) );
  NAND U63 ( .A(n44), .B(n676), .Z(n45) );
  NAND U64 ( .A(n43), .B(n45), .Z(n684) );
  NAND U65 ( .A(n699), .B(n698), .Z(n46) );
  XOR U66 ( .A(n698), .B(n699), .Z(n47) );
  NAND U67 ( .A(n47), .B(n697), .Z(n48) );
  NAND U68 ( .A(n46), .B(n48), .Z(n705) );
  NAND U69 ( .A(n720), .B(n719), .Z(n49) );
  XOR U70 ( .A(n719), .B(n720), .Z(n50) );
  NAND U71 ( .A(n50), .B(n718), .Z(n51) );
  NAND U72 ( .A(n49), .B(n51), .Z(n726) );
  NAND U73 ( .A(n741), .B(n740), .Z(n52) );
  XOR U74 ( .A(n740), .B(n741), .Z(n53) );
  NAND U75 ( .A(n53), .B(n739), .Z(n54) );
  NAND U76 ( .A(n52), .B(n54), .Z(n747) );
  NAND U77 ( .A(n762), .B(n761), .Z(n55) );
  XOR U78 ( .A(n761), .B(n762), .Z(n56) );
  NAND U79 ( .A(n56), .B(n760), .Z(n57) );
  NAND U80 ( .A(n55), .B(n57), .Z(n768) );
  NAND U81 ( .A(n783), .B(n782), .Z(n58) );
  XOR U82 ( .A(n782), .B(n783), .Z(n59) );
  NAND U83 ( .A(n59), .B(n781), .Z(n60) );
  NAND U84 ( .A(n58), .B(n60), .Z(n789) );
  XOR U85 ( .A(n805), .B(n803), .Z(n61) );
  NAND U86 ( .A(n61), .B(n804), .Z(n62) );
  NAND U87 ( .A(n805), .B(n803), .Z(n63) );
  AND U88 ( .A(n62), .B(n63), .Z(n814) );
  NAND U89 ( .A(sreg[66]), .B(n401), .Z(n64) );
  XOR U90 ( .A(n401), .B(sreg[66]), .Z(n65) );
  NAND U91 ( .A(n65), .B(n400), .Z(n66) );
  NAND U92 ( .A(n64), .B(n66), .Z(n407) );
  NAND U93 ( .A(sreg[69]), .B(n422), .Z(n67) );
  XOR U94 ( .A(n422), .B(sreg[69]), .Z(n68) );
  NAND U95 ( .A(n68), .B(n421), .Z(n69) );
  NAND U96 ( .A(n67), .B(n69), .Z(n428) );
  NAND U97 ( .A(sreg[72]), .B(n443), .Z(n70) );
  XOR U98 ( .A(n443), .B(sreg[72]), .Z(n71) );
  NAND U99 ( .A(n71), .B(n442), .Z(n72) );
  NAND U100 ( .A(n70), .B(n72), .Z(n449) );
  NAND U101 ( .A(sreg[75]), .B(n463), .Z(n73) );
  XOR U102 ( .A(n463), .B(sreg[75]), .Z(n74) );
  NANDN U103 ( .A(n464), .B(n74), .Z(n75) );
  NAND U104 ( .A(n73), .B(n75), .Z(n470) );
  NAND U105 ( .A(sreg[78]), .B(n485), .Z(n76) );
  XOR U106 ( .A(n485), .B(sreg[78]), .Z(n77) );
  NAND U107 ( .A(n77), .B(n484), .Z(n78) );
  NAND U108 ( .A(n76), .B(n78), .Z(n491) );
  NAND U109 ( .A(sreg[81]), .B(n506), .Z(n79) );
  XOR U110 ( .A(n506), .B(sreg[81]), .Z(n80) );
  NAND U111 ( .A(n80), .B(n505), .Z(n81) );
  NAND U112 ( .A(n79), .B(n81), .Z(n512) );
  NAND U113 ( .A(sreg[84]), .B(n527), .Z(n82) );
  XOR U114 ( .A(n527), .B(sreg[84]), .Z(n83) );
  NAND U115 ( .A(n83), .B(n526), .Z(n84) );
  NAND U116 ( .A(n82), .B(n84), .Z(n533) );
  NAND U117 ( .A(sreg[87]), .B(n548), .Z(n85) );
  XOR U118 ( .A(n548), .B(sreg[87]), .Z(n86) );
  NAND U119 ( .A(n86), .B(n547), .Z(n87) );
  NAND U120 ( .A(n85), .B(n87), .Z(n554) );
  NAND U121 ( .A(sreg[90]), .B(n569), .Z(n88) );
  XOR U122 ( .A(n569), .B(sreg[90]), .Z(n89) );
  NAND U123 ( .A(n89), .B(n568), .Z(n90) );
  NAND U124 ( .A(n88), .B(n90), .Z(n575) );
  NAND U125 ( .A(sreg[93]), .B(n590), .Z(n91) );
  XOR U126 ( .A(n590), .B(sreg[93]), .Z(n92) );
  NAND U127 ( .A(n92), .B(n589), .Z(n93) );
  NAND U128 ( .A(n91), .B(n93), .Z(n596) );
  NAND U129 ( .A(sreg[96]), .B(n611), .Z(n94) );
  XOR U130 ( .A(n611), .B(sreg[96]), .Z(n95) );
  NAND U131 ( .A(n95), .B(n610), .Z(n96) );
  NAND U132 ( .A(n94), .B(n96), .Z(n617) );
  NAND U133 ( .A(sreg[99]), .B(n632), .Z(n97) );
  XOR U134 ( .A(n632), .B(sreg[99]), .Z(n98) );
  NAND U135 ( .A(n98), .B(n631), .Z(n99) );
  NAND U136 ( .A(n97), .B(n99), .Z(n638) );
  NAND U137 ( .A(sreg[102]), .B(n653), .Z(n100) );
  XOR U138 ( .A(n653), .B(sreg[102]), .Z(n101) );
  NAND U139 ( .A(n101), .B(n652), .Z(n102) );
  NAND U140 ( .A(n100), .B(n102), .Z(n659) );
  NAND U141 ( .A(sreg[105]), .B(n674), .Z(n103) );
  XOR U142 ( .A(n674), .B(sreg[105]), .Z(n104) );
  NAND U143 ( .A(n104), .B(n673), .Z(n105) );
  NAND U144 ( .A(n103), .B(n105), .Z(n680) );
  NAND U145 ( .A(sreg[108]), .B(n695), .Z(n106) );
  XOR U146 ( .A(n695), .B(sreg[108]), .Z(n107) );
  NAND U147 ( .A(n107), .B(n694), .Z(n108) );
  NAND U148 ( .A(n106), .B(n108), .Z(n701) );
  NAND U149 ( .A(sreg[111]), .B(n716), .Z(n109) );
  XOR U150 ( .A(n716), .B(sreg[111]), .Z(n110) );
  NAND U151 ( .A(n110), .B(n715), .Z(n111) );
  NAND U152 ( .A(n109), .B(n111), .Z(n722) );
  NAND U153 ( .A(sreg[114]), .B(n737), .Z(n112) );
  XOR U154 ( .A(n737), .B(sreg[114]), .Z(n113) );
  NAND U155 ( .A(n113), .B(n736), .Z(n114) );
  NAND U156 ( .A(n112), .B(n114), .Z(n743) );
  NAND U157 ( .A(sreg[117]), .B(n758), .Z(n115) );
  XOR U158 ( .A(n758), .B(sreg[117]), .Z(n116) );
  NAND U159 ( .A(n116), .B(n757), .Z(n117) );
  NAND U160 ( .A(n115), .B(n117), .Z(n764) );
  NAND U161 ( .A(sreg[120]), .B(n779), .Z(n118) );
  XOR U162 ( .A(n779), .B(sreg[120]), .Z(n119) );
  NAND U163 ( .A(n119), .B(n778), .Z(n120) );
  NAND U164 ( .A(n118), .B(n120), .Z(n785) );
  NAND U165 ( .A(sreg[123]), .B(n800), .Z(n121) );
  XOR U166 ( .A(n800), .B(sreg[123]), .Z(n122) );
  NAND U167 ( .A(n122), .B(n799), .Z(n123) );
  NAND U168 ( .A(n121), .B(n123), .Z(n806) );
  NAND U169 ( .A(n412), .B(n411), .Z(n124) );
  XOR U170 ( .A(n411), .B(n412), .Z(n125) );
  NAND U171 ( .A(n125), .B(n410), .Z(n126) );
  NAND U172 ( .A(n124), .B(n126), .Z(n418) );
  NAND U173 ( .A(n433), .B(n431), .Z(n127) );
  XOR U174 ( .A(n431), .B(n433), .Z(n128) );
  NAND U175 ( .A(n128), .B(n432), .Z(n129) );
  NAND U176 ( .A(n127), .B(n129), .Z(n439) );
  NAND U177 ( .A(n454), .B(n453), .Z(n130) );
  XOR U178 ( .A(n453), .B(n454), .Z(n131) );
  NAND U179 ( .A(n131), .B(n452), .Z(n132) );
  NAND U180 ( .A(n130), .B(n132), .Z(n460) );
  NAND U181 ( .A(n475), .B(n474), .Z(n133) );
  XOR U182 ( .A(n474), .B(n475), .Z(n134) );
  NAND U183 ( .A(n134), .B(n473), .Z(n135) );
  NAND U184 ( .A(n133), .B(n135), .Z(n481) );
  NAND U185 ( .A(n496), .B(n495), .Z(n136) );
  XOR U186 ( .A(n495), .B(n496), .Z(n137) );
  NAND U187 ( .A(n137), .B(n494), .Z(n138) );
  NAND U188 ( .A(n136), .B(n138), .Z(n502) );
  NAND U189 ( .A(n517), .B(n515), .Z(n139) );
  XOR U190 ( .A(n515), .B(n517), .Z(n140) );
  NAND U191 ( .A(n140), .B(n516), .Z(n141) );
  NAND U192 ( .A(n139), .B(n141), .Z(n523) );
  NAND U193 ( .A(n538), .B(n537), .Z(n142) );
  XOR U194 ( .A(n537), .B(n538), .Z(n143) );
  NAND U195 ( .A(n143), .B(n536), .Z(n144) );
  NAND U196 ( .A(n142), .B(n144), .Z(n544) );
  NAND U197 ( .A(n559), .B(n558), .Z(n145) );
  XOR U198 ( .A(n558), .B(n559), .Z(n146) );
  NAND U199 ( .A(n146), .B(n557), .Z(n147) );
  NAND U200 ( .A(n145), .B(n147), .Z(n565) );
  NAND U201 ( .A(n580), .B(n579), .Z(n148) );
  XOR U202 ( .A(n579), .B(n580), .Z(n149) );
  NAND U203 ( .A(n149), .B(n578), .Z(n150) );
  NAND U204 ( .A(n148), .B(n150), .Z(n586) );
  NAND U205 ( .A(n601), .B(n600), .Z(n151) );
  XOR U206 ( .A(n600), .B(n601), .Z(n152) );
  NAND U207 ( .A(n152), .B(n599), .Z(n153) );
  NAND U208 ( .A(n151), .B(n153), .Z(n607) );
  NAND U209 ( .A(n622), .B(n621), .Z(n154) );
  XOR U210 ( .A(n621), .B(n622), .Z(n155) );
  NAND U211 ( .A(n155), .B(n620), .Z(n156) );
  NAND U212 ( .A(n154), .B(n156), .Z(n628) );
  NAND U213 ( .A(n643), .B(n642), .Z(n157) );
  XOR U214 ( .A(n642), .B(n643), .Z(n158) );
  NAND U215 ( .A(n158), .B(n641), .Z(n159) );
  NAND U216 ( .A(n157), .B(n159), .Z(n649) );
  NAND U217 ( .A(n664), .B(n663), .Z(n160) );
  XOR U218 ( .A(n663), .B(n664), .Z(n161) );
  NAND U219 ( .A(n161), .B(n662), .Z(n162) );
  NAND U220 ( .A(n160), .B(n162), .Z(n670) );
  NAND U221 ( .A(n685), .B(n684), .Z(n163) );
  XOR U222 ( .A(n684), .B(n685), .Z(n164) );
  NAND U223 ( .A(n164), .B(n683), .Z(n165) );
  NAND U224 ( .A(n163), .B(n165), .Z(n691) );
  NAND U225 ( .A(n706), .B(n705), .Z(n166) );
  XOR U226 ( .A(n705), .B(n706), .Z(n167) );
  NAND U227 ( .A(n167), .B(n704), .Z(n168) );
  NAND U228 ( .A(n166), .B(n168), .Z(n712) );
  NAND U229 ( .A(n727), .B(n726), .Z(n169) );
  XOR U230 ( .A(n726), .B(n727), .Z(n170) );
  NAND U231 ( .A(n170), .B(n725), .Z(n171) );
  NAND U232 ( .A(n169), .B(n171), .Z(n733) );
  NAND U233 ( .A(n748), .B(n747), .Z(n172) );
  XOR U234 ( .A(n747), .B(n748), .Z(n173) );
  NAND U235 ( .A(n173), .B(n746), .Z(n174) );
  NAND U236 ( .A(n172), .B(n174), .Z(n754) );
  NAND U237 ( .A(n769), .B(n768), .Z(n175) );
  XOR U238 ( .A(n768), .B(n769), .Z(n176) );
  NAND U239 ( .A(n176), .B(n767), .Z(n177) );
  NAND U240 ( .A(n175), .B(n177), .Z(n775) );
  NAND U241 ( .A(n790), .B(n789), .Z(n178) );
  XOR U242 ( .A(n789), .B(n790), .Z(n179) );
  NAND U243 ( .A(n179), .B(n788), .Z(n180) );
  NAND U244 ( .A(n178), .B(n180), .Z(n796) );
  NAND U245 ( .A(sreg[64]), .B(n380), .Z(n181) );
  XOR U246 ( .A(n380), .B(sreg[64]), .Z(n182) );
  NANDN U247 ( .A(n381), .B(n182), .Z(n183) );
  NAND U248 ( .A(n181), .B(n183), .Z(n393) );
  NAND U249 ( .A(sreg[67]), .B(n407), .Z(n184) );
  XOR U250 ( .A(n407), .B(sreg[67]), .Z(n185) );
  NANDN U251 ( .A(n408), .B(n185), .Z(n186) );
  NAND U252 ( .A(n184), .B(n186), .Z(n414) );
  NAND U253 ( .A(sreg[70]), .B(n429), .Z(n187) );
  XOR U254 ( .A(n429), .B(sreg[70]), .Z(n188) );
  NAND U255 ( .A(n188), .B(n428), .Z(n189) );
  NAND U256 ( .A(n187), .B(n189), .Z(n435) );
  NAND U257 ( .A(sreg[73]), .B(n450), .Z(n190) );
  XOR U258 ( .A(n450), .B(sreg[73]), .Z(n191) );
  NAND U259 ( .A(n191), .B(n449), .Z(n192) );
  NAND U260 ( .A(n190), .B(n192), .Z(n456) );
  NAND U261 ( .A(sreg[76]), .B(n471), .Z(n193) );
  XOR U262 ( .A(n471), .B(sreg[76]), .Z(n194) );
  NAND U263 ( .A(n194), .B(n470), .Z(n195) );
  NAND U264 ( .A(n193), .B(n195), .Z(n477) );
  NAND U265 ( .A(sreg[79]), .B(n491), .Z(n196) );
  XOR U266 ( .A(n491), .B(sreg[79]), .Z(n197) );
  NANDN U267 ( .A(n492), .B(n197), .Z(n198) );
  NAND U268 ( .A(n196), .B(n198), .Z(n498) );
  NAND U269 ( .A(sreg[82]), .B(n513), .Z(n199) );
  XOR U270 ( .A(n513), .B(sreg[82]), .Z(n200) );
  NAND U271 ( .A(n200), .B(n512), .Z(n201) );
  NAND U272 ( .A(n199), .B(n201), .Z(n519) );
  NAND U273 ( .A(sreg[85]), .B(n534), .Z(n202) );
  XOR U274 ( .A(n534), .B(sreg[85]), .Z(n203) );
  NAND U275 ( .A(n203), .B(n533), .Z(n204) );
  NAND U276 ( .A(n202), .B(n204), .Z(n540) );
  NAND U277 ( .A(sreg[88]), .B(n555), .Z(n205) );
  XOR U278 ( .A(n555), .B(sreg[88]), .Z(n206) );
  NAND U279 ( .A(n206), .B(n554), .Z(n207) );
  NAND U280 ( .A(n205), .B(n207), .Z(n561) );
  NAND U281 ( .A(sreg[91]), .B(n576), .Z(n208) );
  XOR U282 ( .A(n576), .B(sreg[91]), .Z(n209) );
  NAND U283 ( .A(n209), .B(n575), .Z(n210) );
  NAND U284 ( .A(n208), .B(n210), .Z(n582) );
  NAND U285 ( .A(sreg[94]), .B(n597), .Z(n211) );
  XOR U286 ( .A(n597), .B(sreg[94]), .Z(n212) );
  NAND U287 ( .A(n212), .B(n596), .Z(n213) );
  NAND U288 ( .A(n211), .B(n213), .Z(n603) );
  NAND U289 ( .A(sreg[97]), .B(n618), .Z(n214) );
  XOR U290 ( .A(n618), .B(sreg[97]), .Z(n215) );
  NAND U291 ( .A(n215), .B(n617), .Z(n216) );
  NAND U292 ( .A(n214), .B(n216), .Z(n624) );
  NAND U293 ( .A(sreg[100]), .B(n639), .Z(n217) );
  XOR U294 ( .A(n639), .B(sreg[100]), .Z(n218) );
  NAND U295 ( .A(n218), .B(n638), .Z(n219) );
  NAND U296 ( .A(n217), .B(n219), .Z(n645) );
  NAND U297 ( .A(sreg[103]), .B(n660), .Z(n220) );
  XOR U298 ( .A(n660), .B(sreg[103]), .Z(n221) );
  NAND U299 ( .A(n221), .B(n659), .Z(n222) );
  NAND U300 ( .A(n220), .B(n222), .Z(n666) );
  NAND U301 ( .A(sreg[106]), .B(n681), .Z(n223) );
  XOR U302 ( .A(n681), .B(sreg[106]), .Z(n224) );
  NAND U303 ( .A(n224), .B(n680), .Z(n225) );
  NAND U304 ( .A(n223), .B(n225), .Z(n687) );
  NAND U305 ( .A(sreg[109]), .B(n702), .Z(n226) );
  XOR U306 ( .A(n702), .B(sreg[109]), .Z(n227) );
  NAND U307 ( .A(n227), .B(n701), .Z(n228) );
  NAND U308 ( .A(n226), .B(n228), .Z(n708) );
  NAND U309 ( .A(sreg[112]), .B(n723), .Z(n229) );
  XOR U310 ( .A(n723), .B(sreg[112]), .Z(n230) );
  NAND U311 ( .A(n230), .B(n722), .Z(n231) );
  NAND U312 ( .A(n229), .B(n231), .Z(n729) );
  NAND U313 ( .A(sreg[115]), .B(n744), .Z(n232) );
  XOR U314 ( .A(n744), .B(sreg[115]), .Z(n233) );
  NAND U315 ( .A(n233), .B(n743), .Z(n234) );
  NAND U316 ( .A(n232), .B(n234), .Z(n750) );
  NAND U317 ( .A(sreg[118]), .B(n765), .Z(n235) );
  XOR U318 ( .A(n765), .B(sreg[118]), .Z(n236) );
  NAND U319 ( .A(n236), .B(n764), .Z(n237) );
  NAND U320 ( .A(n235), .B(n237), .Z(n771) );
  NAND U321 ( .A(sreg[121]), .B(n786), .Z(n238) );
  XOR U322 ( .A(n786), .B(sreg[121]), .Z(n239) );
  NAND U323 ( .A(n239), .B(n785), .Z(n240) );
  NAND U324 ( .A(n238), .B(n240), .Z(n792) );
  NAND U325 ( .A(sreg[124]), .B(n806), .Z(n241) );
  XOR U326 ( .A(n806), .B(sreg[124]), .Z(n242) );
  NANDN U327 ( .A(n807), .B(n242), .Z(n243) );
  NAND U328 ( .A(n241), .B(n243), .Z(n809) );
  NAND U329 ( .A(n398), .B(n397), .Z(n244) );
  XOR U330 ( .A(n397), .B(n398), .Z(n245) );
  NANDN U331 ( .A(n396), .B(n245), .Z(n246) );
  NAND U332 ( .A(n244), .B(n246), .Z(n404) );
  NAND U333 ( .A(n419), .B(n418), .Z(n247) );
  XOR U334 ( .A(n418), .B(n419), .Z(n248) );
  NAND U335 ( .A(n248), .B(n417), .Z(n249) );
  NAND U336 ( .A(n247), .B(n249), .Z(n425) );
  NAND U337 ( .A(n440), .B(n439), .Z(n250) );
  XOR U338 ( .A(n439), .B(n440), .Z(n251) );
  NAND U339 ( .A(n251), .B(n438), .Z(n252) );
  NAND U340 ( .A(n250), .B(n252), .Z(n446) );
  NAND U341 ( .A(n461), .B(n459), .Z(n253) );
  XOR U342 ( .A(n459), .B(n461), .Z(n254) );
  NAND U343 ( .A(n254), .B(n460), .Z(n255) );
  NAND U344 ( .A(n253), .B(n255), .Z(n467) );
  NAND U345 ( .A(n482), .B(n481), .Z(n256) );
  XOR U346 ( .A(n481), .B(n482), .Z(n257) );
  NAND U347 ( .A(n257), .B(n480), .Z(n258) );
  NAND U348 ( .A(n256), .B(n258), .Z(n488) );
  NAND U349 ( .A(n503), .B(n502), .Z(n259) );
  XOR U350 ( .A(n502), .B(n503), .Z(n260) );
  NAND U351 ( .A(n260), .B(n501), .Z(n261) );
  NAND U352 ( .A(n259), .B(n261), .Z(n509) );
  NAND U353 ( .A(n524), .B(n523), .Z(n262) );
  XOR U354 ( .A(n523), .B(n524), .Z(n263) );
  NAND U355 ( .A(n263), .B(n522), .Z(n264) );
  NAND U356 ( .A(n262), .B(n264), .Z(n530) );
  NAND U357 ( .A(n545), .B(n544), .Z(n265) );
  XOR U358 ( .A(n544), .B(n545), .Z(n266) );
  NAND U359 ( .A(n266), .B(n543), .Z(n267) );
  NAND U360 ( .A(n265), .B(n267), .Z(n551) );
  NAND U361 ( .A(n566), .B(n565), .Z(n268) );
  XOR U362 ( .A(n565), .B(n566), .Z(n269) );
  NAND U363 ( .A(n269), .B(n564), .Z(n270) );
  NAND U364 ( .A(n268), .B(n270), .Z(n572) );
  NAND U365 ( .A(n587), .B(n586), .Z(n271) );
  XOR U366 ( .A(n586), .B(n587), .Z(n272) );
  NAND U367 ( .A(n272), .B(n585), .Z(n273) );
  NAND U368 ( .A(n271), .B(n273), .Z(n593) );
  NAND U369 ( .A(n608), .B(n607), .Z(n274) );
  XOR U370 ( .A(n607), .B(n608), .Z(n275) );
  NAND U371 ( .A(n275), .B(n606), .Z(n276) );
  NAND U372 ( .A(n274), .B(n276), .Z(n614) );
  NAND U373 ( .A(n629), .B(n628), .Z(n277) );
  XOR U374 ( .A(n628), .B(n629), .Z(n278) );
  NAND U375 ( .A(n278), .B(n627), .Z(n279) );
  NAND U376 ( .A(n277), .B(n279), .Z(n635) );
  NAND U377 ( .A(n650), .B(n649), .Z(n280) );
  XOR U378 ( .A(n649), .B(n650), .Z(n281) );
  NAND U379 ( .A(n281), .B(n648), .Z(n282) );
  NAND U380 ( .A(n280), .B(n282), .Z(n656) );
  NAND U381 ( .A(n671), .B(n670), .Z(n283) );
  XOR U382 ( .A(n670), .B(n671), .Z(n284) );
  NAND U383 ( .A(n284), .B(n669), .Z(n285) );
  NAND U384 ( .A(n283), .B(n285), .Z(n677) );
  NAND U385 ( .A(n692), .B(n691), .Z(n286) );
  XOR U386 ( .A(n691), .B(n692), .Z(n287) );
  NAND U387 ( .A(n287), .B(n690), .Z(n288) );
  NAND U388 ( .A(n286), .B(n288), .Z(n698) );
  NAND U389 ( .A(n713), .B(n712), .Z(n289) );
  XOR U390 ( .A(n712), .B(n713), .Z(n290) );
  NAND U391 ( .A(n290), .B(n711), .Z(n291) );
  NAND U392 ( .A(n289), .B(n291), .Z(n719) );
  NAND U393 ( .A(n734), .B(n733), .Z(n292) );
  XOR U394 ( .A(n733), .B(n734), .Z(n293) );
  NAND U395 ( .A(n293), .B(n732), .Z(n294) );
  NAND U396 ( .A(n292), .B(n294), .Z(n740) );
  NAND U397 ( .A(n755), .B(n754), .Z(n295) );
  XOR U398 ( .A(n754), .B(n755), .Z(n296) );
  NAND U399 ( .A(n296), .B(n753), .Z(n297) );
  NAND U400 ( .A(n295), .B(n297), .Z(n761) );
  NAND U401 ( .A(n776), .B(n775), .Z(n298) );
  XOR U402 ( .A(n775), .B(n776), .Z(n299) );
  NAND U403 ( .A(n299), .B(n774), .Z(n300) );
  NAND U404 ( .A(n298), .B(n300), .Z(n782) );
  NAND U405 ( .A(sreg[65]), .B(n393), .Z(n301) );
  XOR U406 ( .A(n393), .B(sreg[65]), .Z(n302) );
  NANDN U407 ( .A(n394), .B(n302), .Z(n303) );
  NAND U408 ( .A(n301), .B(n303), .Z(n400) );
  NAND U409 ( .A(sreg[68]), .B(n415), .Z(n304) );
  XOR U410 ( .A(n415), .B(sreg[68]), .Z(n305) );
  NAND U411 ( .A(n305), .B(n414), .Z(n306) );
  NAND U412 ( .A(n304), .B(n306), .Z(n421) );
  NAND U413 ( .A(sreg[71]), .B(n435), .Z(n307) );
  XOR U414 ( .A(n435), .B(sreg[71]), .Z(n308) );
  NANDN U415 ( .A(n436), .B(n308), .Z(n309) );
  NAND U416 ( .A(n307), .B(n309), .Z(n442) );
  NAND U417 ( .A(sreg[74]), .B(n457), .Z(n310) );
  XOR U418 ( .A(n457), .B(sreg[74]), .Z(n311) );
  NAND U419 ( .A(n311), .B(n456), .Z(n312) );
  NAND U420 ( .A(n310), .B(n312), .Z(n463) );
  NAND U421 ( .A(sreg[77]), .B(n478), .Z(n313) );
  XOR U422 ( .A(n478), .B(sreg[77]), .Z(n314) );
  NAND U423 ( .A(n314), .B(n477), .Z(n315) );
  NAND U424 ( .A(n313), .B(n315), .Z(n484) );
  NAND U425 ( .A(sreg[80]), .B(n499), .Z(n316) );
  XOR U426 ( .A(n499), .B(sreg[80]), .Z(n317) );
  NAND U427 ( .A(n317), .B(n498), .Z(n318) );
  NAND U428 ( .A(n316), .B(n318), .Z(n505) );
  NAND U429 ( .A(sreg[83]), .B(n519), .Z(n319) );
  XOR U430 ( .A(n519), .B(sreg[83]), .Z(n320) );
  NANDN U431 ( .A(n520), .B(n320), .Z(n321) );
  NAND U432 ( .A(n319), .B(n321), .Z(n526) );
  NAND U433 ( .A(sreg[86]), .B(n541), .Z(n322) );
  XOR U434 ( .A(n541), .B(sreg[86]), .Z(n323) );
  NAND U435 ( .A(n323), .B(n540), .Z(n324) );
  NAND U436 ( .A(n322), .B(n324), .Z(n547) );
  NAND U437 ( .A(sreg[89]), .B(n562), .Z(n325) );
  XOR U438 ( .A(n562), .B(sreg[89]), .Z(n326) );
  NAND U439 ( .A(n326), .B(n561), .Z(n327) );
  NAND U440 ( .A(n325), .B(n327), .Z(n568) );
  NAND U441 ( .A(sreg[92]), .B(n583), .Z(n328) );
  XOR U442 ( .A(n583), .B(sreg[92]), .Z(n329) );
  NAND U443 ( .A(n329), .B(n582), .Z(n330) );
  NAND U444 ( .A(n328), .B(n330), .Z(n589) );
  NAND U445 ( .A(sreg[95]), .B(n604), .Z(n331) );
  XOR U446 ( .A(n604), .B(sreg[95]), .Z(n332) );
  NAND U447 ( .A(n332), .B(n603), .Z(n333) );
  NAND U448 ( .A(n331), .B(n333), .Z(n610) );
  NAND U449 ( .A(sreg[98]), .B(n625), .Z(n334) );
  XOR U450 ( .A(n625), .B(sreg[98]), .Z(n335) );
  NAND U451 ( .A(n335), .B(n624), .Z(n336) );
  NAND U452 ( .A(n334), .B(n336), .Z(n631) );
  NAND U453 ( .A(sreg[101]), .B(n646), .Z(n337) );
  XOR U454 ( .A(n646), .B(sreg[101]), .Z(n338) );
  NAND U455 ( .A(n338), .B(n645), .Z(n339) );
  NAND U456 ( .A(n337), .B(n339), .Z(n652) );
  NAND U457 ( .A(sreg[104]), .B(n667), .Z(n340) );
  XOR U458 ( .A(n667), .B(sreg[104]), .Z(n341) );
  NAND U459 ( .A(n341), .B(n666), .Z(n342) );
  NAND U460 ( .A(n340), .B(n342), .Z(n673) );
  NAND U461 ( .A(sreg[107]), .B(n688), .Z(n343) );
  XOR U462 ( .A(n688), .B(sreg[107]), .Z(n344) );
  NAND U463 ( .A(n344), .B(n687), .Z(n345) );
  NAND U464 ( .A(n343), .B(n345), .Z(n694) );
  NAND U465 ( .A(sreg[110]), .B(n709), .Z(n346) );
  XOR U466 ( .A(n709), .B(sreg[110]), .Z(n347) );
  NAND U467 ( .A(n347), .B(n708), .Z(n348) );
  NAND U468 ( .A(n346), .B(n348), .Z(n715) );
  NAND U469 ( .A(sreg[113]), .B(n730), .Z(n349) );
  XOR U470 ( .A(n730), .B(sreg[113]), .Z(n350) );
  NAND U471 ( .A(n350), .B(n729), .Z(n351) );
  NAND U472 ( .A(n349), .B(n351), .Z(n736) );
  NAND U473 ( .A(sreg[116]), .B(n751), .Z(n352) );
  XOR U474 ( .A(n751), .B(sreg[116]), .Z(n353) );
  NAND U475 ( .A(n353), .B(n750), .Z(n354) );
  NAND U476 ( .A(n352), .B(n354), .Z(n757) );
  NAND U477 ( .A(sreg[119]), .B(n772), .Z(n355) );
  XOR U478 ( .A(n772), .B(sreg[119]), .Z(n356) );
  NAND U479 ( .A(n356), .B(n771), .Z(n357) );
  NAND U480 ( .A(n355), .B(n357), .Z(n778) );
  NAND U481 ( .A(sreg[122]), .B(n793), .Z(n358) );
  XOR U482 ( .A(n793), .B(sreg[122]), .Z(n359) );
  NAND U483 ( .A(n359), .B(n792), .Z(n360) );
  NAND U484 ( .A(n358), .B(n360), .Z(n799) );
  NAND U485 ( .A(sreg[125]), .B(n810), .Z(n361) );
  XOR U486 ( .A(n810), .B(sreg[125]), .Z(n362) );
  NAND U487 ( .A(n362), .B(n809), .Z(n363) );
  NAND U488 ( .A(n361), .B(n363), .Z(n820) );
  IV U489 ( .A(b[1]), .Z(n364) );
  IV U490 ( .A(b[0]), .Z(n802) );
  NANDN U491 ( .A(n802), .B(a[0]), .Z(n365) );
  XNOR U492 ( .A(n365), .B(sreg[62]), .Z(c[62]) );
  ANDN U493 ( .B(a[0]), .A(n364), .Z(n376) );
  ANDN U494 ( .B(a[1]), .A(n802), .Z(n389) );
  XNOR U495 ( .A(n376), .B(n389), .Z(n369) );
  XOR U496 ( .A(sreg[63]), .B(n369), .Z(n371) );
  NANDN U497 ( .A(n365), .B(sreg[62]), .Z(n370) );
  XOR U498 ( .A(n371), .B(n370), .Z(c[63]) );
  IV U499 ( .A(n389), .Z(n375) );
  ANDN U500 ( .B(n376), .A(n375), .Z(n386) );
  IV U501 ( .A(n386), .Z(n383) );
  ANDN U502 ( .B(a[2]), .A(n802), .Z(n367) );
  NANDN U503 ( .A(n364), .B(a[1]), .Z(n366) );
  XNOR U504 ( .A(n367), .B(n366), .Z(n368) );
  XOR U505 ( .A(n383), .B(n368), .Z(n381) );
  NANDN U506 ( .A(n369), .B(sreg[63]), .Z(n373) );
  OR U507 ( .A(n371), .B(n370), .Z(n372) );
  NAND U508 ( .A(n373), .B(n372), .Z(n380) );
  XOR U509 ( .A(n380), .B(sreg[64]), .Z(n374) );
  XNOR U510 ( .A(n381), .B(n374), .Z(c[64]) );
  NANDN U511 ( .A(n802), .B(a[3]), .Z(n387) );
  AND U512 ( .A(a[2]), .B(b[1]), .Z(n385) );
  XNOR U513 ( .A(n375), .B(n385), .Z(n378) );
  NANDN U514 ( .A(n376), .B(n389), .Z(n377) );
  NAND U515 ( .A(n378), .B(n377), .Z(n379) );
  XNOR U516 ( .A(n387), .B(n379), .Z(n394) );
  XOR U517 ( .A(n393), .B(sreg[65]), .Z(n382) );
  XNOR U518 ( .A(n394), .B(n382), .Z(c[65]) );
  OR U519 ( .A(n387), .B(n383), .Z(n384) );
  NANDN U520 ( .A(n385), .B(n384), .Z(n391) );
  ANDN U521 ( .B(n387), .A(n386), .Z(n388) );
  NANDN U522 ( .A(n389), .B(n388), .Z(n390) );
  NAND U523 ( .A(n391), .B(n390), .Z(n396) );
  AND U524 ( .A(a[3]), .B(b[1]), .Z(n398) );
  ANDN U525 ( .B(a[4]), .A(n802), .Z(n397) );
  XNOR U526 ( .A(n398), .B(n397), .Z(n392) );
  XOR U527 ( .A(n396), .B(n392), .Z(n401) );
  XOR U528 ( .A(n400), .B(sreg[66]), .Z(n395) );
  XOR U529 ( .A(n401), .B(n395), .Z(c[66]) );
  AND U530 ( .A(a[4]), .B(b[1]), .Z(n405) );
  ANDN U531 ( .B(a[5]), .A(n802), .Z(n403) );
  XOR U532 ( .A(n404), .B(n403), .Z(n399) );
  XNOR U533 ( .A(n405), .B(n399), .Z(n408) );
  XOR U534 ( .A(n407), .B(sreg[67]), .Z(n402) );
  XNOR U535 ( .A(n408), .B(n402), .Z(c[67]) );
  ANDN U536 ( .B(a[6]), .A(n802), .Z(n410) );
  AND U537 ( .A(a[5]), .B(b[1]), .Z(n412) );
  XNOR U538 ( .A(n412), .B(n411), .Z(n406) );
  XNOR U539 ( .A(n410), .B(n406), .Z(n415) );
  XOR U540 ( .A(n414), .B(sreg[68]), .Z(n409) );
  XOR U541 ( .A(n415), .B(n409), .Z(c[68]) );
  ANDN U542 ( .B(a[7]), .A(n802), .Z(n417) );
  AND U543 ( .A(a[6]), .B(b[1]), .Z(n419) );
  XNOR U544 ( .A(n419), .B(n418), .Z(n413) );
  XNOR U545 ( .A(n417), .B(n413), .Z(n422) );
  XOR U546 ( .A(n421), .B(sreg[69]), .Z(n416) );
  XOR U547 ( .A(n422), .B(n416), .Z(c[69]) );
  ANDN U548 ( .B(a[8]), .A(n802), .Z(n424) );
  AND U549 ( .A(a[7]), .B(b[1]), .Z(n426) );
  XNOR U550 ( .A(n426), .B(n425), .Z(n420) );
  XNOR U551 ( .A(n424), .B(n420), .Z(n429) );
  XOR U552 ( .A(n428), .B(sreg[70]), .Z(n423) );
  XOR U553 ( .A(n429), .B(n423), .Z(c[70]) );
  AND U554 ( .A(a[8]), .B(b[1]), .Z(n433) );
  ANDN U555 ( .B(a[9]), .A(n802), .Z(n431) );
  XOR U556 ( .A(n432), .B(n431), .Z(n427) );
  XNOR U557 ( .A(n433), .B(n427), .Z(n436) );
  XOR U558 ( .A(n435), .B(sreg[71]), .Z(n430) );
  XNOR U559 ( .A(n436), .B(n430), .Z(c[71]) );
  ANDN U560 ( .B(a[10]), .A(n802), .Z(n438) );
  AND U561 ( .A(a[9]), .B(b[1]), .Z(n440) );
  XNOR U562 ( .A(n440), .B(n439), .Z(n434) );
  XNOR U563 ( .A(n438), .B(n434), .Z(n443) );
  XOR U564 ( .A(n442), .B(sreg[72]), .Z(n437) );
  XOR U565 ( .A(n443), .B(n437), .Z(c[72]) );
  ANDN U566 ( .B(a[11]), .A(n802), .Z(n445) );
  AND U567 ( .A(a[10]), .B(b[1]), .Z(n447) );
  XNOR U568 ( .A(n447), .B(n446), .Z(n441) );
  XNOR U569 ( .A(n445), .B(n441), .Z(n450) );
  XOR U570 ( .A(n449), .B(sreg[73]), .Z(n444) );
  XOR U571 ( .A(n450), .B(n444), .Z(c[73]) );
  ANDN U572 ( .B(a[12]), .A(n802), .Z(n452) );
  AND U573 ( .A(a[11]), .B(b[1]), .Z(n454) );
  XNOR U574 ( .A(n454), .B(n453), .Z(n448) );
  XNOR U575 ( .A(n452), .B(n448), .Z(n457) );
  XOR U576 ( .A(n456), .B(sreg[74]), .Z(n451) );
  XOR U577 ( .A(n457), .B(n451), .Z(c[74]) );
  AND U578 ( .A(a[12]), .B(b[1]), .Z(n461) );
  ANDN U579 ( .B(a[13]), .A(n802), .Z(n459) );
  XOR U580 ( .A(n460), .B(n459), .Z(n455) );
  XNOR U581 ( .A(n461), .B(n455), .Z(n464) );
  XOR U582 ( .A(n463), .B(sreg[75]), .Z(n458) );
  XNOR U583 ( .A(n464), .B(n458), .Z(c[75]) );
  ANDN U584 ( .B(a[14]), .A(n802), .Z(n466) );
  AND U585 ( .A(a[13]), .B(b[1]), .Z(n468) );
  XNOR U586 ( .A(n468), .B(n467), .Z(n462) );
  XNOR U587 ( .A(n466), .B(n462), .Z(n471) );
  XOR U588 ( .A(n470), .B(sreg[76]), .Z(n465) );
  XOR U589 ( .A(n471), .B(n465), .Z(c[76]) );
  ANDN U590 ( .B(a[15]), .A(n802), .Z(n473) );
  AND U591 ( .A(a[14]), .B(b[1]), .Z(n475) );
  XNOR U592 ( .A(n475), .B(n474), .Z(n469) );
  XNOR U593 ( .A(n473), .B(n469), .Z(n478) );
  XOR U594 ( .A(n477), .B(sreg[77]), .Z(n472) );
  XOR U595 ( .A(n478), .B(n472), .Z(c[77]) );
  ANDN U596 ( .B(a[16]), .A(n802), .Z(n480) );
  AND U597 ( .A(a[15]), .B(b[1]), .Z(n482) );
  XNOR U598 ( .A(n482), .B(n481), .Z(n476) );
  XNOR U599 ( .A(n480), .B(n476), .Z(n485) );
  XOR U600 ( .A(n484), .B(sreg[78]), .Z(n479) );
  XOR U601 ( .A(n485), .B(n479), .Z(c[78]) );
  AND U602 ( .A(a[16]), .B(b[1]), .Z(n489) );
  ANDN U603 ( .B(a[17]), .A(n802), .Z(n487) );
  XOR U604 ( .A(n488), .B(n487), .Z(n483) );
  XNOR U605 ( .A(n489), .B(n483), .Z(n492) );
  XOR U606 ( .A(n491), .B(sreg[79]), .Z(n486) );
  XNOR U607 ( .A(n492), .B(n486), .Z(c[79]) );
  ANDN U608 ( .B(a[18]), .A(n802), .Z(n494) );
  AND U609 ( .A(a[17]), .B(b[1]), .Z(n496) );
  XNOR U610 ( .A(n496), .B(n495), .Z(n490) );
  XNOR U611 ( .A(n494), .B(n490), .Z(n499) );
  XOR U612 ( .A(n498), .B(sreg[80]), .Z(n493) );
  XOR U613 ( .A(n499), .B(n493), .Z(c[80]) );
  ANDN U614 ( .B(a[19]), .A(n802), .Z(n501) );
  AND U615 ( .A(a[18]), .B(b[1]), .Z(n503) );
  XNOR U616 ( .A(n503), .B(n502), .Z(n497) );
  XNOR U617 ( .A(n501), .B(n497), .Z(n506) );
  XOR U618 ( .A(n505), .B(sreg[81]), .Z(n500) );
  XOR U619 ( .A(n506), .B(n500), .Z(c[81]) );
  ANDN U620 ( .B(a[20]), .A(n802), .Z(n508) );
  AND U621 ( .A(a[19]), .B(b[1]), .Z(n510) );
  XNOR U622 ( .A(n510), .B(n509), .Z(n504) );
  XNOR U623 ( .A(n508), .B(n504), .Z(n513) );
  XOR U624 ( .A(n512), .B(sreg[82]), .Z(n507) );
  XOR U625 ( .A(n513), .B(n507), .Z(c[82]) );
  AND U626 ( .A(a[20]), .B(b[1]), .Z(n517) );
  ANDN U627 ( .B(a[21]), .A(n802), .Z(n515) );
  XOR U628 ( .A(n516), .B(n515), .Z(n511) );
  XNOR U629 ( .A(n517), .B(n511), .Z(n520) );
  XOR U630 ( .A(n519), .B(sreg[83]), .Z(n514) );
  XNOR U631 ( .A(n520), .B(n514), .Z(c[83]) );
  ANDN U632 ( .B(a[22]), .A(n802), .Z(n522) );
  AND U633 ( .A(a[21]), .B(b[1]), .Z(n524) );
  XNOR U634 ( .A(n524), .B(n523), .Z(n518) );
  XNOR U635 ( .A(n522), .B(n518), .Z(n527) );
  XOR U636 ( .A(n526), .B(sreg[84]), .Z(n521) );
  XOR U637 ( .A(n527), .B(n521), .Z(c[84]) );
  ANDN U638 ( .B(a[23]), .A(n802), .Z(n529) );
  AND U639 ( .A(a[22]), .B(b[1]), .Z(n531) );
  XNOR U640 ( .A(n530), .B(n531), .Z(n525) );
  XNOR U641 ( .A(n529), .B(n525), .Z(n534) );
  XOR U642 ( .A(n533), .B(sreg[85]), .Z(n528) );
  XOR U643 ( .A(n534), .B(n528), .Z(c[85]) );
  ANDN U644 ( .B(a[24]), .A(n802), .Z(n536) );
  AND U645 ( .A(a[23]), .B(b[1]), .Z(n538) );
  XNOR U646 ( .A(n538), .B(n537), .Z(n532) );
  XNOR U647 ( .A(n536), .B(n532), .Z(n541) );
  XOR U648 ( .A(n540), .B(sreg[86]), .Z(n535) );
  XOR U649 ( .A(n541), .B(n535), .Z(c[86]) );
  ANDN U650 ( .B(a[25]), .A(n802), .Z(n543) );
  AND U651 ( .A(a[24]), .B(b[1]), .Z(n545) );
  XNOR U652 ( .A(n544), .B(n545), .Z(n539) );
  XNOR U653 ( .A(n543), .B(n539), .Z(n548) );
  XOR U654 ( .A(n547), .B(sreg[87]), .Z(n542) );
  XOR U655 ( .A(n548), .B(n542), .Z(c[87]) );
  ANDN U656 ( .B(a[26]), .A(n802), .Z(n550) );
  AND U657 ( .A(a[25]), .B(b[1]), .Z(n552) );
  XNOR U658 ( .A(n552), .B(n551), .Z(n546) );
  XNOR U659 ( .A(n550), .B(n546), .Z(n555) );
  XOR U660 ( .A(n554), .B(sreg[88]), .Z(n549) );
  XOR U661 ( .A(n555), .B(n549), .Z(c[88]) );
  ANDN U662 ( .B(a[27]), .A(n802), .Z(n557) );
  AND U663 ( .A(a[26]), .B(b[1]), .Z(n559) );
  XNOR U664 ( .A(n559), .B(n558), .Z(n553) );
  XNOR U665 ( .A(n557), .B(n553), .Z(n562) );
  XOR U666 ( .A(n561), .B(sreg[89]), .Z(n556) );
  XOR U667 ( .A(n562), .B(n556), .Z(c[89]) );
  ANDN U668 ( .B(a[28]), .A(n802), .Z(n564) );
  AND U669 ( .A(a[27]), .B(b[1]), .Z(n566) );
  XNOR U670 ( .A(n566), .B(n565), .Z(n560) );
  XNOR U671 ( .A(n564), .B(n560), .Z(n569) );
  XOR U672 ( .A(n568), .B(sreg[90]), .Z(n563) );
  XOR U673 ( .A(n569), .B(n563), .Z(c[90]) );
  ANDN U674 ( .B(a[29]), .A(n802), .Z(n571) );
  AND U675 ( .A(a[28]), .B(b[1]), .Z(n573) );
  XNOR U676 ( .A(n573), .B(n572), .Z(n567) );
  XNOR U677 ( .A(n571), .B(n567), .Z(n576) );
  XOR U678 ( .A(n575), .B(sreg[91]), .Z(n570) );
  XOR U679 ( .A(n576), .B(n570), .Z(c[91]) );
  ANDN U680 ( .B(a[30]), .A(n802), .Z(n578) );
  AND U681 ( .A(a[29]), .B(b[1]), .Z(n580) );
  XNOR U682 ( .A(n580), .B(n579), .Z(n574) );
  XNOR U683 ( .A(n578), .B(n574), .Z(n583) );
  XOR U684 ( .A(n582), .B(sreg[92]), .Z(n577) );
  XOR U685 ( .A(n583), .B(n577), .Z(c[92]) );
  ANDN U686 ( .B(a[31]), .A(n802), .Z(n585) );
  AND U687 ( .A(a[30]), .B(b[1]), .Z(n587) );
  XNOR U688 ( .A(n587), .B(n586), .Z(n581) );
  XNOR U689 ( .A(n585), .B(n581), .Z(n590) );
  XOR U690 ( .A(n589), .B(sreg[93]), .Z(n584) );
  XOR U691 ( .A(n590), .B(n584), .Z(c[93]) );
  ANDN U692 ( .B(a[32]), .A(n802), .Z(n592) );
  AND U693 ( .A(a[31]), .B(b[1]), .Z(n594) );
  XNOR U694 ( .A(n594), .B(n593), .Z(n588) );
  XNOR U695 ( .A(n592), .B(n588), .Z(n597) );
  XOR U696 ( .A(n596), .B(sreg[94]), .Z(n591) );
  XOR U697 ( .A(n597), .B(n591), .Z(c[94]) );
  ANDN U698 ( .B(a[33]), .A(n802), .Z(n599) );
  AND U699 ( .A(a[32]), .B(b[1]), .Z(n601) );
  XNOR U700 ( .A(n601), .B(n600), .Z(n595) );
  XNOR U701 ( .A(n599), .B(n595), .Z(n604) );
  XOR U702 ( .A(n603), .B(sreg[95]), .Z(n598) );
  XOR U703 ( .A(n604), .B(n598), .Z(c[95]) );
  ANDN U704 ( .B(a[34]), .A(n802), .Z(n606) );
  AND U705 ( .A(a[33]), .B(b[1]), .Z(n608) );
  XNOR U706 ( .A(n608), .B(n607), .Z(n602) );
  XNOR U707 ( .A(n606), .B(n602), .Z(n611) );
  XOR U708 ( .A(n610), .B(sreg[96]), .Z(n605) );
  XOR U709 ( .A(n611), .B(n605), .Z(c[96]) );
  ANDN U710 ( .B(a[35]), .A(n802), .Z(n613) );
  AND U711 ( .A(a[34]), .B(b[1]), .Z(n615) );
  XNOR U712 ( .A(n615), .B(n614), .Z(n609) );
  XNOR U713 ( .A(n613), .B(n609), .Z(n618) );
  XOR U714 ( .A(n617), .B(sreg[97]), .Z(n612) );
  XOR U715 ( .A(n618), .B(n612), .Z(c[97]) );
  ANDN U716 ( .B(a[36]), .A(n802), .Z(n620) );
  AND U717 ( .A(a[35]), .B(b[1]), .Z(n622) );
  XNOR U718 ( .A(n622), .B(n621), .Z(n616) );
  XNOR U719 ( .A(n620), .B(n616), .Z(n625) );
  XOR U720 ( .A(n624), .B(sreg[98]), .Z(n619) );
  XOR U721 ( .A(n625), .B(n619), .Z(c[98]) );
  ANDN U722 ( .B(a[37]), .A(n802), .Z(n627) );
  AND U723 ( .A(a[36]), .B(b[1]), .Z(n629) );
  XNOR U724 ( .A(n629), .B(n628), .Z(n623) );
  XNOR U725 ( .A(n627), .B(n623), .Z(n632) );
  XOR U726 ( .A(n631), .B(sreg[99]), .Z(n626) );
  XOR U727 ( .A(n632), .B(n626), .Z(c[99]) );
  ANDN U728 ( .B(a[38]), .A(n802), .Z(n634) );
  AND U729 ( .A(a[37]), .B(b[1]), .Z(n636) );
  XNOR U730 ( .A(n636), .B(n635), .Z(n630) );
  XNOR U731 ( .A(n634), .B(n630), .Z(n639) );
  XOR U732 ( .A(n638), .B(sreg[100]), .Z(n633) );
  XOR U733 ( .A(n639), .B(n633), .Z(c[100]) );
  ANDN U734 ( .B(a[39]), .A(n802), .Z(n641) );
  AND U735 ( .A(a[38]), .B(b[1]), .Z(n643) );
  XNOR U736 ( .A(n643), .B(n642), .Z(n637) );
  XNOR U737 ( .A(n641), .B(n637), .Z(n646) );
  XOR U738 ( .A(n645), .B(sreg[101]), .Z(n640) );
  XOR U739 ( .A(n646), .B(n640), .Z(c[101]) );
  ANDN U740 ( .B(a[40]), .A(n802), .Z(n648) );
  AND U741 ( .A(a[39]), .B(b[1]), .Z(n650) );
  XNOR U742 ( .A(n650), .B(n649), .Z(n644) );
  XNOR U743 ( .A(n648), .B(n644), .Z(n653) );
  XOR U744 ( .A(n652), .B(sreg[102]), .Z(n647) );
  XOR U745 ( .A(n653), .B(n647), .Z(c[102]) );
  ANDN U746 ( .B(a[41]), .A(n802), .Z(n655) );
  AND U747 ( .A(a[40]), .B(b[1]), .Z(n657) );
  XNOR U748 ( .A(n657), .B(n656), .Z(n651) );
  XNOR U749 ( .A(n655), .B(n651), .Z(n660) );
  XOR U750 ( .A(n659), .B(sreg[103]), .Z(n654) );
  XOR U751 ( .A(n660), .B(n654), .Z(c[103]) );
  ANDN U752 ( .B(a[42]), .A(n802), .Z(n662) );
  AND U753 ( .A(a[41]), .B(b[1]), .Z(n664) );
  XNOR U754 ( .A(n664), .B(n663), .Z(n658) );
  XNOR U755 ( .A(n662), .B(n658), .Z(n667) );
  XOR U756 ( .A(n666), .B(sreg[104]), .Z(n661) );
  XOR U757 ( .A(n667), .B(n661), .Z(c[104]) );
  ANDN U758 ( .B(a[43]), .A(n802), .Z(n669) );
  AND U759 ( .A(a[42]), .B(b[1]), .Z(n671) );
  XNOR U760 ( .A(n671), .B(n670), .Z(n665) );
  XNOR U761 ( .A(n669), .B(n665), .Z(n674) );
  XOR U762 ( .A(n673), .B(sreg[105]), .Z(n668) );
  XOR U763 ( .A(n674), .B(n668), .Z(c[105]) );
  ANDN U764 ( .B(a[44]), .A(n802), .Z(n676) );
  AND U765 ( .A(a[43]), .B(b[1]), .Z(n678) );
  XNOR U766 ( .A(n678), .B(n677), .Z(n672) );
  XNOR U767 ( .A(n676), .B(n672), .Z(n681) );
  XOR U768 ( .A(n680), .B(sreg[106]), .Z(n675) );
  XOR U769 ( .A(n681), .B(n675), .Z(c[106]) );
  ANDN U770 ( .B(a[45]), .A(n802), .Z(n683) );
  AND U771 ( .A(a[44]), .B(b[1]), .Z(n685) );
  XNOR U772 ( .A(n685), .B(n684), .Z(n679) );
  XNOR U773 ( .A(n683), .B(n679), .Z(n688) );
  XOR U774 ( .A(n687), .B(sreg[107]), .Z(n682) );
  XOR U775 ( .A(n688), .B(n682), .Z(c[107]) );
  ANDN U776 ( .B(a[46]), .A(n802), .Z(n690) );
  AND U777 ( .A(a[45]), .B(b[1]), .Z(n692) );
  XNOR U778 ( .A(n692), .B(n691), .Z(n686) );
  XNOR U779 ( .A(n690), .B(n686), .Z(n695) );
  XOR U780 ( .A(n694), .B(sreg[108]), .Z(n689) );
  XOR U781 ( .A(n695), .B(n689), .Z(c[108]) );
  ANDN U782 ( .B(a[47]), .A(n802), .Z(n697) );
  AND U783 ( .A(a[46]), .B(b[1]), .Z(n699) );
  XNOR U784 ( .A(n699), .B(n698), .Z(n693) );
  XNOR U785 ( .A(n697), .B(n693), .Z(n702) );
  XOR U786 ( .A(n701), .B(sreg[109]), .Z(n696) );
  XOR U787 ( .A(n702), .B(n696), .Z(c[109]) );
  ANDN U788 ( .B(a[48]), .A(n802), .Z(n704) );
  AND U789 ( .A(a[47]), .B(b[1]), .Z(n706) );
  XNOR U790 ( .A(n706), .B(n705), .Z(n700) );
  XNOR U791 ( .A(n704), .B(n700), .Z(n709) );
  XOR U792 ( .A(n708), .B(sreg[110]), .Z(n703) );
  XOR U793 ( .A(n709), .B(n703), .Z(c[110]) );
  ANDN U794 ( .B(a[49]), .A(n802), .Z(n711) );
  AND U795 ( .A(a[48]), .B(b[1]), .Z(n713) );
  XNOR U796 ( .A(n713), .B(n712), .Z(n707) );
  XNOR U797 ( .A(n711), .B(n707), .Z(n716) );
  XOR U798 ( .A(n715), .B(sreg[111]), .Z(n710) );
  XOR U799 ( .A(n716), .B(n710), .Z(c[111]) );
  ANDN U800 ( .B(a[50]), .A(n802), .Z(n718) );
  AND U801 ( .A(a[49]), .B(b[1]), .Z(n720) );
  XNOR U802 ( .A(n720), .B(n719), .Z(n714) );
  XNOR U803 ( .A(n718), .B(n714), .Z(n723) );
  XOR U804 ( .A(n722), .B(sreg[112]), .Z(n717) );
  XOR U805 ( .A(n723), .B(n717), .Z(c[112]) );
  ANDN U806 ( .B(a[51]), .A(n802), .Z(n725) );
  AND U807 ( .A(a[50]), .B(b[1]), .Z(n727) );
  XNOR U808 ( .A(n727), .B(n726), .Z(n721) );
  XNOR U809 ( .A(n725), .B(n721), .Z(n730) );
  XOR U810 ( .A(n729), .B(sreg[113]), .Z(n724) );
  XOR U811 ( .A(n730), .B(n724), .Z(c[113]) );
  ANDN U812 ( .B(a[52]), .A(n802), .Z(n732) );
  AND U813 ( .A(a[51]), .B(b[1]), .Z(n734) );
  XNOR U814 ( .A(n734), .B(n733), .Z(n728) );
  XNOR U815 ( .A(n732), .B(n728), .Z(n737) );
  XOR U816 ( .A(n736), .B(sreg[114]), .Z(n731) );
  XOR U817 ( .A(n737), .B(n731), .Z(c[114]) );
  ANDN U818 ( .B(a[53]), .A(n802), .Z(n739) );
  AND U819 ( .A(a[52]), .B(b[1]), .Z(n741) );
  XNOR U820 ( .A(n741), .B(n740), .Z(n735) );
  XNOR U821 ( .A(n739), .B(n735), .Z(n744) );
  XOR U822 ( .A(n743), .B(sreg[115]), .Z(n738) );
  XOR U823 ( .A(n744), .B(n738), .Z(c[115]) );
  ANDN U824 ( .B(a[54]), .A(n802), .Z(n746) );
  AND U825 ( .A(a[53]), .B(b[1]), .Z(n748) );
  XNOR U826 ( .A(n748), .B(n747), .Z(n742) );
  XNOR U827 ( .A(n746), .B(n742), .Z(n751) );
  XOR U828 ( .A(n750), .B(sreg[116]), .Z(n745) );
  XOR U829 ( .A(n751), .B(n745), .Z(c[116]) );
  ANDN U830 ( .B(a[55]), .A(n802), .Z(n753) );
  AND U831 ( .A(a[54]), .B(b[1]), .Z(n755) );
  XNOR U832 ( .A(n755), .B(n754), .Z(n749) );
  XNOR U833 ( .A(n753), .B(n749), .Z(n758) );
  XOR U834 ( .A(n757), .B(sreg[117]), .Z(n752) );
  XOR U835 ( .A(n758), .B(n752), .Z(c[117]) );
  ANDN U836 ( .B(a[56]), .A(n802), .Z(n760) );
  AND U837 ( .A(a[55]), .B(b[1]), .Z(n762) );
  XNOR U838 ( .A(n762), .B(n761), .Z(n756) );
  XNOR U839 ( .A(n760), .B(n756), .Z(n765) );
  XOR U840 ( .A(n764), .B(sreg[118]), .Z(n759) );
  XOR U841 ( .A(n765), .B(n759), .Z(c[118]) );
  ANDN U842 ( .B(a[57]), .A(n802), .Z(n767) );
  AND U843 ( .A(a[56]), .B(b[1]), .Z(n769) );
  XNOR U844 ( .A(n769), .B(n768), .Z(n763) );
  XNOR U845 ( .A(n767), .B(n763), .Z(n772) );
  XOR U846 ( .A(n771), .B(sreg[119]), .Z(n766) );
  XOR U847 ( .A(n772), .B(n766), .Z(c[119]) );
  ANDN U848 ( .B(a[58]), .A(n802), .Z(n774) );
  AND U849 ( .A(a[57]), .B(b[1]), .Z(n776) );
  XNOR U850 ( .A(n776), .B(n775), .Z(n770) );
  XNOR U851 ( .A(n774), .B(n770), .Z(n779) );
  XOR U852 ( .A(n778), .B(sreg[120]), .Z(n773) );
  XOR U853 ( .A(n779), .B(n773), .Z(c[120]) );
  ANDN U854 ( .B(a[59]), .A(n802), .Z(n781) );
  AND U855 ( .A(a[58]), .B(b[1]), .Z(n783) );
  XNOR U856 ( .A(n783), .B(n782), .Z(n777) );
  XNOR U857 ( .A(n781), .B(n777), .Z(n786) );
  XOR U858 ( .A(n785), .B(sreg[121]), .Z(n780) );
  XOR U859 ( .A(n786), .B(n780), .Z(c[121]) );
  ANDN U860 ( .B(a[60]), .A(n802), .Z(n788) );
  AND U861 ( .A(a[59]), .B(b[1]), .Z(n790) );
  XNOR U862 ( .A(n790), .B(n789), .Z(n784) );
  XNOR U863 ( .A(n788), .B(n784), .Z(n793) );
  XOR U864 ( .A(n792), .B(sreg[122]), .Z(n787) );
  XOR U865 ( .A(n793), .B(n787), .Z(c[122]) );
  ANDN U866 ( .B(a[61]), .A(n802), .Z(n795) );
  AND U867 ( .A(a[60]), .B(b[1]), .Z(n797) );
  XNOR U868 ( .A(n797), .B(n796), .Z(n791) );
  XNOR U869 ( .A(n795), .B(n791), .Z(n800) );
  XOR U870 ( .A(n799), .B(sreg[123]), .Z(n794) );
  XOR U871 ( .A(n800), .B(n794), .Z(c[123]) );
  AND U872 ( .A(a[61]), .B(b[1]), .Z(n805) );
  AND U873 ( .A(a[62]), .B(b[0]), .Z(n803) );
  XNOR U874 ( .A(n803), .B(n804), .Z(n798) );
  XOR U875 ( .A(n805), .B(n798), .Z(n807) );
  XOR U876 ( .A(n806), .B(sreg[124]), .Z(n801) );
  XNOR U877 ( .A(n807), .B(n801), .Z(c[124]) );
  NANDN U878 ( .A(n364), .B(a[62]), .Z(n812) );
  NANDN U879 ( .A(n802), .B(a[63]), .Z(n811) );
  XOR U880 ( .A(n812), .B(n811), .Z(n813) );
  XNOR U881 ( .A(n813), .B(n814), .Z(n810) );
  XOR U882 ( .A(n809), .B(sreg[125]), .Z(n808) );
  XOR U883 ( .A(n810), .B(n808), .Z(c[125]) );
  AND U884 ( .A(a[63]), .B(b[1]), .Z(n818) );
  OR U885 ( .A(n812), .B(n811), .Z(n816) );
  NANDN U886 ( .A(n814), .B(n813), .Z(n815) );
  AND U887 ( .A(n816), .B(n815), .Z(n819) );
  XNOR U888 ( .A(n820), .B(n819), .Z(n817) );
  XOR U889 ( .A(n818), .B(n817), .Z(c[126]) );
  NANDN U890 ( .A(n818), .B(n817), .Z(n822) );
  NANDN U891 ( .A(n820), .B(n819), .Z(n821) );
  AND U892 ( .A(n822), .B(n821), .Z(c[127]) );
endmodule

