
module mult_N128_CC4 ( clk, rst, a, b, c );
  input [127:0] a;
  input [31:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452;
  wire   [255:0] sreg;

  DFF \sreg_reg[223]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U35 ( .A(n19407), .B(n19408), .Z(n1) );
  NAND U36 ( .A(n19406), .B(n19422), .Z(n2) );
  NAND U37 ( .A(n1), .B(n2), .Z(n19433) );
  NAND U38 ( .A(n18318), .B(n18223), .Z(n3) );
  NANDN U39 ( .A(n18225), .B(n18224), .Z(n4) );
  AND U40 ( .A(n3), .B(n4), .Z(n18338) );
  NAND U41 ( .A(n19018), .B(n19017), .Z(n5) );
  NANDN U42 ( .A(n19016), .B(n19015), .Z(n6) );
  NAND U43 ( .A(n5), .B(n6), .Z(n19079) );
  NAND U44 ( .A(n19420), .B(n19421), .Z(n7) );
  NANDN U45 ( .A(n19422), .B(n19423), .Z(n8) );
  AND U46 ( .A(n7), .B(n8), .Z(n19446) );
  XOR U47 ( .A(n16420), .B(n16419), .Z(n16468) );
  XNOR U48 ( .A(n18134), .B(n18135), .Z(n18137) );
  NAND U49 ( .A(n18341), .B(n18342), .Z(n9) );
  NANDN U50 ( .A(n18344), .B(n18343), .Z(n10) );
  AND U51 ( .A(n9), .B(n10), .Z(n18398) );
  NAND U52 ( .A(n18482), .B(n18445), .Z(n11) );
  NANDN U53 ( .A(n18447), .B(n18446), .Z(n12) );
  AND U54 ( .A(n11), .B(n12), .Z(n18534) );
  NAND U55 ( .A(n18978), .B(n18911), .Z(n13) );
  NANDN U56 ( .A(n18913), .B(n18912), .Z(n14) );
  NAND U57 ( .A(n13), .B(n14), .Z(n19019) );
  NAND U58 ( .A(n1250), .B(n1249), .Z(n15) );
  NAND U59 ( .A(n1247), .B(n1248), .Z(n16) );
  AND U60 ( .A(n15), .B(n16), .Z(n1433) );
  NAND U61 ( .A(n19078), .B(n19079), .Z(n17) );
  NANDN U62 ( .A(n19081), .B(n19080), .Z(n18) );
  NAND U63 ( .A(n17), .B(n18), .Z(n19093) );
  NAND U64 ( .A(n185), .B(n186), .Z(n19) );
  NANDN U65 ( .A(n188), .B(n187), .Z(n20) );
  AND U66 ( .A(n19), .B(n20), .Z(n219) );
  XOR U67 ( .A(n1051), .B(sreg[115]), .Z(n21) );
  NANDN U68 ( .A(n1052), .B(n21), .Z(n22) );
  NAND U69 ( .A(n1051), .B(sreg[115]), .Z(n23) );
  AND U70 ( .A(n22), .B(n23), .Z(n1235) );
  NAND U71 ( .A(n1243), .B(n1244), .Z(n24) );
  NANDN U72 ( .A(n1246), .B(n1245), .Z(n25) );
  AND U73 ( .A(n24), .B(n25), .Z(n1336) );
  XOR U74 ( .A(n796), .B(sreg[112]), .Z(n26) );
  NANDN U75 ( .A(n797), .B(n26), .Z(n27) );
  NAND U76 ( .A(n796), .B(sreg[112]), .Z(n28) );
  AND U77 ( .A(n27), .B(n28), .Z(n878) );
  NAND U78 ( .A(n19437), .B(n19438), .Z(n29) );
  NANDN U79 ( .A(n19440), .B(n19439), .Z(n30) );
  NAND U80 ( .A(n29), .B(n30), .Z(n19452) );
  NANDN U81 ( .A(b[0]), .B(a[127]), .Z(n31) );
  NAND U82 ( .A(b[1]), .B(n31), .Z(n16893) );
  NAND U83 ( .A(n3573), .B(n3572), .Z(n32) );
  NANDN U84 ( .A(n3571), .B(n3570), .Z(n33) );
  AND U85 ( .A(n32), .B(n33), .Z(n3768) );
  NAND U86 ( .A(n4316), .B(n4315), .Z(n34) );
  NANDN U87 ( .A(n4314), .B(n4313), .Z(n35) );
  AND U88 ( .A(n34), .B(n35), .Z(n4517) );
  NAND U89 ( .A(n4916), .B(n4915), .Z(n36) );
  NANDN U90 ( .A(n4914), .B(n4913), .Z(n37) );
  AND U91 ( .A(n36), .B(n37), .Z(n5111) );
  NAND U92 ( .A(n5212), .B(n5211), .Z(n38) );
  NANDN U93 ( .A(n5210), .B(n5209), .Z(n39) );
  AND U94 ( .A(n38), .B(n39), .Z(n5405) );
  NAND U95 ( .A(n5347), .B(n5346), .Z(n40) );
  NANDN U96 ( .A(n5345), .B(n5344), .Z(n41) );
  AND U97 ( .A(n40), .B(n41), .Z(n5554) );
  NAND U98 ( .A(n6251), .B(n6250), .Z(n42) );
  NANDN U99 ( .A(n6249), .B(n6248), .Z(n43) );
  AND U100 ( .A(n42), .B(n43), .Z(n6440) );
  NAND U101 ( .A(n7882), .B(n7881), .Z(n44) );
  NANDN U102 ( .A(n7880), .B(n7879), .Z(n45) );
  AND U103 ( .A(n44), .B(n45), .Z(n8083) );
  NAND U104 ( .A(n9376), .B(n9375), .Z(n46) );
  NANDN U105 ( .A(n9374), .B(n9373), .Z(n47) );
  AND U106 ( .A(n46), .B(n47), .Z(n9563) );
  NAND U107 ( .A(n9505), .B(n9504), .Z(n48) );
  NANDN U108 ( .A(n9503), .B(n9502), .Z(n49) );
  AND U109 ( .A(n48), .B(n49), .Z(n9716) );
  NAND U110 ( .A(n9658), .B(n9657), .Z(n50) );
  NANDN U111 ( .A(n9656), .B(n9655), .Z(n51) );
  AND U112 ( .A(n50), .B(n51), .Z(n9865) );
  NAND U113 ( .A(n9966), .B(n9965), .Z(n52) );
  NANDN U114 ( .A(n9964), .B(n9963), .Z(n53) );
  AND U115 ( .A(n52), .B(n53), .Z(n10153) );
  NAND U116 ( .A(n10095), .B(n10094), .Z(n54) );
  NANDN U117 ( .A(n10093), .B(n10092), .Z(n55) );
  AND U118 ( .A(n54), .B(n55), .Z(n10306) );
  NAND U119 ( .A(n10248), .B(n10247), .Z(n56) );
  NANDN U120 ( .A(n10246), .B(n10245), .Z(n57) );
  AND U121 ( .A(n56), .B(n57), .Z(n10455) );
  NAND U122 ( .A(n10556), .B(n10555), .Z(n58) );
  NANDN U123 ( .A(n10554), .B(n10553), .Z(n59) );
  AND U124 ( .A(n58), .B(n59), .Z(n10751) );
  NAND U125 ( .A(n12187), .B(n12186), .Z(n60) );
  NANDN U126 ( .A(n12185), .B(n12184), .Z(n61) );
  AND U127 ( .A(n60), .B(n61), .Z(n12380) );
  NAND U128 ( .A(n12322), .B(n12321), .Z(n62) );
  NANDN U129 ( .A(n12320), .B(n12319), .Z(n63) );
  AND U130 ( .A(n62), .B(n63), .Z(n12535) );
  NAND U131 ( .A(n12785), .B(n12784), .Z(n64) );
  NANDN U132 ( .A(n12783), .B(n12782), .Z(n65) );
  AND U133 ( .A(n64), .B(n65), .Z(n12974) );
  NAND U134 ( .A(n13820), .B(n13819), .Z(n66) );
  NANDN U135 ( .A(n13818), .B(n13817), .Z(n67) );
  AND U136 ( .A(n66), .B(n67), .Z(n14015) );
  NAND U137 ( .A(n14122), .B(n14121), .Z(n68) );
  NANDN U138 ( .A(n14120), .B(n14119), .Z(n69) );
  AND U139 ( .A(n68), .B(n69), .Z(n14315) );
  NAND U140 ( .A(n14257), .B(n14256), .Z(n70) );
  NANDN U141 ( .A(n14255), .B(n14254), .Z(n71) );
  AND U142 ( .A(n70), .B(n71), .Z(n14464) );
  NAND U143 ( .A(n14708), .B(n14707), .Z(n72) );
  NANDN U144 ( .A(n14706), .B(n14705), .Z(n73) );
  AND U145 ( .A(n72), .B(n73), .Z(n14903) );
  XOR U146 ( .A(n17081), .B(n17080), .Z(n17093) );
  NAND U147 ( .A(n1628), .B(n1627), .Z(n74) );
  NANDN U148 ( .A(n1626), .B(n1625), .Z(n75) );
  AND U149 ( .A(n74), .B(n75), .Z(n1783) );
  NAND U150 ( .A(n16351), .B(n16350), .Z(n76) );
  NANDN U151 ( .A(n16349), .B(n16348), .Z(n77) );
  AND U152 ( .A(n76), .B(n77), .Z(n16534) );
  NAND U153 ( .A(n18135), .B(n17989), .Z(n78) );
  NANDN U154 ( .A(n17991), .B(n17990), .Z(n79) );
  NAND U155 ( .A(n78), .B(n79), .Z(n18152) );
  NAND U156 ( .A(n18079), .B(n18078), .Z(n80) );
  NANDN U157 ( .A(n18077), .B(n18076), .Z(n81) );
  AND U158 ( .A(n80), .B(n81), .Z(n18186) );
  NAND U159 ( .A(n18494), .B(n18495), .Z(n82) );
  NANDN U160 ( .A(n18497), .B(n18496), .Z(n83) );
  NAND U161 ( .A(n82), .B(n83), .Z(n18634) );
  NAND U162 ( .A(n709), .B(n708), .Z(n84) );
  NANDN U163 ( .A(n707), .B(n706), .Z(n85) );
  NAND U164 ( .A(n84), .B(n85), .Z(n727) );
  NAND U165 ( .A(n1574), .B(n1573), .Z(n86) );
  NANDN U166 ( .A(n1572), .B(n1571), .Z(n87) );
  AND U167 ( .A(n86), .B(n87), .Z(n1691) );
  NAND U168 ( .A(n16689), .B(n16688), .Z(n88) );
  NAND U169 ( .A(n16687), .B(n16686), .Z(n89) );
  AND U170 ( .A(n88), .B(n89), .Z(n16719) );
  NAND U171 ( .A(n18362), .B(n18361), .Z(n90) );
  NAND U172 ( .A(n18359), .B(n18360), .Z(n91) );
  AND U173 ( .A(n90), .B(n91), .Z(n18455) );
  NAND U174 ( .A(n18395), .B(n18396), .Z(n92) );
  NANDN U175 ( .A(n18398), .B(n18397), .Z(n93) );
  NAND U176 ( .A(n92), .B(n93), .Z(n18469) );
  NAND U177 ( .A(n18979), .B(n18980), .Z(n94) );
  NANDN U178 ( .A(n18978), .B(n18977), .Z(n95) );
  AND U179 ( .A(n94), .B(n95), .Z(n19037) );
  NAND U180 ( .A(n19105), .B(n19104), .Z(n96) );
  NANDN U181 ( .A(n19103), .B(n19102), .Z(n97) );
  AND U182 ( .A(n96), .B(n97), .Z(n19156) );
  NAND U183 ( .A(n1329), .B(n1330), .Z(n98) );
  NANDN U184 ( .A(n1332), .B(n1331), .Z(n99) );
  AND U185 ( .A(n98), .B(n99), .Z(n1333) );
  NAND U186 ( .A(n19033), .B(n19034), .Z(n100) );
  NANDN U187 ( .A(n19036), .B(n19035), .Z(n101) );
  AND U188 ( .A(n100), .B(n101), .Z(n19085) );
  XOR U189 ( .A(n175), .B(n173), .Z(n102) );
  NANDN U190 ( .A(n174), .B(n102), .Z(n103) );
  NAND U191 ( .A(n175), .B(n173), .Z(n104) );
  AND U192 ( .A(n103), .B(n104), .Z(n188) );
  NAND U193 ( .A(n1241), .B(n1242), .Z(n105) );
  XOR U194 ( .A(n1241), .B(n1242), .Z(n106) );
  NAND U195 ( .A(n106), .B(sreg[117]), .Z(n107) );
  NAND U196 ( .A(n105), .B(n107), .Z(n1438) );
  NAND U197 ( .A(sreg[125]), .B(n2177), .Z(n108) );
  XOR U198 ( .A(sreg[125]), .B(n2177), .Z(n109) );
  NANDN U199 ( .A(n2176), .B(n109), .Z(n110) );
  NAND U200 ( .A(n108), .B(n110), .Z(n2310) );
  XOR U201 ( .A(n960), .B(sreg[114]), .Z(n111) );
  NANDN U202 ( .A(n961), .B(n111), .Z(n112) );
  NAND U203 ( .A(n960), .B(sreg[114]), .Z(n113) );
  AND U204 ( .A(n112), .B(n113), .Z(n1052) );
  XOR U205 ( .A(n1787), .B(sreg[122]), .Z(n114) );
  NANDN U206 ( .A(n1788), .B(n114), .Z(n115) );
  NAND U207 ( .A(n1787), .B(sreg[122]), .Z(n116) );
  AND U208 ( .A(n115), .B(n116), .Z(n1913) );
  XOR U209 ( .A(n2602), .B(sreg[128]), .Z(n117) );
  NANDN U210 ( .A(n2603), .B(n117), .Z(n118) );
  NAND U211 ( .A(n2602), .B(sreg[128]), .Z(n119) );
  AND U212 ( .A(n118), .B(n119), .Z(n2895) );
  NAND U213 ( .A(sreg[131]), .B(n3049), .Z(n120) );
  XOR U214 ( .A(sreg[131]), .B(n3049), .Z(n121) );
  NANDN U215 ( .A(n3048), .B(n121), .Z(n122) );
  NAND U216 ( .A(n120), .B(n122), .Z(n3340) );
  XNOR U217 ( .A(a[127]), .B(a[126]), .Z(n123) );
  XNOR U218 ( .A(n19443), .B(n123), .Z(n124) );
  AND U219 ( .A(n124), .B(b[31]), .Z(n125) );
  NANDN U220 ( .A(n19446), .B(n19447), .Z(n126) );
  NANDN U221 ( .A(n19444), .B(n19445), .Z(n127) );
  AND U222 ( .A(n126), .B(n127), .Z(n128) );
  NOR U223 ( .A(n19452), .B(n19451), .Z(n129) );
  NANDN U224 ( .A(n19448), .B(n19451), .Z(n130) );
  OR U225 ( .A(n129), .B(n19449), .Z(n131) );
  NAND U226 ( .A(n130), .B(n131), .Z(n132) );
  OR U227 ( .A(n19449), .B(n130), .Z(n133) );
  NANDN U228 ( .A(n19450), .B(n133), .Z(n134) );
  NAND U229 ( .A(n132), .B(n134), .Z(n135) );
  XNOR U230 ( .A(n125), .B(n128), .Z(n136) );
  XNOR U231 ( .A(n135), .B(n136), .Z(c[255]) );
  AND U232 ( .A(b[0]), .B(a[0]), .Z(n138) );
  XOR U233 ( .A(n138), .B(sreg[96]), .Z(c[96]) );
  AND U234 ( .A(b[0]), .B(a[1]), .Z(n145) );
  NAND U235 ( .A(a[0]), .B(b[1]), .Z(n137) );
  XOR U236 ( .A(n145), .B(n137), .Z(n139) );
  XNOR U237 ( .A(sreg[97]), .B(n139), .Z(n141) );
  AND U238 ( .A(n138), .B(sreg[96]), .Z(n140) );
  XOR U239 ( .A(n141), .B(n140), .Z(c[97]) );
  NANDN U240 ( .A(n139), .B(sreg[97]), .Z(n143) );
  NAND U241 ( .A(n141), .B(n140), .Z(n142) );
  AND U242 ( .A(n143), .B(n142), .Z(n163) );
  XNOR U243 ( .A(n163), .B(sreg[98]), .Z(n165) );
  NAND U244 ( .A(a[0]), .B(b[2]), .Z(n144) );
  XNOR U245 ( .A(b[1]), .B(n144), .Z(n147) );
  NANDN U246 ( .A(a[0]), .B(n145), .Z(n146) );
  NAND U247 ( .A(n147), .B(n146), .Z(n152) );
  NAND U248 ( .A(b[0]), .B(a[2]), .Z(n148) );
  XNOR U249 ( .A(b[1]), .B(n148), .Z(n150) );
  NANDN U250 ( .A(b[0]), .B(a[1]), .Z(n149) );
  NAND U251 ( .A(n150), .B(n149), .Z(n151) );
  XOR U252 ( .A(n152), .B(n151), .Z(n164) );
  XOR U253 ( .A(n165), .B(n164), .Z(c[98]) );
  NOR U254 ( .A(n152), .B(n151), .Z(n175) );
  XOR U255 ( .A(b[3]), .B(b[2]), .Z(n176) );
  XOR U256 ( .A(b[3]), .B(a[0]), .Z(n153) );
  NAND U257 ( .A(n176), .B(n153), .Z(n154) );
  XOR U258 ( .A(b[1]), .B(b[2]), .Z(n2512) );
  OR U259 ( .A(n154), .B(n2512), .Z(n156) );
  XOR U260 ( .A(b[3]), .B(a[1]), .Z(n177) );
  NAND U261 ( .A(n2512), .B(n177), .Z(n155) );
  AND U262 ( .A(n156), .B(n155), .Z(n184) );
  NAND U263 ( .A(b[0]), .B(a[3]), .Z(n157) );
  XNOR U264 ( .A(b[1]), .B(n157), .Z(n159) );
  NANDN U265 ( .A(b[0]), .B(a[2]), .Z(n158) );
  NAND U266 ( .A(n159), .B(n158), .Z(n183) );
  XNOR U267 ( .A(n184), .B(n183), .Z(n174) );
  NAND U268 ( .A(b[1]), .B(b[2]), .Z(n160) );
  AND U269 ( .A(b[3]), .B(n160), .Z(n17335) );
  IV U270 ( .A(n2512), .Z(n17068) );
  NANDN U271 ( .A(n17068), .B(a[0]), .Z(n161) );
  AND U272 ( .A(n17335), .B(n161), .Z(n173) );
  XOR U273 ( .A(n174), .B(n173), .Z(n162) );
  XOR U274 ( .A(n175), .B(n162), .Z(n168) );
  XNOR U275 ( .A(sreg[99]), .B(n168), .Z(n170) );
  NANDN U276 ( .A(n163), .B(sreg[98]), .Z(n167) );
  NAND U277 ( .A(n165), .B(n164), .Z(n166) );
  NAND U278 ( .A(n167), .B(n166), .Z(n169) );
  XOR U279 ( .A(n170), .B(n169), .Z(c[99]) );
  NANDN U280 ( .A(n168), .B(sreg[99]), .Z(n172) );
  NAND U281 ( .A(n170), .B(n169), .Z(n171) );
  AND U282 ( .A(n172), .B(n171), .Z(n206) );
  XNOR U283 ( .A(n206), .B(sreg[100]), .Z(n208) );
  ANDN U284 ( .B(n176), .A(n2512), .Z(n2664) );
  IV U285 ( .A(n2664), .Z(n17067) );
  NANDN U286 ( .A(n17067), .B(n177), .Z(n179) );
  XOR U287 ( .A(b[3]), .B(a[2]), .Z(n189) );
  NANDN U288 ( .A(n17068), .B(n189), .Z(n178) );
  AND U289 ( .A(n179), .B(n178), .Z(n203) );
  XOR U290 ( .A(b[4]), .B(b[3]), .Z(n17391) );
  IV U291 ( .A(n17391), .Z(n17223) );
  ANDN U292 ( .B(a[0]), .A(n17223), .Z(n200) );
  NAND U293 ( .A(b[0]), .B(a[4]), .Z(n180) );
  XNOR U294 ( .A(b[1]), .B(n180), .Z(n182) );
  NANDN U295 ( .A(b[0]), .B(a[3]), .Z(n181) );
  NAND U296 ( .A(n182), .B(n181), .Z(n201) );
  XNOR U297 ( .A(n200), .B(n201), .Z(n202) );
  XNOR U298 ( .A(n203), .B(n202), .Z(n186) );
  NOR U299 ( .A(n184), .B(n183), .Z(n185) );
  XOR U300 ( .A(n186), .B(n185), .Z(n187) );
  XNOR U301 ( .A(n188), .B(n187), .Z(n207) );
  XOR U302 ( .A(n208), .B(n207), .Z(c[100]) );
  NANDN U303 ( .A(n17067), .B(n189), .Z(n191) );
  XOR U304 ( .A(b[3]), .B(a[3]), .Z(n228) );
  NANDN U305 ( .A(n17068), .B(n228), .Z(n190) );
  AND U306 ( .A(n191), .B(n190), .Z(n235) );
  NAND U307 ( .A(b[3]), .B(b[4]), .Z(n192) );
  AND U308 ( .A(b[5]), .B(n192), .Z(n17658) );
  ANDN U309 ( .B(n17658), .A(n200), .Z(n234) );
  XNOR U310 ( .A(n235), .B(n234), .Z(n237) );
  NAND U311 ( .A(b[0]), .B(a[5]), .Z(n193) );
  XNOR U312 ( .A(b[1]), .B(n193), .Z(n195) );
  NANDN U313 ( .A(b[0]), .B(a[4]), .Z(n194) );
  NAND U314 ( .A(n195), .B(n194), .Z(n226) );
  XOR U315 ( .A(b[5]), .B(b[4]), .Z(n222) );
  XOR U316 ( .A(b[5]), .B(a[0]), .Z(n196) );
  NAND U317 ( .A(n222), .B(n196), .Z(n197) );
  OR U318 ( .A(n197), .B(n17391), .Z(n199) );
  XOR U319 ( .A(b[5]), .B(a[1]), .Z(n223) );
  NAND U320 ( .A(n17391), .B(n223), .Z(n198) );
  NAND U321 ( .A(n199), .B(n198), .Z(n227) );
  XNOR U322 ( .A(n226), .B(n227), .Z(n236) );
  XOR U323 ( .A(n237), .B(n236), .Z(n217) );
  NANDN U324 ( .A(n201), .B(n200), .Z(n205) );
  NANDN U325 ( .A(n203), .B(n202), .Z(n204) );
  AND U326 ( .A(n205), .B(n204), .Z(n216) );
  XNOR U327 ( .A(n217), .B(n216), .Z(n218) );
  XOR U328 ( .A(n219), .B(n218), .Z(n211) );
  XNOR U329 ( .A(n211), .B(sreg[101]), .Z(n213) );
  NANDN U330 ( .A(n206), .B(sreg[100]), .Z(n210) );
  NAND U331 ( .A(n208), .B(n207), .Z(n209) );
  NAND U332 ( .A(n210), .B(n209), .Z(n212) );
  XOR U333 ( .A(n213), .B(n212), .Z(c[101]) );
  NANDN U334 ( .A(n211), .B(sreg[101]), .Z(n215) );
  NAND U335 ( .A(n213), .B(n212), .Z(n214) );
  AND U336 ( .A(n215), .B(n214), .Z(n272) );
  XNOR U337 ( .A(n272), .B(sreg[102]), .Z(n274) );
  NANDN U338 ( .A(n217), .B(n216), .Z(n221) );
  NAND U339 ( .A(n219), .B(n218), .Z(n220) );
  AND U340 ( .A(n221), .B(n220), .Z(n242) );
  ANDN U341 ( .B(n222), .A(n17391), .Z(n17390) );
  IV U342 ( .A(n17390), .Z(n17072) );
  NANDN U343 ( .A(n17072), .B(n223), .Z(n225) );
  XOR U344 ( .A(b[5]), .B(a[2]), .Z(n250) );
  NANDN U345 ( .A(n17223), .B(n250), .Z(n224) );
  AND U346 ( .A(n225), .B(n224), .Z(n267) );
  ANDN U347 ( .B(n227), .A(n226), .Z(n266) );
  XNOR U348 ( .A(n267), .B(n266), .Z(n269) );
  NANDN U349 ( .A(n17067), .B(n228), .Z(n230) );
  XOR U350 ( .A(b[3]), .B(a[4]), .Z(n257) );
  NANDN U351 ( .A(n17068), .B(n257), .Z(n229) );
  AND U352 ( .A(n230), .B(n229), .Z(n263) );
  XOR U353 ( .A(b[6]), .B(b[5]), .Z(n17624) );
  IV U354 ( .A(n17624), .Z(n17522) );
  ANDN U355 ( .B(a[0]), .A(n17522), .Z(n260) );
  NAND U356 ( .A(b[0]), .B(a[6]), .Z(n231) );
  XNOR U357 ( .A(b[1]), .B(n231), .Z(n233) );
  NANDN U358 ( .A(b[0]), .B(a[5]), .Z(n232) );
  NAND U359 ( .A(n233), .B(n232), .Z(n261) );
  XNOR U360 ( .A(n260), .B(n261), .Z(n262) );
  XNOR U361 ( .A(n263), .B(n262), .Z(n268) );
  XOR U362 ( .A(n269), .B(n268), .Z(n241) );
  NANDN U363 ( .A(n235), .B(n234), .Z(n239) );
  NAND U364 ( .A(n237), .B(n236), .Z(n238) );
  AND U365 ( .A(n239), .B(n238), .Z(n240) );
  XOR U366 ( .A(n241), .B(n240), .Z(n243) );
  XNOR U367 ( .A(n242), .B(n243), .Z(n273) );
  XOR U368 ( .A(n274), .B(n273), .Z(c[102]) );
  NANDN U369 ( .A(n241), .B(n240), .Z(n245) );
  OR U370 ( .A(n243), .B(n242), .Z(n244) );
  AND U371 ( .A(n245), .B(n244), .Z(n284) );
  XOR U372 ( .A(b[7]), .B(b[6]), .Z(n300) );
  XOR U373 ( .A(b[7]), .B(a[0]), .Z(n246) );
  NAND U374 ( .A(n300), .B(n246), .Z(n247) );
  OR U375 ( .A(n247), .B(n17624), .Z(n249) );
  XOR U376 ( .A(b[7]), .B(a[1]), .Z(n301) );
  NAND U377 ( .A(n17624), .B(n301), .Z(n248) );
  AND U378 ( .A(n249), .B(n248), .Z(n308) );
  NANDN U379 ( .A(n17072), .B(n250), .Z(n252) );
  XOR U380 ( .A(b[5]), .B(a[3]), .Z(n312) );
  NANDN U381 ( .A(n17223), .B(n312), .Z(n251) );
  AND U382 ( .A(n252), .B(n251), .Z(n307) );
  XOR U383 ( .A(n308), .B(n307), .Z(n297) );
  NAND U384 ( .A(b[5]), .B(b[6]), .Z(n253) );
  NAND U385 ( .A(b[7]), .B(n253), .Z(n17746) );
  NOR U386 ( .A(n17746), .B(n260), .Z(n295) );
  NAND U387 ( .A(b[0]), .B(a[7]), .Z(n254) );
  XNOR U388 ( .A(b[1]), .B(n254), .Z(n256) );
  NANDN U389 ( .A(b[0]), .B(a[6]), .Z(n255) );
  NAND U390 ( .A(n256), .B(n255), .Z(n294) );
  XNOR U391 ( .A(n295), .B(n294), .Z(n296) );
  XNOR U392 ( .A(n297), .B(n296), .Z(n288) );
  NAND U393 ( .A(n2664), .B(n257), .Z(n259) );
  XNOR U394 ( .A(b[3]), .B(a[5]), .Z(n304) );
  NANDN U395 ( .A(n304), .B(n2512), .Z(n258) );
  NAND U396 ( .A(n259), .B(n258), .Z(n289) );
  XNOR U397 ( .A(n288), .B(n289), .Z(n290) );
  NANDN U398 ( .A(n261), .B(n260), .Z(n265) );
  NANDN U399 ( .A(n263), .B(n262), .Z(n264) );
  NAND U400 ( .A(n265), .B(n264), .Z(n291) );
  XNOR U401 ( .A(n290), .B(n291), .Z(n282) );
  NANDN U402 ( .A(n267), .B(n266), .Z(n271) );
  NAND U403 ( .A(n269), .B(n268), .Z(n270) );
  NAND U404 ( .A(n271), .B(n270), .Z(n283) );
  XOR U405 ( .A(n282), .B(n283), .Z(n285) );
  XOR U406 ( .A(n284), .B(n285), .Z(n277) );
  XNOR U407 ( .A(n277), .B(sreg[103]), .Z(n279) );
  NANDN U408 ( .A(n272), .B(sreg[102]), .Z(n276) );
  NAND U409 ( .A(n274), .B(n273), .Z(n275) );
  NAND U410 ( .A(n276), .B(n275), .Z(n278) );
  XOR U411 ( .A(n279), .B(n278), .Z(c[103]) );
  NANDN U412 ( .A(n277), .B(sreg[103]), .Z(n281) );
  NAND U413 ( .A(n279), .B(n278), .Z(n280) );
  AND U414 ( .A(n281), .B(n280), .Z(n358) );
  XNOR U415 ( .A(n358), .B(sreg[104]), .Z(n360) );
  NANDN U416 ( .A(n283), .B(n282), .Z(n287) );
  OR U417 ( .A(n285), .B(n284), .Z(n286) );
  AND U418 ( .A(n287), .B(n286), .Z(n354) );
  NANDN U419 ( .A(n289), .B(n288), .Z(n293) );
  NANDN U420 ( .A(n291), .B(n290), .Z(n292) );
  AND U421 ( .A(n293), .B(n292), .Z(n353) );
  NANDN U422 ( .A(n295), .B(n294), .Z(n299) );
  NANDN U423 ( .A(n297), .B(n296), .Z(n298) );
  AND U424 ( .A(n299), .B(n298), .Z(n318) );
  ANDN U425 ( .B(n300), .A(n17624), .Z(n17623) );
  IV U426 ( .A(n17623), .Z(n17362) );
  NANDN U427 ( .A(n17362), .B(n301), .Z(n303) );
  XOR U428 ( .A(b[7]), .B(a[2]), .Z(n332) );
  NANDN U429 ( .A(n17522), .B(n332), .Z(n302) );
  AND U430 ( .A(n303), .B(n302), .Z(n322) );
  NANDN U431 ( .A(n304), .B(n2664), .Z(n306) );
  XOR U432 ( .A(b[3]), .B(a[6]), .Z(n349) );
  NANDN U433 ( .A(n17068), .B(n349), .Z(n305) );
  NAND U434 ( .A(n306), .B(n305), .Z(n321) );
  XNOR U435 ( .A(n322), .B(n321), .Z(n324) );
  NOR U436 ( .A(n308), .B(n307), .Z(n323) );
  XOR U437 ( .A(n324), .B(n323), .Z(n316) );
  NAND U438 ( .A(b[0]), .B(a[8]), .Z(n309) );
  XNOR U439 ( .A(b[1]), .B(n309), .Z(n311) );
  NANDN U440 ( .A(b[0]), .B(a[7]), .Z(n310) );
  NAND U441 ( .A(n311), .B(n310), .Z(n329) );
  XOR U442 ( .A(b[7]), .B(b[8]), .Z(n17879) );
  IV U443 ( .A(n17879), .Z(n17739) );
  ANDN U444 ( .B(a[0]), .A(n17739), .Z(n342) );
  NANDN U445 ( .A(n17072), .B(n312), .Z(n314) );
  XOR U446 ( .A(b[5]), .B(a[4]), .Z(n343) );
  NANDN U447 ( .A(n17223), .B(n343), .Z(n313) );
  AND U448 ( .A(n314), .B(n313), .Z(n327) );
  XOR U449 ( .A(n342), .B(n327), .Z(n328) );
  XNOR U450 ( .A(n329), .B(n328), .Z(n315) );
  XNOR U451 ( .A(n316), .B(n315), .Z(n317) );
  XNOR U452 ( .A(n318), .B(n317), .Z(n352) );
  XOR U453 ( .A(n353), .B(n352), .Z(n355) );
  XNOR U454 ( .A(n354), .B(n355), .Z(n359) );
  XOR U455 ( .A(n360), .B(n359), .Z(c[104]) );
  NANDN U456 ( .A(n316), .B(n315), .Z(n320) );
  NANDN U457 ( .A(n318), .B(n317), .Z(n319) );
  AND U458 ( .A(n320), .B(n319), .Z(n368) );
  NANDN U459 ( .A(n322), .B(n321), .Z(n326) );
  NAND U460 ( .A(n324), .B(n323), .Z(n325) );
  AND U461 ( .A(n326), .B(n325), .Z(n407) );
  NANDN U462 ( .A(n327), .B(n342), .Z(n331) );
  OR U463 ( .A(n329), .B(n328), .Z(n330) );
  AND U464 ( .A(n331), .B(n330), .Z(n405) );
  NANDN U465 ( .A(n17362), .B(n332), .Z(n334) );
  XOR U466 ( .A(b[7]), .B(a[3]), .Z(n389) );
  NANDN U467 ( .A(n17522), .B(n389), .Z(n333) );
  AND U468 ( .A(n334), .B(n333), .Z(n399) );
  XOR U469 ( .A(b[9]), .B(a[1]), .Z(n396) );
  NANDN U470 ( .A(n17739), .B(n396), .Z(n341) );
  ANDN U471 ( .B(b[8]), .A(b[9]), .Z(n335) );
  NAND U472 ( .A(n335), .B(a[0]), .Z(n338) );
  NAND U473 ( .A(b[7]), .B(b[8]), .Z(n336) );
  NAND U474 ( .A(b[9]), .B(n336), .Z(n18134) );
  OR U475 ( .A(a[0]), .B(n18134), .Z(n337) );
  NAND U476 ( .A(n338), .B(n337), .Z(n339) );
  NAND U477 ( .A(n17739), .B(n339), .Z(n340) );
  NAND U478 ( .A(n341), .B(n340), .Z(n400) );
  XOR U479 ( .A(n399), .B(n400), .Z(n376) );
  NOR U480 ( .A(n18134), .B(n342), .Z(n375) );
  NANDN U481 ( .A(n17072), .B(n343), .Z(n345) );
  XOR U482 ( .A(b[5]), .B(a[5]), .Z(n392) );
  NANDN U483 ( .A(n17223), .B(n392), .Z(n344) );
  AND U484 ( .A(n345), .B(n344), .Z(n374) );
  XOR U485 ( .A(n375), .B(n374), .Z(n377) );
  XOR U486 ( .A(n376), .B(n377), .Z(n383) );
  NAND U487 ( .A(b[0]), .B(a[9]), .Z(n346) );
  XNOR U488 ( .A(b[1]), .B(n346), .Z(n348) );
  NANDN U489 ( .A(b[0]), .B(a[8]), .Z(n347) );
  NAND U490 ( .A(n348), .B(n347), .Z(n381) );
  NANDN U491 ( .A(n17067), .B(n349), .Z(n351) );
  XOR U492 ( .A(b[3]), .B(a[7]), .Z(n401) );
  NANDN U493 ( .A(n17068), .B(n401), .Z(n350) );
  NAND U494 ( .A(n351), .B(n350), .Z(n380) );
  XNOR U495 ( .A(n381), .B(n380), .Z(n382) );
  XOR U496 ( .A(n383), .B(n382), .Z(n404) );
  XNOR U497 ( .A(n405), .B(n404), .Z(n406) );
  XOR U498 ( .A(n407), .B(n406), .Z(n369) );
  XNOR U499 ( .A(n368), .B(n369), .Z(n370) );
  NANDN U500 ( .A(n353), .B(n352), .Z(n357) );
  OR U501 ( .A(n355), .B(n354), .Z(n356) );
  NAND U502 ( .A(n357), .B(n356), .Z(n371) );
  XOR U503 ( .A(n370), .B(n371), .Z(n363) );
  XNOR U504 ( .A(sreg[105]), .B(n363), .Z(n365) );
  NANDN U505 ( .A(n358), .B(sreg[104]), .Z(n362) );
  NAND U506 ( .A(n360), .B(n359), .Z(n361) );
  NAND U507 ( .A(n362), .B(n361), .Z(n364) );
  XOR U508 ( .A(n365), .B(n364), .Z(c[105]) );
  NANDN U509 ( .A(n363), .B(sreg[105]), .Z(n367) );
  NAND U510 ( .A(n365), .B(n364), .Z(n366) );
  AND U511 ( .A(n367), .B(n366), .Z(n410) );
  XNOR U512 ( .A(n410), .B(sreg[106]), .Z(n412) );
  NANDN U513 ( .A(n369), .B(n368), .Z(n373) );
  NANDN U514 ( .A(n371), .B(n370), .Z(n372) );
  AND U515 ( .A(n373), .B(n372), .Z(n418) );
  NANDN U516 ( .A(n375), .B(n374), .Z(n379) );
  NANDN U517 ( .A(n377), .B(n376), .Z(n378) );
  AND U518 ( .A(n379), .B(n378), .Z(n422) );
  NANDN U519 ( .A(n381), .B(n380), .Z(n385) );
  NAND U520 ( .A(n383), .B(n382), .Z(n384) );
  AND U521 ( .A(n385), .B(n384), .Z(n421) );
  XNOR U522 ( .A(n422), .B(n421), .Z(n423) );
  NAND U523 ( .A(b[0]), .B(a[10]), .Z(n386) );
  XNOR U524 ( .A(b[1]), .B(n386), .Z(n388) );
  NANDN U525 ( .A(b[0]), .B(a[9]), .Z(n387) );
  NAND U526 ( .A(n388), .B(n387), .Z(n429) );
  XOR U527 ( .A(b[10]), .B(b[9]), .Z(n18085) );
  IV U528 ( .A(n18085), .Z(n18025) );
  ANDN U529 ( .B(a[0]), .A(n18025), .Z(n452) );
  NANDN U530 ( .A(n17362), .B(n389), .Z(n391) );
  XOR U531 ( .A(b[7]), .B(a[4]), .Z(n453) );
  NANDN U532 ( .A(n17522), .B(n453), .Z(n390) );
  AND U533 ( .A(n391), .B(n390), .Z(n427) );
  XOR U534 ( .A(n452), .B(n427), .Z(n428) );
  XOR U535 ( .A(n429), .B(n428), .Z(n462) );
  NANDN U536 ( .A(n17072), .B(n392), .Z(n394) );
  XOR U537 ( .A(b[5]), .B(a[6]), .Z(n448) );
  NANDN U538 ( .A(n17223), .B(n448), .Z(n393) );
  AND U539 ( .A(n394), .B(n393), .Z(n433) );
  XOR U540 ( .A(b[8]), .B(b[9]), .Z(n395) );
  ANDN U541 ( .B(n395), .A(n17879), .Z(n17881) );
  IV U542 ( .A(n17881), .Z(n17613) );
  NANDN U543 ( .A(n17613), .B(n396), .Z(n398) );
  XOR U544 ( .A(b[9]), .B(a[2]), .Z(n438) );
  NANDN U545 ( .A(n17739), .B(n438), .Z(n397) );
  NAND U546 ( .A(n398), .B(n397), .Z(n432) );
  XNOR U547 ( .A(n433), .B(n432), .Z(n435) );
  ANDN U548 ( .B(n400), .A(n399), .Z(n434) );
  XOR U549 ( .A(n435), .B(n434), .Z(n460) );
  NAND U550 ( .A(n2664), .B(n401), .Z(n403) );
  XNOR U551 ( .A(b[3]), .B(a[8]), .Z(n456) );
  NANDN U552 ( .A(n456), .B(n2512), .Z(n402) );
  AND U553 ( .A(n403), .B(n402), .Z(n459) );
  XNOR U554 ( .A(n460), .B(n459), .Z(n461) );
  XOR U555 ( .A(n462), .B(n461), .Z(n424) );
  XNOR U556 ( .A(n423), .B(n424), .Z(n415) );
  NANDN U557 ( .A(n405), .B(n404), .Z(n409) );
  NANDN U558 ( .A(n407), .B(n406), .Z(n408) );
  NAND U559 ( .A(n409), .B(n408), .Z(n416) );
  XNOR U560 ( .A(n415), .B(n416), .Z(n417) );
  XNOR U561 ( .A(n418), .B(n417), .Z(n411) );
  XOR U562 ( .A(n412), .B(n411), .Z(c[106]) );
  NANDN U563 ( .A(n410), .B(sreg[106]), .Z(n414) );
  NAND U564 ( .A(n412), .B(n411), .Z(n413) );
  AND U565 ( .A(n414), .B(n413), .Z(n467) );
  NANDN U566 ( .A(n416), .B(n415), .Z(n420) );
  NAND U567 ( .A(n418), .B(n417), .Z(n419) );
  AND U568 ( .A(n420), .B(n419), .Z(n473) );
  NANDN U569 ( .A(n422), .B(n421), .Z(n426) );
  NANDN U570 ( .A(n424), .B(n423), .Z(n425) );
  AND U571 ( .A(n426), .B(n425), .Z(n471) );
  NANDN U572 ( .A(n427), .B(n452), .Z(n431) );
  OR U573 ( .A(n429), .B(n428), .Z(n430) );
  AND U574 ( .A(n431), .B(n430), .Z(n516) );
  NANDN U575 ( .A(n433), .B(n432), .Z(n437) );
  NAND U576 ( .A(n435), .B(n434), .Z(n436) );
  AND U577 ( .A(n437), .B(n436), .Z(n479) );
  NANDN U578 ( .A(n17613), .B(n438), .Z(n440) );
  XOR U579 ( .A(b[9]), .B(a[3]), .Z(n491) );
  NANDN U580 ( .A(n17739), .B(n491), .Z(n439) );
  AND U581 ( .A(n440), .B(n439), .Z(n507) );
  XOR U582 ( .A(b[11]), .B(b[10]), .Z(n500) );
  XOR U583 ( .A(b[11]), .B(a[0]), .Z(n441) );
  NAND U584 ( .A(n500), .B(n441), .Z(n442) );
  OR U585 ( .A(n442), .B(n18085), .Z(n444) );
  XOR U586 ( .A(b[11]), .B(a[1]), .Z(n501) );
  NAND U587 ( .A(n18085), .B(n501), .Z(n443) );
  AND U588 ( .A(n444), .B(n443), .Z(n508) );
  XOR U589 ( .A(n507), .B(n508), .Z(n496) );
  NAND U590 ( .A(b[0]), .B(a[11]), .Z(n445) );
  XNOR U591 ( .A(b[1]), .B(n445), .Z(n447) );
  NANDN U592 ( .A(b[0]), .B(a[10]), .Z(n446) );
  NAND U593 ( .A(n447), .B(n446), .Z(n494) );
  NAND U594 ( .A(n17390), .B(n448), .Z(n450) );
  XNOR U595 ( .A(b[5]), .B(a[7]), .Z(n504) );
  NANDN U596 ( .A(n504), .B(n17391), .Z(n449) );
  NAND U597 ( .A(n450), .B(n449), .Z(n495) );
  XOR U598 ( .A(n494), .B(n495), .Z(n497) );
  XOR U599 ( .A(n496), .B(n497), .Z(n477) );
  NAND U600 ( .A(b[9]), .B(b[10]), .Z(n451) );
  AND U601 ( .A(b[11]), .B(n451), .Z(n18319) );
  ANDN U602 ( .B(n18319), .A(n452), .Z(n483) );
  NAND U603 ( .A(n17623), .B(n453), .Z(n455) );
  XNOR U604 ( .A(b[7]), .B(a[5]), .Z(n512) );
  NANDN U605 ( .A(n512), .B(n17624), .Z(n454) );
  NAND U606 ( .A(n455), .B(n454), .Z(n482) );
  XOR U607 ( .A(n483), .B(n482), .Z(n485) );
  NANDN U608 ( .A(n456), .B(n2664), .Z(n458) );
  XNOR U609 ( .A(b[3]), .B(a[9]), .Z(n509) );
  NANDN U610 ( .A(n509), .B(n2512), .Z(n457) );
  NAND U611 ( .A(n458), .B(n457), .Z(n484) );
  XOR U612 ( .A(n485), .B(n484), .Z(n476) );
  XNOR U613 ( .A(n477), .B(n476), .Z(n478) );
  XNOR U614 ( .A(n479), .B(n478), .Z(n515) );
  XNOR U615 ( .A(n516), .B(n515), .Z(n518) );
  NANDN U616 ( .A(n460), .B(n459), .Z(n464) );
  NANDN U617 ( .A(n462), .B(n461), .Z(n463) );
  AND U618 ( .A(n464), .B(n463), .Z(n517) );
  XNOR U619 ( .A(n518), .B(n517), .Z(n470) );
  XNOR U620 ( .A(n471), .B(n470), .Z(n472) );
  XNOR U621 ( .A(n473), .B(n472), .Z(n465) );
  XNOR U622 ( .A(sreg[107]), .B(n465), .Z(n466) );
  XNOR U623 ( .A(n467), .B(n466), .Z(c[107]) );
  NANDN U624 ( .A(sreg[107]), .B(n465), .Z(n469) );
  NAND U625 ( .A(n467), .B(n466), .Z(n468) );
  NAND U626 ( .A(n469), .B(n468), .Z(n580) );
  XNOR U627 ( .A(sreg[108]), .B(n580), .Z(n582) );
  NANDN U628 ( .A(n471), .B(n470), .Z(n475) );
  NANDN U629 ( .A(n473), .B(n472), .Z(n474) );
  AND U630 ( .A(n475), .B(n474), .Z(n523) );
  NANDN U631 ( .A(n477), .B(n476), .Z(n481) );
  NANDN U632 ( .A(n479), .B(n478), .Z(n480) );
  AND U633 ( .A(n481), .B(n480), .Z(n575) );
  NAND U634 ( .A(n483), .B(n482), .Z(n487) );
  NAND U635 ( .A(n485), .B(n484), .Z(n486) );
  NAND U636 ( .A(n487), .B(n486), .Z(n574) );
  XNOR U637 ( .A(n575), .B(n574), .Z(n577) );
  NAND U638 ( .A(b[0]), .B(a[12]), .Z(n488) );
  XNOR U639 ( .A(b[1]), .B(n488), .Z(n490) );
  NANDN U640 ( .A(b[0]), .B(a[11]), .Z(n489) );
  NAND U641 ( .A(n490), .B(n489), .Z(n565) );
  XOR U642 ( .A(b[11]), .B(b[12]), .Z(n18345) );
  IV U643 ( .A(n18345), .Z(n18229) );
  ANDN U644 ( .B(a[0]), .A(n18229), .Z(n562) );
  NANDN U645 ( .A(n17613), .B(n491), .Z(n493) );
  XOR U646 ( .A(b[9]), .B(a[4]), .Z(n555) );
  NANDN U647 ( .A(n17739), .B(n555), .Z(n492) );
  AND U648 ( .A(n493), .B(n492), .Z(n563) );
  XNOR U649 ( .A(n562), .B(n563), .Z(n564) );
  XNOR U650 ( .A(n565), .B(n564), .Z(n527) );
  NANDN U651 ( .A(n495), .B(n494), .Z(n499) );
  OR U652 ( .A(n497), .B(n496), .Z(n498) );
  NAND U653 ( .A(n499), .B(n498), .Z(n528) );
  XNOR U654 ( .A(n527), .B(n528), .Z(n529) );
  ANDN U655 ( .B(n500), .A(n18085), .Z(n18084) );
  IV U656 ( .A(n18084), .Z(n17888) );
  NANDN U657 ( .A(n17888), .B(n501), .Z(n503) );
  XOR U658 ( .A(b[11]), .B(a[2]), .Z(n549) );
  NANDN U659 ( .A(n18025), .B(n549), .Z(n502) );
  AND U660 ( .A(n503), .B(n502), .Z(n536) );
  NANDN U661 ( .A(n504), .B(n17390), .Z(n506) );
  XOR U662 ( .A(b[5]), .B(a[8]), .Z(n559) );
  NANDN U663 ( .A(n17223), .B(n559), .Z(n505) );
  AND U664 ( .A(n506), .B(n505), .Z(n534) );
  NOR U665 ( .A(n508), .B(n507), .Z(n570) );
  NANDN U666 ( .A(n509), .B(n2664), .Z(n511) );
  XNOR U667 ( .A(b[3]), .B(a[10]), .Z(n552) );
  NANDN U668 ( .A(n552), .B(n2512), .Z(n510) );
  AND U669 ( .A(n511), .B(n510), .Z(n568) );
  NANDN U670 ( .A(n512), .B(n17623), .Z(n514) );
  XNOR U671 ( .A(b[7]), .B(a[6]), .Z(n539) );
  NANDN U672 ( .A(n539), .B(n17624), .Z(n513) );
  NAND U673 ( .A(n514), .B(n513), .Z(n569) );
  XOR U674 ( .A(n568), .B(n569), .Z(n571) );
  XNOR U675 ( .A(n570), .B(n571), .Z(n533) );
  XNOR U676 ( .A(n534), .B(n533), .Z(n535) );
  XOR U677 ( .A(n536), .B(n535), .Z(n530) );
  XNOR U678 ( .A(n529), .B(n530), .Z(n576) );
  XOR U679 ( .A(n577), .B(n576), .Z(n522) );
  NANDN U680 ( .A(n516), .B(n515), .Z(n520) );
  NAND U681 ( .A(n518), .B(n517), .Z(n519) );
  AND U682 ( .A(n520), .B(n519), .Z(n521) );
  XOR U683 ( .A(n522), .B(n521), .Z(n524) );
  XNOR U684 ( .A(n523), .B(n524), .Z(n581) );
  XOR U685 ( .A(n582), .B(n581), .Z(c[108]) );
  NANDN U686 ( .A(n522), .B(n521), .Z(n526) );
  OR U687 ( .A(n524), .B(n523), .Z(n525) );
  AND U688 ( .A(n526), .B(n525), .Z(n592) );
  NANDN U689 ( .A(n528), .B(n527), .Z(n532) );
  NANDN U690 ( .A(n530), .B(n529), .Z(n531) );
  AND U691 ( .A(n532), .B(n531), .Z(n646) );
  NANDN U692 ( .A(n534), .B(n533), .Z(n538) );
  NANDN U693 ( .A(n536), .B(n535), .Z(n537) );
  AND U694 ( .A(n538), .B(n537), .Z(n645) );
  NANDN U695 ( .A(n539), .B(n17623), .Z(n541) );
  XOR U696 ( .A(b[7]), .B(a[7]), .Z(n623) );
  NANDN U697 ( .A(n17522), .B(n623), .Z(n540) );
  NAND U698 ( .A(n541), .B(n540), .Z(n629) );
  NAND U699 ( .A(b[0]), .B(a[13]), .Z(n542) );
  XNOR U700 ( .A(b[1]), .B(n542), .Z(n544) );
  NANDN U701 ( .A(b[0]), .B(a[12]), .Z(n543) );
  NAND U702 ( .A(n544), .B(n543), .Z(n630) );
  XNOR U703 ( .A(n629), .B(n630), .Z(n632) );
  XOR U704 ( .A(b[13]), .B(b[12]), .Z(n635) );
  XOR U705 ( .A(b[13]), .B(a[0]), .Z(n545) );
  NAND U706 ( .A(n635), .B(n545), .Z(n546) );
  OR U707 ( .A(n546), .B(n18345), .Z(n548) );
  XOR U708 ( .A(b[13]), .B(a[1]), .Z(n636) );
  NAND U709 ( .A(n18345), .B(n636), .Z(n547) );
  AND U710 ( .A(n548), .B(n547), .Z(n642) );
  NANDN U711 ( .A(n17888), .B(n549), .Z(n551) );
  XOR U712 ( .A(b[11]), .B(a[3]), .Z(n617) );
  NANDN U713 ( .A(n18025), .B(n617), .Z(n550) );
  NAND U714 ( .A(n551), .B(n550), .Z(n643) );
  XNOR U715 ( .A(n642), .B(n643), .Z(n631) );
  XOR U716 ( .A(n632), .B(n631), .Z(n604) );
  NANDN U717 ( .A(n552), .B(n2664), .Z(n554) );
  XOR U718 ( .A(b[3]), .B(a[11]), .Z(n626) );
  NANDN U719 ( .A(n17068), .B(n626), .Z(n553) );
  AND U720 ( .A(n554), .B(n553), .Z(n609) );
  NANDN U721 ( .A(n17613), .B(n555), .Z(n557) );
  XOR U722 ( .A(b[9]), .B(a[5]), .Z(n639) );
  NANDN U723 ( .A(n17739), .B(n639), .Z(n556) );
  NAND U724 ( .A(n557), .B(n556), .Z(n608) );
  XNOR U725 ( .A(n609), .B(n608), .Z(n611) );
  NAND U726 ( .A(b[11]), .B(b[12]), .Z(n558) );
  AND U727 ( .A(b[13]), .B(n558), .Z(n18481) );
  ANDN U728 ( .B(n18481), .A(n562), .Z(n610) );
  XOR U729 ( .A(n611), .B(n610), .Z(n603) );
  NAND U730 ( .A(n17390), .B(n559), .Z(n561) );
  XNOR U731 ( .A(b[5]), .B(a[9]), .Z(n620) );
  NANDN U732 ( .A(n620), .B(n17391), .Z(n560) );
  AND U733 ( .A(n561), .B(n560), .Z(n602) );
  XOR U734 ( .A(n603), .B(n602), .Z(n605) );
  XOR U735 ( .A(n604), .B(n605), .Z(n599) );
  NANDN U736 ( .A(n563), .B(n562), .Z(n567) );
  NANDN U737 ( .A(n565), .B(n564), .Z(n566) );
  AND U738 ( .A(n567), .B(n566), .Z(n597) );
  NANDN U739 ( .A(n569), .B(n568), .Z(n573) );
  OR U740 ( .A(n571), .B(n570), .Z(n572) );
  AND U741 ( .A(n573), .B(n572), .Z(n596) );
  XNOR U742 ( .A(n597), .B(n596), .Z(n598) );
  XNOR U743 ( .A(n599), .B(n598), .Z(n644) );
  XOR U744 ( .A(n645), .B(n644), .Z(n647) );
  XOR U745 ( .A(n646), .B(n647), .Z(n591) );
  NANDN U746 ( .A(n575), .B(n574), .Z(n579) );
  NAND U747 ( .A(n577), .B(n576), .Z(n578) );
  AND U748 ( .A(n579), .B(n578), .Z(n590) );
  XOR U749 ( .A(n591), .B(n590), .Z(n593) );
  XOR U750 ( .A(n592), .B(n593), .Z(n585) );
  XNOR U751 ( .A(n585), .B(sreg[109]), .Z(n587) );
  NANDN U752 ( .A(n580), .B(sreg[108]), .Z(n584) );
  NAND U753 ( .A(n582), .B(n581), .Z(n583) );
  NAND U754 ( .A(n584), .B(n583), .Z(n586) );
  XOR U755 ( .A(n587), .B(n586), .Z(c[109]) );
  NANDN U756 ( .A(n585), .B(sreg[109]), .Z(n589) );
  NAND U757 ( .A(n587), .B(n586), .Z(n588) );
  AND U758 ( .A(n589), .B(n588), .Z(n716) );
  XNOR U759 ( .A(sreg[110]), .B(n716), .Z(n718) );
  NANDN U760 ( .A(n591), .B(n590), .Z(n595) );
  OR U761 ( .A(n593), .B(n592), .Z(n594) );
  AND U762 ( .A(n595), .B(n594), .Z(n653) );
  NANDN U763 ( .A(n597), .B(n596), .Z(n601) );
  NANDN U764 ( .A(n599), .B(n598), .Z(n600) );
  AND U765 ( .A(n601), .B(n600), .Z(n712) );
  NANDN U766 ( .A(n603), .B(n602), .Z(n607) );
  OR U767 ( .A(n605), .B(n604), .Z(n606) );
  AND U768 ( .A(n607), .B(n606), .Z(n710) );
  NANDN U769 ( .A(n609), .B(n608), .Z(n613) );
  NAND U770 ( .A(n611), .B(n610), .Z(n612) );
  AND U771 ( .A(n613), .B(n612), .Z(n697) );
  NAND U772 ( .A(b[0]), .B(a[14]), .Z(n614) );
  XNOR U773 ( .A(b[1]), .B(n614), .Z(n616) );
  NANDN U774 ( .A(b[0]), .B(a[13]), .Z(n615) );
  NAND U775 ( .A(n616), .B(n615), .Z(n703) );
  XOR U776 ( .A(b[13]), .B(b[14]), .Z(n18486) );
  IV U777 ( .A(n18486), .Z(n18311) );
  ANDN U778 ( .B(a[0]), .A(n18311), .Z(n700) );
  NANDN U779 ( .A(n17888), .B(n617), .Z(n619) );
  XOR U780 ( .A(b[11]), .B(a[4]), .Z(n671) );
  NANDN U781 ( .A(n18025), .B(n671), .Z(n618) );
  AND U782 ( .A(n619), .B(n618), .Z(n701) );
  XNOR U783 ( .A(n700), .B(n701), .Z(n702) );
  XNOR U784 ( .A(n703), .B(n702), .Z(n694) );
  NANDN U785 ( .A(n620), .B(n17390), .Z(n622) );
  XOR U786 ( .A(b[5]), .B(a[10]), .Z(n665) );
  NANDN U787 ( .A(n17223), .B(n665), .Z(n621) );
  AND U788 ( .A(n622), .B(n621), .Z(n691) );
  NANDN U789 ( .A(n17362), .B(n623), .Z(n625) );
  XOR U790 ( .A(b[7]), .B(a[8]), .Z(n662) );
  NANDN U791 ( .A(n17522), .B(n662), .Z(n624) );
  AND U792 ( .A(n625), .B(n624), .Z(n689) );
  NANDN U793 ( .A(n17067), .B(n626), .Z(n628) );
  XOR U794 ( .A(b[3]), .B(a[12]), .Z(n668) );
  NANDN U795 ( .A(n17068), .B(n668), .Z(n627) );
  NAND U796 ( .A(n628), .B(n627), .Z(n688) );
  XNOR U797 ( .A(n689), .B(n688), .Z(n690) );
  XOR U798 ( .A(n691), .B(n690), .Z(n695) );
  XNOR U799 ( .A(n694), .B(n695), .Z(n696) );
  XNOR U800 ( .A(n697), .B(n696), .Z(n658) );
  NANDN U801 ( .A(n630), .B(n629), .Z(n634) );
  NAND U802 ( .A(n632), .B(n631), .Z(n633) );
  AND U803 ( .A(n634), .B(n633), .Z(n657) );
  ANDN U804 ( .B(n635), .A(n18345), .Z(n18347) );
  IV U805 ( .A(n18347), .Z(n18113) );
  NANDN U806 ( .A(n18113), .B(n636), .Z(n638) );
  XOR U807 ( .A(b[13]), .B(a[2]), .Z(n681) );
  NANDN U808 ( .A(n18229), .B(n681), .Z(n637) );
  AND U809 ( .A(n638), .B(n637), .Z(n707) );
  NANDN U810 ( .A(n17613), .B(n639), .Z(n641) );
  XOR U811 ( .A(b[9]), .B(a[6]), .Z(n675) );
  NANDN U812 ( .A(n17739), .B(n675), .Z(n640) );
  NAND U813 ( .A(n641), .B(n640), .Z(n706) );
  XNOR U814 ( .A(n707), .B(n706), .Z(n709) );
  ANDN U815 ( .B(n643), .A(n642), .Z(n708) );
  XOR U816 ( .A(n709), .B(n708), .Z(n656) );
  XOR U817 ( .A(n657), .B(n656), .Z(n659) );
  XOR U818 ( .A(n658), .B(n659), .Z(n711) );
  XOR U819 ( .A(n710), .B(n711), .Z(n713) );
  XOR U820 ( .A(n712), .B(n713), .Z(n651) );
  NANDN U821 ( .A(n645), .B(n644), .Z(n649) );
  OR U822 ( .A(n647), .B(n646), .Z(n648) );
  AND U823 ( .A(n649), .B(n648), .Z(n650) );
  XNOR U824 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U825 ( .A(n653), .B(n652), .Z(n717) );
  XNOR U826 ( .A(n718), .B(n717), .Z(c[110]) );
  NANDN U827 ( .A(n651), .B(n650), .Z(n655) );
  NANDN U828 ( .A(n653), .B(n652), .Z(n654) );
  AND U829 ( .A(n655), .B(n654), .Z(n723) );
  NANDN U830 ( .A(n657), .B(n656), .Z(n661) );
  NANDN U831 ( .A(n659), .B(n658), .Z(n660) );
  AND U832 ( .A(n661), .B(n660), .Z(n785) );
  NANDN U833 ( .A(n17362), .B(n662), .Z(n664) );
  XOR U834 ( .A(b[7]), .B(a[9]), .Z(n747) );
  NANDN U835 ( .A(n17522), .B(n747), .Z(n663) );
  AND U836 ( .A(n664), .B(n663), .Z(n734) );
  NANDN U837 ( .A(n17072), .B(n665), .Z(n667) );
  XOR U838 ( .A(b[5]), .B(a[11]), .Z(n757) );
  NANDN U839 ( .A(n17223), .B(n757), .Z(n666) );
  AND U840 ( .A(n667), .B(n666), .Z(n763) );
  NANDN U841 ( .A(n17067), .B(n668), .Z(n670) );
  XOR U842 ( .A(b[3]), .B(a[13]), .Z(n741) );
  NANDN U843 ( .A(n17068), .B(n741), .Z(n669) );
  AND U844 ( .A(n670), .B(n669), .Z(n761) );
  NANDN U845 ( .A(n17888), .B(n671), .Z(n673) );
  XOR U846 ( .A(b[11]), .B(a[5]), .Z(n750) );
  NANDN U847 ( .A(n18025), .B(n750), .Z(n672) );
  NAND U848 ( .A(n673), .B(n672), .Z(n760) );
  XNOR U849 ( .A(n761), .B(n760), .Z(n762) );
  XNOR U850 ( .A(n763), .B(n762), .Z(n733) );
  XNOR U851 ( .A(n734), .B(n733), .Z(n736) );
  NAND U852 ( .A(b[13]), .B(b[14]), .Z(n674) );
  AND U853 ( .A(b[15]), .B(n674), .Z(n18700) );
  ANDN U854 ( .B(n18700), .A(n700), .Z(n735) );
  XOR U855 ( .A(n736), .B(n735), .Z(n780) );
  NANDN U856 ( .A(n17613), .B(n675), .Z(n677) );
  XOR U857 ( .A(b[9]), .B(a[7]), .Z(n744) );
  NANDN U858 ( .A(n17739), .B(n744), .Z(n676) );
  NAND U859 ( .A(n677), .B(n676), .Z(n766) );
  NAND U860 ( .A(b[0]), .B(a[15]), .Z(n678) );
  XNOR U861 ( .A(b[1]), .B(n678), .Z(n680) );
  NANDN U862 ( .A(b[0]), .B(a[14]), .Z(n679) );
  NAND U863 ( .A(n680), .B(n679), .Z(n767) );
  XNOR U864 ( .A(n766), .B(n767), .Z(n769) );
  NANDN U865 ( .A(n18113), .B(n681), .Z(n683) );
  XOR U866 ( .A(b[13]), .B(a[3]), .Z(n775) );
  NANDN U867 ( .A(n18229), .B(n775), .Z(n682) );
  AND U868 ( .A(n683), .B(n682), .Z(n739) );
  XOR U869 ( .A(b[15]), .B(b[14]), .Z(n753) );
  XOR U870 ( .A(b[15]), .B(a[0]), .Z(n684) );
  NAND U871 ( .A(n753), .B(n684), .Z(n685) );
  OR U872 ( .A(n685), .B(n18486), .Z(n687) );
  XOR U873 ( .A(b[15]), .B(a[1]), .Z(n754) );
  NAND U874 ( .A(n18486), .B(n754), .Z(n686) );
  NAND U875 ( .A(n687), .B(n686), .Z(n740) );
  XNOR U876 ( .A(n739), .B(n740), .Z(n768) );
  XOR U877 ( .A(n769), .B(n768), .Z(n779) );
  NANDN U878 ( .A(n689), .B(n688), .Z(n693) );
  NANDN U879 ( .A(n691), .B(n690), .Z(n692) );
  AND U880 ( .A(n693), .B(n692), .Z(n778) );
  XOR U881 ( .A(n779), .B(n778), .Z(n781) );
  XNOR U882 ( .A(n780), .B(n781), .Z(n784) );
  XNOR U883 ( .A(n785), .B(n784), .Z(n787) );
  NANDN U884 ( .A(n695), .B(n694), .Z(n699) );
  NANDN U885 ( .A(n697), .B(n696), .Z(n698) );
  AND U886 ( .A(n699), .B(n698), .Z(n730) );
  NANDN U887 ( .A(n701), .B(n700), .Z(n705) );
  NANDN U888 ( .A(n703), .B(n702), .Z(n704) );
  AND U889 ( .A(n705), .B(n704), .Z(n728) );
  XNOR U890 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U891 ( .A(n730), .B(n729), .Z(n786) );
  XOR U892 ( .A(n787), .B(n786), .Z(n722) );
  NANDN U893 ( .A(n711), .B(n710), .Z(n715) );
  OR U894 ( .A(n713), .B(n712), .Z(n714) );
  AND U895 ( .A(n715), .B(n714), .Z(n721) );
  XOR U896 ( .A(n722), .B(n721), .Z(n724) );
  XOR U897 ( .A(n723), .B(n724), .Z(n790) );
  XNOR U898 ( .A(n790), .B(sreg[111]), .Z(n792) );
  NANDN U899 ( .A(sreg[110]), .B(n716), .Z(n720) );
  NAND U900 ( .A(n718), .B(n717), .Z(n719) );
  AND U901 ( .A(n720), .B(n719), .Z(n791) );
  XOR U902 ( .A(n792), .B(n791), .Z(c[111]) );
  NANDN U903 ( .A(n722), .B(n721), .Z(n726) );
  OR U904 ( .A(n724), .B(n723), .Z(n725) );
  AND U905 ( .A(n726), .B(n725), .Z(n801) );
  NANDN U906 ( .A(n728), .B(n727), .Z(n732) );
  NANDN U907 ( .A(n730), .B(n729), .Z(n731) );
  AND U908 ( .A(n732), .B(n731), .Z(n872) );
  NANDN U909 ( .A(n734), .B(n733), .Z(n738) );
  NAND U910 ( .A(n736), .B(n735), .Z(n737) );
  AND U911 ( .A(n738), .B(n737), .Z(n865) );
  ANDN U912 ( .B(n740), .A(n739), .Z(n839) );
  NAND U913 ( .A(n2664), .B(n741), .Z(n743) );
  XNOR U914 ( .A(b[3]), .B(a[14]), .Z(n828) );
  NANDN U915 ( .A(n828), .B(n2512), .Z(n742) );
  AND U916 ( .A(n743), .B(n742), .Z(n837) );
  NAND U917 ( .A(n17881), .B(n744), .Z(n746) );
  XNOR U918 ( .A(b[9]), .B(a[8]), .Z(n819) );
  NANDN U919 ( .A(n819), .B(n17879), .Z(n745) );
  NAND U920 ( .A(n746), .B(n745), .Z(n838) );
  XOR U921 ( .A(n837), .B(n838), .Z(n840) );
  XOR U922 ( .A(n839), .B(n840), .Z(n834) );
  NANDN U923 ( .A(n17362), .B(n747), .Z(n749) );
  XOR U924 ( .A(b[7]), .B(a[10]), .Z(n849) );
  NANDN U925 ( .A(n17522), .B(n849), .Z(n748) );
  AND U926 ( .A(n749), .B(n748), .Z(n832) );
  NANDN U927 ( .A(n17888), .B(n750), .Z(n752) );
  XOR U928 ( .A(b[11]), .B(a[6]), .Z(n843) );
  NANDN U929 ( .A(n18025), .B(n843), .Z(n751) );
  AND U930 ( .A(n752), .B(n751), .Z(n855) );
  ANDN U931 ( .B(n753), .A(n18486), .Z(n18439) );
  IV U932 ( .A(n18439), .Z(n18487) );
  NANDN U933 ( .A(n18487), .B(n754), .Z(n756) );
  XOR U934 ( .A(b[15]), .B(a[2]), .Z(n814) );
  NANDN U935 ( .A(n18311), .B(n814), .Z(n755) );
  AND U936 ( .A(n756), .B(n755), .Z(n853) );
  NANDN U937 ( .A(n17072), .B(n757), .Z(n759) );
  XOR U938 ( .A(b[5]), .B(a[12]), .Z(n825) );
  NANDN U939 ( .A(n17223), .B(n825), .Z(n758) );
  NAND U940 ( .A(n759), .B(n758), .Z(n852) );
  XNOR U941 ( .A(n853), .B(n852), .Z(n854) );
  XNOR U942 ( .A(n855), .B(n854), .Z(n831) );
  XNOR U943 ( .A(n832), .B(n831), .Z(n833) );
  XNOR U944 ( .A(n834), .B(n833), .Z(n864) );
  XNOR U945 ( .A(n865), .B(n864), .Z(n866) );
  NANDN U946 ( .A(n761), .B(n760), .Z(n765) );
  NANDN U947 ( .A(n763), .B(n762), .Z(n764) );
  AND U948 ( .A(n765), .B(n764), .Z(n861) );
  NANDN U949 ( .A(n767), .B(n766), .Z(n771) );
  NAND U950 ( .A(n769), .B(n768), .Z(n770) );
  AND U951 ( .A(n771), .B(n770), .Z(n859) );
  NAND U952 ( .A(b[0]), .B(a[16]), .Z(n772) );
  XNOR U953 ( .A(b[1]), .B(n772), .Z(n774) );
  NANDN U954 ( .A(b[0]), .B(a[15]), .Z(n773) );
  NAND U955 ( .A(n774), .B(n773), .Z(n806) );
  XOR U956 ( .A(b[16]), .B(b[15]), .Z(n18684) );
  IV U957 ( .A(n18684), .Z(n18585) );
  ANDN U958 ( .B(a[0]), .A(n18585), .Z(n818) );
  NANDN U959 ( .A(n18113), .B(n775), .Z(n777) );
  XOR U960 ( .A(b[13]), .B(a[4]), .Z(n846) );
  NANDN U961 ( .A(n18229), .B(n846), .Z(n776) );
  AND U962 ( .A(n777), .B(n776), .Z(n804) );
  XNOR U963 ( .A(n818), .B(n804), .Z(n805) );
  XNOR U964 ( .A(n806), .B(n805), .Z(n858) );
  XNOR U965 ( .A(n859), .B(n858), .Z(n860) );
  XOR U966 ( .A(n861), .B(n860), .Z(n867) );
  XNOR U967 ( .A(n866), .B(n867), .Z(n870) );
  NANDN U968 ( .A(n779), .B(n778), .Z(n783) );
  OR U969 ( .A(n781), .B(n780), .Z(n782) );
  NAND U970 ( .A(n783), .B(n782), .Z(n871) );
  XOR U971 ( .A(n870), .B(n871), .Z(n873) );
  XOR U972 ( .A(n872), .B(n873), .Z(n799) );
  NANDN U973 ( .A(n785), .B(n784), .Z(n789) );
  NAND U974 ( .A(n787), .B(n786), .Z(n788) );
  AND U975 ( .A(n789), .B(n788), .Z(n798) );
  XNOR U976 ( .A(n799), .B(n798), .Z(n800) );
  XNOR U977 ( .A(n801), .B(n800), .Z(n797) );
  NANDN U978 ( .A(n790), .B(sreg[111]), .Z(n794) );
  NAND U979 ( .A(n792), .B(n791), .Z(n793) );
  NAND U980 ( .A(n794), .B(n793), .Z(n796) );
  XOR U981 ( .A(n796), .B(sreg[112]), .Z(n795) );
  XNOR U982 ( .A(n797), .B(n795), .Z(c[112]) );
  NANDN U983 ( .A(n799), .B(n798), .Z(n803) );
  NANDN U984 ( .A(n801), .B(n800), .Z(n802) );
  AND U985 ( .A(n803), .B(n802), .Z(n884) );
  NANDN U986 ( .A(n804), .B(n818), .Z(n808) );
  NANDN U987 ( .A(n806), .B(n805), .Z(n807) );
  AND U988 ( .A(n808), .B(n807), .Z(n901) );
  XOR U989 ( .A(b[17]), .B(a[0]), .Z(n811) );
  XOR U990 ( .A(b[17]), .B(b[15]), .Z(n809) );
  XOR U991 ( .A(b[17]), .B(b[16]), .Z(n937) );
  AND U992 ( .A(n809), .B(n937), .Z(n810) );
  NAND U993 ( .A(n811), .B(n810), .Z(n813) );
  XOR U994 ( .A(b[17]), .B(a[1]), .Z(n938) );
  NANDN U995 ( .A(n18585), .B(n938), .Z(n812) );
  AND U996 ( .A(n813), .B(n812), .Z(n933) );
  NANDN U997 ( .A(n18487), .B(n814), .Z(n816) );
  XOR U998 ( .A(b[15]), .B(a[3]), .Z(n944) );
  NANDN U999 ( .A(n18311), .B(n944), .Z(n815) );
  AND U1000 ( .A(n816), .B(n815), .Z(n932) );
  XOR U1001 ( .A(n933), .B(n932), .Z(n949) );
  NAND U1002 ( .A(b[15]), .B(b[16]), .Z(n817) );
  NAND U1003 ( .A(b[17]), .B(n817), .Z(n18765) );
  NOR U1004 ( .A(n18765), .B(n818), .Z(n948) );
  NANDN U1005 ( .A(n819), .B(n17881), .Z(n821) );
  XNOR U1006 ( .A(b[9]), .B(a[9]), .Z(n923) );
  NANDN U1007 ( .A(n923), .B(n17879), .Z(n820) );
  AND U1008 ( .A(n821), .B(n820), .Z(n947) );
  XOR U1009 ( .A(n948), .B(n947), .Z(n950) );
  XOR U1010 ( .A(n949), .B(n950), .Z(n900) );
  NAND U1011 ( .A(b[0]), .B(a[17]), .Z(n822) );
  XNOR U1012 ( .A(b[1]), .B(n822), .Z(n824) );
  NANDN U1013 ( .A(b[0]), .B(a[16]), .Z(n823) );
  NAND U1014 ( .A(n824), .B(n823), .Z(n906) );
  NANDN U1015 ( .A(n17072), .B(n825), .Z(n827) );
  XOR U1016 ( .A(b[5]), .B(a[13]), .Z(n917) );
  NANDN U1017 ( .A(n17223), .B(n917), .Z(n826) );
  NAND U1018 ( .A(n827), .B(n826), .Z(n905) );
  XNOR U1019 ( .A(n906), .B(n905), .Z(n908) );
  NANDN U1020 ( .A(n828), .B(n2664), .Z(n830) );
  XNOR U1021 ( .A(b[3]), .B(a[15]), .Z(n929) );
  NANDN U1022 ( .A(n929), .B(n2512), .Z(n829) );
  NAND U1023 ( .A(n830), .B(n829), .Z(n907) );
  XOR U1024 ( .A(n908), .B(n907), .Z(n899) );
  XOR U1025 ( .A(n900), .B(n899), .Z(n902) );
  XOR U1026 ( .A(n901), .B(n902), .Z(n888) );
  NANDN U1027 ( .A(n832), .B(n831), .Z(n836) );
  NANDN U1028 ( .A(n834), .B(n833), .Z(n835) );
  AND U1029 ( .A(n836), .B(n835), .Z(n887) );
  XNOR U1030 ( .A(n888), .B(n887), .Z(n890) );
  NANDN U1031 ( .A(n838), .B(n837), .Z(n842) );
  OR U1032 ( .A(n840), .B(n839), .Z(n841) );
  AND U1033 ( .A(n842), .B(n841), .Z(n894) );
  NANDN U1034 ( .A(n17888), .B(n843), .Z(n845) );
  XOR U1035 ( .A(b[11]), .B(a[7]), .Z(n934) );
  NANDN U1036 ( .A(n18025), .B(n934), .Z(n844) );
  AND U1037 ( .A(n845), .B(n844), .Z(n913) );
  NANDN U1038 ( .A(n18113), .B(n846), .Z(n848) );
  XOR U1039 ( .A(b[13]), .B(a[5]), .Z(n926) );
  NANDN U1040 ( .A(n18229), .B(n926), .Z(n847) );
  AND U1041 ( .A(n848), .B(n847), .Z(n912) );
  NANDN U1042 ( .A(n17362), .B(n849), .Z(n851) );
  XOR U1043 ( .A(b[7]), .B(a[11]), .Z(n920) );
  NANDN U1044 ( .A(n17522), .B(n920), .Z(n850) );
  NAND U1045 ( .A(n851), .B(n850), .Z(n911) );
  XOR U1046 ( .A(n912), .B(n911), .Z(n914) );
  XNOR U1047 ( .A(n913), .B(n914), .Z(n893) );
  XNOR U1048 ( .A(n894), .B(n893), .Z(n895) );
  NANDN U1049 ( .A(n853), .B(n852), .Z(n857) );
  NANDN U1050 ( .A(n855), .B(n854), .Z(n856) );
  NAND U1051 ( .A(n857), .B(n856), .Z(n896) );
  XNOR U1052 ( .A(n895), .B(n896), .Z(n889) );
  XOR U1053 ( .A(n890), .B(n889), .Z(n955) );
  NANDN U1054 ( .A(n859), .B(n858), .Z(n863) );
  NANDN U1055 ( .A(n861), .B(n860), .Z(n862) );
  AND U1056 ( .A(n863), .B(n862), .Z(n954) );
  NANDN U1057 ( .A(n865), .B(n864), .Z(n869) );
  NANDN U1058 ( .A(n867), .B(n866), .Z(n868) );
  NAND U1059 ( .A(n869), .B(n868), .Z(n953) );
  XOR U1060 ( .A(n954), .B(n953), .Z(n956) );
  XOR U1061 ( .A(n955), .B(n956), .Z(n882) );
  NANDN U1062 ( .A(n871), .B(n870), .Z(n875) );
  OR U1063 ( .A(n873), .B(n872), .Z(n874) );
  AND U1064 ( .A(n875), .B(n874), .Z(n881) );
  XNOR U1065 ( .A(n882), .B(n881), .Z(n883) );
  XNOR U1066 ( .A(n884), .B(n883), .Z(n876) );
  XNOR U1067 ( .A(sreg[113]), .B(n876), .Z(n877) );
  XNOR U1068 ( .A(n878), .B(n877), .Z(c[113]) );
  NANDN U1069 ( .A(sreg[113]), .B(n876), .Z(n880) );
  NAND U1070 ( .A(n878), .B(n877), .Z(n879) );
  AND U1071 ( .A(n880), .B(n879), .Z(n960) );
  NANDN U1072 ( .A(n882), .B(n881), .Z(n886) );
  NANDN U1073 ( .A(n884), .B(n883), .Z(n885) );
  AND U1074 ( .A(n886), .B(n885), .Z(n965) );
  NANDN U1075 ( .A(n888), .B(n887), .Z(n892) );
  NAND U1076 ( .A(n890), .B(n889), .Z(n891) );
  AND U1077 ( .A(n892), .B(n891), .Z(n1047) );
  NANDN U1078 ( .A(n894), .B(n893), .Z(n898) );
  NANDN U1079 ( .A(n896), .B(n895), .Z(n897) );
  AND U1080 ( .A(n898), .B(n897), .Z(n1044) );
  NANDN U1081 ( .A(n900), .B(n899), .Z(n904) );
  OR U1082 ( .A(n902), .B(n901), .Z(n903) );
  AND U1083 ( .A(n904), .B(n903), .Z(n1039) );
  NANDN U1084 ( .A(n906), .B(n905), .Z(n910) );
  NAND U1085 ( .A(n908), .B(n907), .Z(n909) );
  NAND U1086 ( .A(n910), .B(n909), .Z(n1038) );
  XNOR U1087 ( .A(n1039), .B(n1038), .Z(n1040) );
  NANDN U1088 ( .A(n912), .B(n911), .Z(n916) );
  OR U1089 ( .A(n914), .B(n913), .Z(n915) );
  AND U1090 ( .A(n916), .B(n915), .Z(n1033) );
  NANDN U1091 ( .A(n17072), .B(n917), .Z(n919) );
  XOR U1092 ( .A(b[5]), .B(a[14]), .Z(n1020) );
  NANDN U1093 ( .A(n17223), .B(n1020), .Z(n918) );
  AND U1094 ( .A(n919), .B(n918), .Z(n1000) );
  NANDN U1095 ( .A(n17362), .B(n920), .Z(n922) );
  XOR U1096 ( .A(b[7]), .B(a[12]), .Z(n1011) );
  NANDN U1097 ( .A(n17522), .B(n1011), .Z(n921) );
  NAND U1098 ( .A(n922), .B(n921), .Z(n999) );
  XNOR U1099 ( .A(n1000), .B(n999), .Z(n1001) );
  NANDN U1100 ( .A(n923), .B(n17881), .Z(n925) );
  XOR U1101 ( .A(b[9]), .B(a[10]), .Z(n984) );
  NANDN U1102 ( .A(n17739), .B(n984), .Z(n924) );
  AND U1103 ( .A(n925), .B(n924), .Z(n990) );
  NANDN U1104 ( .A(n18113), .B(n926), .Z(n928) );
  XOR U1105 ( .A(b[13]), .B(a[6]), .Z(n1014) );
  NANDN U1106 ( .A(n18229), .B(n1014), .Z(n927) );
  AND U1107 ( .A(n928), .B(n927), .Z(n988) );
  NANDN U1108 ( .A(n929), .B(n2664), .Z(n931) );
  XOR U1109 ( .A(b[3]), .B(a[16]), .Z(n1023) );
  NANDN U1110 ( .A(n17068), .B(n1023), .Z(n930) );
  NAND U1111 ( .A(n931), .B(n930), .Z(n987) );
  XNOR U1112 ( .A(n988), .B(n987), .Z(n989) );
  XOR U1113 ( .A(n990), .B(n989), .Z(n1002) );
  XNOR U1114 ( .A(n1001), .B(n1002), .Z(n1032) );
  XNOR U1115 ( .A(n1033), .B(n1032), .Z(n1034) );
  NOR U1116 ( .A(n933), .B(n932), .Z(n995) );
  NAND U1117 ( .A(n18084), .B(n934), .Z(n936) );
  XNOR U1118 ( .A(b[11]), .B(a[8]), .Z(n1026) );
  NANDN U1119 ( .A(n1026), .B(n18085), .Z(n935) );
  AND U1120 ( .A(n936), .B(n935), .Z(n993) );
  ANDN U1121 ( .B(n937), .A(n18684), .Z(n18683) );
  NAND U1122 ( .A(n18683), .B(n938), .Z(n940) );
  XNOR U1123 ( .A(b[17]), .B(a[2]), .Z(n974) );
  NANDN U1124 ( .A(n974), .B(n18684), .Z(n939) );
  NAND U1125 ( .A(n940), .B(n939), .Z(n994) );
  XOR U1126 ( .A(n993), .B(n994), .Z(n996) );
  XOR U1127 ( .A(n995), .B(n996), .Z(n969) );
  NAND U1128 ( .A(b[0]), .B(a[18]), .Z(n941) );
  XNOR U1129 ( .A(b[1]), .B(n941), .Z(n943) );
  NANDN U1130 ( .A(b[0]), .B(a[17]), .Z(n942) );
  NAND U1131 ( .A(n943), .B(n942), .Z(n1008) );
  XOR U1132 ( .A(b[18]), .B(b[17]), .Z(n18882) );
  IV U1133 ( .A(n18882), .Z(n18758) );
  ANDN U1134 ( .B(a[0]), .A(n18758), .Z(n1005) );
  NANDN U1135 ( .A(n18487), .B(n944), .Z(n946) );
  XOR U1136 ( .A(b[15]), .B(a[4]), .Z(n1017) );
  NANDN U1137 ( .A(n18311), .B(n1017), .Z(n945) );
  AND U1138 ( .A(n946), .B(n945), .Z(n1006) );
  XNOR U1139 ( .A(n1005), .B(n1006), .Z(n1007) );
  XNOR U1140 ( .A(n1008), .B(n1007), .Z(n968) );
  XNOR U1141 ( .A(n969), .B(n968), .Z(n970) );
  NANDN U1142 ( .A(n948), .B(n947), .Z(n952) );
  OR U1143 ( .A(n950), .B(n949), .Z(n951) );
  NAND U1144 ( .A(n952), .B(n951), .Z(n971) );
  XOR U1145 ( .A(n970), .B(n971), .Z(n1035) );
  XOR U1146 ( .A(n1034), .B(n1035), .Z(n1041) );
  XOR U1147 ( .A(n1040), .B(n1041), .Z(n1045) );
  XNOR U1148 ( .A(n1044), .B(n1045), .Z(n1046) );
  XOR U1149 ( .A(n1047), .B(n1046), .Z(n963) );
  NANDN U1150 ( .A(n954), .B(n953), .Z(n958) );
  OR U1151 ( .A(n956), .B(n955), .Z(n957) );
  AND U1152 ( .A(n958), .B(n957), .Z(n962) );
  XNOR U1153 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U1154 ( .A(n965), .B(n964), .Z(n961) );
  XNOR U1155 ( .A(sreg[114]), .B(n961), .Z(n959) );
  XOR U1156 ( .A(n960), .B(n959), .Z(c[114]) );
  NANDN U1157 ( .A(n963), .B(n962), .Z(n967) );
  NANDN U1158 ( .A(n965), .B(n964), .Z(n966) );
  AND U1159 ( .A(n967), .B(n966), .Z(n1056) );
  NANDN U1160 ( .A(n969), .B(n968), .Z(n973) );
  NANDN U1161 ( .A(n971), .B(n970), .Z(n972) );
  AND U1162 ( .A(n973), .B(n972), .Z(n1066) );
  NANDN U1163 ( .A(n974), .B(n18683), .Z(n976) );
  XOR U1164 ( .A(b[17]), .B(a[3]), .Z(n1080) );
  NANDN U1165 ( .A(n18585), .B(n1080), .Z(n975) );
  AND U1166 ( .A(n976), .B(n975), .Z(n1104) );
  XOR U1167 ( .A(b[19]), .B(a[1]), .Z(n1110) );
  NANDN U1168 ( .A(n18758), .B(n1110), .Z(n983) );
  ANDN U1169 ( .B(b[18]), .A(b[19]), .Z(n977) );
  NAND U1170 ( .A(n977), .B(a[0]), .Z(n980) );
  NAND U1171 ( .A(b[17]), .B(b[18]), .Z(n978) );
  NAND U1172 ( .A(b[19]), .B(n978), .Z(n18979) );
  OR U1173 ( .A(a[0]), .B(n18979), .Z(n979) );
  NAND U1174 ( .A(n980), .B(n979), .Z(n981) );
  NAND U1175 ( .A(n18758), .B(n981), .Z(n982) );
  AND U1176 ( .A(n983), .B(n982), .Z(n1105) );
  XOR U1177 ( .A(n1104), .B(n1105), .Z(n1094) );
  NOR U1178 ( .A(n18979), .B(n1005), .Z(n1093) );
  NAND U1179 ( .A(n17881), .B(n984), .Z(n986) );
  XNOR U1180 ( .A(b[9]), .B(a[11]), .Z(n1113) );
  NANDN U1181 ( .A(n1113), .B(n17879), .Z(n985) );
  AND U1182 ( .A(n986), .B(n985), .Z(n1092) );
  XOR U1183 ( .A(n1093), .B(n1092), .Z(n1095) );
  XOR U1184 ( .A(n1094), .B(n1095), .Z(n1123) );
  NANDN U1185 ( .A(n988), .B(n987), .Z(n992) );
  NANDN U1186 ( .A(n990), .B(n989), .Z(n991) );
  NAND U1187 ( .A(n992), .B(n991), .Z(n1122) );
  XNOR U1188 ( .A(n1123), .B(n1122), .Z(n1124) );
  NANDN U1189 ( .A(n994), .B(n993), .Z(n998) );
  OR U1190 ( .A(n996), .B(n995), .Z(n997) );
  NAND U1191 ( .A(n998), .B(n997), .Z(n1125) );
  XNOR U1192 ( .A(n1124), .B(n1125), .Z(n1065) );
  XNOR U1193 ( .A(n1066), .B(n1065), .Z(n1068) );
  NANDN U1194 ( .A(n1000), .B(n999), .Z(n1004) );
  NANDN U1195 ( .A(n1002), .B(n1001), .Z(n1003) );
  AND U1196 ( .A(n1004), .B(n1003), .Z(n1060) );
  NANDN U1197 ( .A(n1006), .B(n1005), .Z(n1010) );
  NANDN U1198 ( .A(n1008), .B(n1007), .Z(n1009) );
  NAND U1199 ( .A(n1010), .B(n1009), .Z(n1059) );
  XNOR U1200 ( .A(n1060), .B(n1059), .Z(n1061) );
  NANDN U1201 ( .A(n17362), .B(n1011), .Z(n1013) );
  XOR U1202 ( .A(b[7]), .B(a[13]), .Z(n1086) );
  NANDN U1203 ( .A(n17522), .B(n1086), .Z(n1012) );
  AND U1204 ( .A(n1013), .B(n1012), .Z(n1129) );
  NANDN U1205 ( .A(n18113), .B(n1014), .Z(n1016) );
  XOR U1206 ( .A(b[13]), .B(a[7]), .Z(n1119) );
  NANDN U1207 ( .A(n18229), .B(n1119), .Z(n1015) );
  AND U1208 ( .A(n1016), .B(n1015), .Z(n1074) );
  NANDN U1209 ( .A(n18487), .B(n1017), .Z(n1019) );
  XOR U1210 ( .A(b[15]), .B(a[5]), .Z(n1116) );
  NANDN U1211 ( .A(n18311), .B(n1116), .Z(n1018) );
  AND U1212 ( .A(n1019), .B(n1018), .Z(n1072) );
  NANDN U1213 ( .A(n17072), .B(n1020), .Z(n1022) );
  XOR U1214 ( .A(b[5]), .B(a[15]), .Z(n1083) );
  NANDN U1215 ( .A(n17223), .B(n1083), .Z(n1021) );
  NAND U1216 ( .A(n1022), .B(n1021), .Z(n1071) );
  XNOR U1217 ( .A(n1072), .B(n1071), .Z(n1073) );
  XNOR U1218 ( .A(n1074), .B(n1073), .Z(n1128) );
  XNOR U1219 ( .A(n1129), .B(n1128), .Z(n1130) );
  NANDN U1220 ( .A(n17067), .B(n1023), .Z(n1025) );
  XOR U1221 ( .A(b[3]), .B(a[17]), .Z(n1089) );
  NANDN U1222 ( .A(n17068), .B(n1089), .Z(n1024) );
  AND U1223 ( .A(n1025), .B(n1024), .Z(n1101) );
  NANDN U1224 ( .A(n1026), .B(n18084), .Z(n1028) );
  XOR U1225 ( .A(b[11]), .B(a[9]), .Z(n1106) );
  NANDN U1226 ( .A(n18025), .B(n1106), .Z(n1027) );
  NAND U1227 ( .A(n1028), .B(n1027), .Z(n1098) );
  NAND U1228 ( .A(b[0]), .B(a[19]), .Z(n1029) );
  XNOR U1229 ( .A(b[1]), .B(n1029), .Z(n1031) );
  NANDN U1230 ( .A(b[0]), .B(a[18]), .Z(n1030) );
  NAND U1231 ( .A(n1031), .B(n1030), .Z(n1099) );
  XNOR U1232 ( .A(n1098), .B(n1099), .Z(n1100) );
  XOR U1233 ( .A(n1101), .B(n1100), .Z(n1131) );
  XOR U1234 ( .A(n1130), .B(n1131), .Z(n1062) );
  XNOR U1235 ( .A(n1061), .B(n1062), .Z(n1067) );
  XOR U1236 ( .A(n1068), .B(n1067), .Z(n1135) );
  NANDN U1237 ( .A(n1033), .B(n1032), .Z(n1037) );
  NANDN U1238 ( .A(n1035), .B(n1034), .Z(n1036) );
  AND U1239 ( .A(n1037), .B(n1036), .Z(n1134) );
  XNOR U1240 ( .A(n1135), .B(n1134), .Z(n1136) );
  NANDN U1241 ( .A(n1039), .B(n1038), .Z(n1043) );
  NANDN U1242 ( .A(n1041), .B(n1040), .Z(n1042) );
  NAND U1243 ( .A(n1043), .B(n1042), .Z(n1137) );
  XNOR U1244 ( .A(n1136), .B(n1137), .Z(n1053) );
  NANDN U1245 ( .A(n1045), .B(n1044), .Z(n1049) );
  NAND U1246 ( .A(n1047), .B(n1046), .Z(n1048) );
  NAND U1247 ( .A(n1049), .B(n1048), .Z(n1054) );
  XNOR U1248 ( .A(n1053), .B(n1054), .Z(n1055) );
  XOR U1249 ( .A(n1056), .B(n1055), .Z(n1051) );
  XOR U1250 ( .A(n1051), .B(sreg[115]), .Z(n1050) );
  XNOR U1251 ( .A(n1052), .B(n1050), .Z(c[115]) );
  XNOR U1252 ( .A(sreg[116]), .B(n1235), .Z(n1237) );
  NANDN U1253 ( .A(n1054), .B(n1053), .Z(n1058) );
  NANDN U1254 ( .A(n1056), .B(n1055), .Z(n1057) );
  AND U1255 ( .A(n1058), .B(n1057), .Z(n1143) );
  NANDN U1256 ( .A(n1060), .B(n1059), .Z(n1064) );
  NANDN U1257 ( .A(n1062), .B(n1061), .Z(n1063) );
  AND U1258 ( .A(n1064), .B(n1063), .Z(n1230) );
  NANDN U1259 ( .A(n1066), .B(n1065), .Z(n1070) );
  NAND U1260 ( .A(n1068), .B(n1067), .Z(n1069) );
  NAND U1261 ( .A(n1070), .B(n1069), .Z(n1229) );
  XNOR U1262 ( .A(n1230), .B(n1229), .Z(n1232) );
  NANDN U1263 ( .A(n1072), .B(n1071), .Z(n1076) );
  NANDN U1264 ( .A(n1074), .B(n1073), .Z(n1075) );
  AND U1265 ( .A(n1076), .B(n1075), .Z(n1225) );
  NAND U1266 ( .A(b[0]), .B(a[20]), .Z(n1077) );
  XNOR U1267 ( .A(b[1]), .B(n1077), .Z(n1079) );
  NANDN U1268 ( .A(b[0]), .B(a[19]), .Z(n1078) );
  NAND U1269 ( .A(n1079), .B(n1078), .Z(n1160) );
  XOR U1270 ( .A(b[20]), .B(b[19]), .Z(n18998) );
  IV U1271 ( .A(n18998), .Z(n18926) );
  ANDN U1272 ( .B(a[0]), .A(n18926), .Z(n1171) );
  IV U1273 ( .A(n18683), .Z(n18514) );
  NANDN U1274 ( .A(n18514), .B(n1080), .Z(n1082) );
  XOR U1275 ( .A(b[17]), .B(a[4]), .Z(n1199) );
  NANDN U1276 ( .A(n18585), .B(n1199), .Z(n1081) );
  AND U1277 ( .A(n1082), .B(n1081), .Z(n1158) );
  XNOR U1278 ( .A(n1171), .B(n1158), .Z(n1159) );
  XNOR U1279 ( .A(n1160), .B(n1159), .Z(n1223) );
  NANDN U1280 ( .A(n17072), .B(n1083), .Z(n1085) );
  XOR U1281 ( .A(b[5]), .B(a[16]), .Z(n1193) );
  NANDN U1282 ( .A(n17223), .B(n1193), .Z(n1084) );
  AND U1283 ( .A(n1085), .B(n1084), .Z(n1220) );
  NANDN U1284 ( .A(n17362), .B(n1086), .Z(n1088) );
  XOR U1285 ( .A(b[7]), .B(a[14]), .Z(n1190) );
  NANDN U1286 ( .A(n17522), .B(n1190), .Z(n1087) );
  AND U1287 ( .A(n1088), .B(n1087), .Z(n1218) );
  NANDN U1288 ( .A(n17067), .B(n1089), .Z(n1091) );
  XOR U1289 ( .A(b[3]), .B(a[18]), .Z(n1175) );
  NANDN U1290 ( .A(n17068), .B(n1175), .Z(n1090) );
  NAND U1291 ( .A(n1091), .B(n1090), .Z(n1217) );
  XNOR U1292 ( .A(n1218), .B(n1217), .Z(n1219) );
  XOR U1293 ( .A(n1220), .B(n1219), .Z(n1224) );
  XOR U1294 ( .A(n1223), .B(n1224), .Z(n1226) );
  XOR U1295 ( .A(n1225), .B(n1226), .Z(n1154) );
  NANDN U1296 ( .A(n1093), .B(n1092), .Z(n1097) );
  OR U1297 ( .A(n1095), .B(n1094), .Z(n1096) );
  AND U1298 ( .A(n1097), .B(n1096), .Z(n1153) );
  NANDN U1299 ( .A(n1099), .B(n1098), .Z(n1103) );
  NANDN U1300 ( .A(n1101), .B(n1100), .Z(n1102) );
  AND U1301 ( .A(n1103), .B(n1102), .Z(n1207) );
  NOR U1302 ( .A(n1105), .B(n1104), .Z(n1186) );
  NAND U1303 ( .A(n18084), .B(n1106), .Z(n1108) );
  XNOR U1304 ( .A(b[11]), .B(a[10]), .Z(n1172) );
  NANDN U1305 ( .A(n1172), .B(n18085), .Z(n1107) );
  AND U1306 ( .A(n1108), .B(n1107), .Z(n1184) );
  XOR U1307 ( .A(b[18]), .B(b[19]), .Z(n1109) );
  ANDN U1308 ( .B(n1109), .A(n18882), .Z(n18881) );
  NAND U1309 ( .A(n18881), .B(n1110), .Z(n1112) );
  XNOR U1310 ( .A(b[19]), .B(a[2]), .Z(n1163) );
  NANDN U1311 ( .A(n1163), .B(n18882), .Z(n1111) );
  NAND U1312 ( .A(n1112), .B(n1111), .Z(n1185) );
  XOR U1313 ( .A(n1184), .B(n1185), .Z(n1187) );
  XOR U1314 ( .A(n1186), .B(n1187), .Z(n1206) );
  NANDN U1315 ( .A(n1113), .B(n17881), .Z(n1115) );
  XNOR U1316 ( .A(b[9]), .B(a[12]), .Z(n1181) );
  NANDN U1317 ( .A(n1181), .B(n17879), .Z(n1114) );
  NAND U1318 ( .A(n1115), .B(n1114), .Z(n1212) );
  NANDN U1319 ( .A(n18487), .B(n1116), .Z(n1118) );
  XOR U1320 ( .A(b[15]), .B(a[6]), .Z(n1202) );
  NANDN U1321 ( .A(n18311), .B(n1202), .Z(n1117) );
  NAND U1322 ( .A(n1118), .B(n1117), .Z(n1211) );
  XOR U1323 ( .A(n1212), .B(n1211), .Z(n1214) );
  NAND U1324 ( .A(n18347), .B(n1119), .Z(n1121) );
  XNOR U1325 ( .A(b[13]), .B(a[8]), .Z(n1196) );
  NANDN U1326 ( .A(n1196), .B(n18345), .Z(n1120) );
  NAND U1327 ( .A(n1121), .B(n1120), .Z(n1213) );
  XOR U1328 ( .A(n1214), .B(n1213), .Z(n1205) );
  XOR U1329 ( .A(n1206), .B(n1205), .Z(n1208) );
  XNOR U1330 ( .A(n1207), .B(n1208), .Z(n1152) );
  XOR U1331 ( .A(n1153), .B(n1152), .Z(n1155) );
  XOR U1332 ( .A(n1154), .B(n1155), .Z(n1149) );
  NANDN U1333 ( .A(n1123), .B(n1122), .Z(n1127) );
  NANDN U1334 ( .A(n1125), .B(n1124), .Z(n1126) );
  AND U1335 ( .A(n1127), .B(n1126), .Z(n1147) );
  NANDN U1336 ( .A(n1129), .B(n1128), .Z(n1133) );
  NANDN U1337 ( .A(n1131), .B(n1130), .Z(n1132) );
  NAND U1338 ( .A(n1133), .B(n1132), .Z(n1146) );
  XNOR U1339 ( .A(n1147), .B(n1146), .Z(n1148) );
  XNOR U1340 ( .A(n1149), .B(n1148), .Z(n1231) );
  XOR U1341 ( .A(n1232), .B(n1231), .Z(n1141) );
  NANDN U1342 ( .A(n1135), .B(n1134), .Z(n1139) );
  NANDN U1343 ( .A(n1137), .B(n1136), .Z(n1138) );
  NAND U1344 ( .A(n1139), .B(n1138), .Z(n1140) );
  XNOR U1345 ( .A(n1141), .B(n1140), .Z(n1142) );
  XNOR U1346 ( .A(n1143), .B(n1142), .Z(n1236) );
  XNOR U1347 ( .A(n1237), .B(n1236), .Z(c[116]) );
  NANDN U1348 ( .A(n1141), .B(n1140), .Z(n1145) );
  NANDN U1349 ( .A(n1143), .B(n1142), .Z(n1144) );
  AND U1350 ( .A(n1145), .B(n1144), .Z(n1246) );
  NANDN U1351 ( .A(n1147), .B(n1146), .Z(n1151) );
  NANDN U1352 ( .A(n1149), .B(n1148), .Z(n1150) );
  AND U1353 ( .A(n1151), .B(n1150), .Z(n1332) );
  NANDN U1354 ( .A(n1153), .B(n1152), .Z(n1157) );
  OR U1355 ( .A(n1155), .B(n1154), .Z(n1156) );
  AND U1356 ( .A(n1157), .B(n1156), .Z(n1330) );
  NANDN U1357 ( .A(n1158), .B(n1171), .Z(n1162) );
  NANDN U1358 ( .A(n1160), .B(n1159), .Z(n1161) );
  NAND U1359 ( .A(n1162), .B(n1161), .Z(n1259) );
  NANDN U1360 ( .A(n1163), .B(n18881), .Z(n1165) );
  XOR U1361 ( .A(b[19]), .B(a[3]), .Z(n1292) );
  NANDN U1362 ( .A(n18758), .B(n1292), .Z(n1164) );
  AND U1363 ( .A(n1165), .B(n1164), .Z(n1287) );
  XOR U1364 ( .A(b[21]), .B(b[20]), .Z(n1307) );
  XOR U1365 ( .A(b[21]), .B(a[0]), .Z(n1166) );
  NAND U1366 ( .A(n1307), .B(n1166), .Z(n1167) );
  OR U1367 ( .A(n1167), .B(n18998), .Z(n1169) );
  XOR U1368 ( .A(b[21]), .B(a[1]), .Z(n1308) );
  NAND U1369 ( .A(n18998), .B(n1308), .Z(n1168) );
  AND U1370 ( .A(n1169), .B(n1168), .Z(n1288) );
  XOR U1371 ( .A(n1287), .B(n1288), .Z(n1278) );
  NAND U1372 ( .A(b[19]), .B(b[20]), .Z(n1170) );
  NAND U1373 ( .A(b[21]), .B(n1170), .Z(n19106) );
  NOR U1374 ( .A(n19106), .B(n1171), .Z(n1276) );
  NANDN U1375 ( .A(n1172), .B(n18084), .Z(n1174) );
  XNOR U1376 ( .A(b[11]), .B(a[11]), .Z(n1314) );
  NANDN U1377 ( .A(n1314), .B(n18085), .Z(n1173) );
  AND U1378 ( .A(n1174), .B(n1173), .Z(n1275) );
  XNOR U1379 ( .A(n1276), .B(n1275), .Z(n1277) );
  XOR U1380 ( .A(n1278), .B(n1277), .Z(n1257) );
  NANDN U1381 ( .A(n17067), .B(n1175), .Z(n1177) );
  XOR U1382 ( .A(b[3]), .B(a[19]), .Z(n1281) );
  NANDN U1383 ( .A(n17068), .B(n1281), .Z(n1176) );
  AND U1384 ( .A(n1177), .B(n1176), .Z(n1325) );
  NAND U1385 ( .A(b[0]), .B(a[21]), .Z(n1178) );
  XNOR U1386 ( .A(b[1]), .B(n1178), .Z(n1180) );
  NANDN U1387 ( .A(b[0]), .B(a[20]), .Z(n1179) );
  NAND U1388 ( .A(n1180), .B(n1179), .Z(n1324) );
  NANDN U1389 ( .A(n1181), .B(n17881), .Z(n1183) );
  XOR U1390 ( .A(b[9]), .B(a[13]), .Z(n1311) );
  NANDN U1391 ( .A(n17739), .B(n1311), .Z(n1182) );
  NAND U1392 ( .A(n1183), .B(n1182), .Z(n1323) );
  XOR U1393 ( .A(n1324), .B(n1323), .Z(n1326) );
  XOR U1394 ( .A(n1325), .B(n1326), .Z(n1258) );
  XOR U1395 ( .A(n1257), .B(n1258), .Z(n1260) );
  XNOR U1396 ( .A(n1259), .B(n1260), .Z(n1265) );
  NANDN U1397 ( .A(n1185), .B(n1184), .Z(n1189) );
  OR U1398 ( .A(n1187), .B(n1186), .Z(n1188) );
  AND U1399 ( .A(n1189), .B(n1188), .Z(n1264) );
  NANDN U1400 ( .A(n17362), .B(n1190), .Z(n1192) );
  XOR U1401 ( .A(b[7]), .B(a[15]), .Z(n1295) );
  NANDN U1402 ( .A(n17522), .B(n1295), .Z(n1191) );
  AND U1403 ( .A(n1192), .B(n1191), .Z(n1270) );
  NANDN U1404 ( .A(n17072), .B(n1193), .Z(n1195) );
  XOR U1405 ( .A(b[5]), .B(a[17]), .Z(n1298) );
  NANDN U1406 ( .A(n17223), .B(n1298), .Z(n1194) );
  NAND U1407 ( .A(n1195), .B(n1194), .Z(n1269) );
  XNOR U1408 ( .A(n1270), .B(n1269), .Z(n1272) );
  NANDN U1409 ( .A(n1196), .B(n18347), .Z(n1198) );
  XOR U1410 ( .A(b[13]), .B(a[9]), .Z(n1284) );
  NANDN U1411 ( .A(n18229), .B(n1284), .Z(n1197) );
  AND U1412 ( .A(n1198), .B(n1197), .Z(n1320) );
  NANDN U1413 ( .A(n18514), .B(n1199), .Z(n1201) );
  XOR U1414 ( .A(b[17]), .B(a[5]), .Z(n1304) );
  NANDN U1415 ( .A(n18585), .B(n1304), .Z(n1200) );
  AND U1416 ( .A(n1201), .B(n1200), .Z(n1318) );
  NANDN U1417 ( .A(n18487), .B(n1202), .Z(n1204) );
  XOR U1418 ( .A(b[15]), .B(a[7]), .Z(n1301) );
  NANDN U1419 ( .A(n18311), .B(n1301), .Z(n1203) );
  NAND U1420 ( .A(n1204), .B(n1203), .Z(n1317) );
  XNOR U1421 ( .A(n1318), .B(n1317), .Z(n1319) );
  XNOR U1422 ( .A(n1320), .B(n1319), .Z(n1271) );
  XNOR U1423 ( .A(n1272), .B(n1271), .Z(n1263) );
  XOR U1424 ( .A(n1264), .B(n1263), .Z(n1266) );
  XOR U1425 ( .A(n1265), .B(n1266), .Z(n1247) );
  NANDN U1426 ( .A(n1206), .B(n1205), .Z(n1210) );
  OR U1427 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1428 ( .A(n1210), .B(n1209), .Z(n1248) );
  XOR U1429 ( .A(n1247), .B(n1248), .Z(n1250) );
  NAND U1430 ( .A(n1212), .B(n1211), .Z(n1216) );
  NAND U1431 ( .A(n1214), .B(n1213), .Z(n1215) );
  NAND U1432 ( .A(n1216), .B(n1215), .Z(n1252) );
  NANDN U1433 ( .A(n1218), .B(n1217), .Z(n1222) );
  NANDN U1434 ( .A(n1220), .B(n1219), .Z(n1221) );
  NAND U1435 ( .A(n1222), .B(n1221), .Z(n1251) );
  XOR U1436 ( .A(n1252), .B(n1251), .Z(n1254) );
  NANDN U1437 ( .A(n1224), .B(n1223), .Z(n1228) );
  OR U1438 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U1439 ( .A(n1228), .B(n1227), .Z(n1253) );
  XOR U1440 ( .A(n1254), .B(n1253), .Z(n1249) );
  XOR U1441 ( .A(n1250), .B(n1249), .Z(n1329) );
  XOR U1442 ( .A(n1330), .B(n1329), .Z(n1331) );
  XOR U1443 ( .A(n1332), .B(n1331), .Z(n1243) );
  NANDN U1444 ( .A(n1230), .B(n1229), .Z(n1234) );
  NAND U1445 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U1446 ( .A(n1234), .B(n1233), .Z(n1244) );
  XOR U1447 ( .A(n1243), .B(n1244), .Z(n1245) );
  XOR U1448 ( .A(n1246), .B(n1245), .Z(n1241) );
  NANDN U1449 ( .A(sreg[116]), .B(n1235), .Z(n1239) );
  NAND U1450 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U1451 ( .A(n1239), .B(n1238), .Z(n1242) );
  XNOR U1452 ( .A(sreg[117]), .B(n1242), .Z(n1240) );
  XNOR U1453 ( .A(n1241), .B(n1240), .Z(c[117]) );
  XOR U1454 ( .A(sreg[118]), .B(n1438), .Z(n1440) );
  NAND U1455 ( .A(n1252), .B(n1251), .Z(n1256) );
  NAND U1456 ( .A(n1254), .B(n1253), .Z(n1255) );
  NAND U1457 ( .A(n1256), .B(n1255), .Z(n1432) );
  XNOR U1458 ( .A(n1433), .B(n1432), .Z(n1435) );
  NAND U1459 ( .A(n1258), .B(n1257), .Z(n1262) );
  NAND U1460 ( .A(n1260), .B(n1259), .Z(n1261) );
  AND U1461 ( .A(n1262), .B(n1261), .Z(n1340) );
  NANDN U1462 ( .A(n1264), .B(n1263), .Z(n1268) );
  NANDN U1463 ( .A(n1266), .B(n1265), .Z(n1267) );
  AND U1464 ( .A(n1268), .B(n1267), .Z(n1339) );
  XNOR U1465 ( .A(n1340), .B(n1339), .Z(n1341) );
  NANDN U1466 ( .A(n1270), .B(n1269), .Z(n1274) );
  NAND U1467 ( .A(n1272), .B(n1271), .Z(n1273) );
  AND U1468 ( .A(n1274), .B(n1273), .Z(n1346) );
  NANDN U1469 ( .A(n1276), .B(n1275), .Z(n1280) );
  NANDN U1470 ( .A(n1278), .B(n1277), .Z(n1279) );
  AND U1471 ( .A(n1280), .B(n1279), .Z(n1353) );
  NANDN U1472 ( .A(n17067), .B(n1281), .Z(n1283) );
  XOR U1473 ( .A(b[3]), .B(a[20]), .Z(n1374) );
  NANDN U1474 ( .A(n17068), .B(n1374), .Z(n1282) );
  AND U1475 ( .A(n1283), .B(n1282), .Z(n1415) );
  NANDN U1476 ( .A(n18113), .B(n1284), .Z(n1286) );
  XOR U1477 ( .A(b[13]), .B(a[10]), .Z(n1388) );
  NANDN U1478 ( .A(n18229), .B(n1388), .Z(n1285) );
  NAND U1479 ( .A(n1286), .B(n1285), .Z(n1414) );
  XNOR U1480 ( .A(n1415), .B(n1414), .Z(n1417) );
  NOR U1481 ( .A(n1288), .B(n1287), .Z(n1416) );
  XOR U1482 ( .A(n1417), .B(n1416), .Z(n1352) );
  NAND U1483 ( .A(b[0]), .B(a[22]), .Z(n1289) );
  XNOR U1484 ( .A(b[1]), .B(n1289), .Z(n1291) );
  NANDN U1485 ( .A(b[0]), .B(a[21]), .Z(n1290) );
  NAND U1486 ( .A(n1291), .B(n1290), .Z(n1371) );
  XOR U1487 ( .A(b[22]), .B(b[21]), .Z(n19127) );
  IV U1488 ( .A(n19127), .Z(n19055) );
  ANDN U1489 ( .B(a[0]), .A(n19055), .Z(n1381) );
  IV U1490 ( .A(n18881), .Z(n18673) );
  NANDN U1491 ( .A(n18673), .B(n1292), .Z(n1294) );
  XOR U1492 ( .A(b[19]), .B(a[4]), .Z(n1385) );
  NANDN U1493 ( .A(n18758), .B(n1385), .Z(n1293) );
  AND U1494 ( .A(n1294), .B(n1293), .Z(n1369) );
  XOR U1495 ( .A(n1381), .B(n1369), .Z(n1370) );
  XNOR U1496 ( .A(n1371), .B(n1370), .Z(n1351) );
  XOR U1497 ( .A(n1352), .B(n1351), .Z(n1354) );
  XNOR U1498 ( .A(n1353), .B(n1354), .Z(n1345) );
  XNOR U1499 ( .A(n1346), .B(n1345), .Z(n1347) );
  NANDN U1500 ( .A(n17362), .B(n1295), .Z(n1297) );
  XOR U1501 ( .A(b[7]), .B(a[16]), .Z(n1405) );
  NANDN U1502 ( .A(n17522), .B(n1405), .Z(n1296) );
  AND U1503 ( .A(n1297), .B(n1296), .Z(n1428) );
  NANDN U1504 ( .A(n17072), .B(n1298), .Z(n1300) );
  XOR U1505 ( .A(b[5]), .B(a[18]), .Z(n1411) );
  NANDN U1506 ( .A(n17223), .B(n1411), .Z(n1299) );
  AND U1507 ( .A(n1300), .B(n1299), .Z(n1427) );
  NANDN U1508 ( .A(n18487), .B(n1301), .Z(n1303) );
  XOR U1509 ( .A(b[15]), .B(a[8]), .Z(n1377) );
  NANDN U1510 ( .A(n18311), .B(n1377), .Z(n1302) );
  NAND U1511 ( .A(n1303), .B(n1302), .Z(n1426) );
  XOR U1512 ( .A(n1427), .B(n1426), .Z(n1429) );
  XOR U1513 ( .A(n1428), .B(n1429), .Z(n1365) );
  NANDN U1514 ( .A(n18514), .B(n1304), .Z(n1306) );
  XOR U1515 ( .A(b[17]), .B(a[6]), .Z(n1382) );
  NANDN U1516 ( .A(n18585), .B(n1382), .Z(n1305) );
  AND U1517 ( .A(n1306), .B(n1305), .Z(n1422) );
  ANDN U1518 ( .B(n1307), .A(n18998), .Z(n18997) );
  IV U1519 ( .A(n18997), .Z(n18853) );
  NANDN U1520 ( .A(n18853), .B(n1308), .Z(n1310) );
  XOR U1521 ( .A(b[21]), .B(a[2]), .Z(n1402) );
  NANDN U1522 ( .A(n18926), .B(n1402), .Z(n1309) );
  AND U1523 ( .A(n1310), .B(n1309), .Z(n1421) );
  NANDN U1524 ( .A(n17613), .B(n1311), .Z(n1313) );
  XOR U1525 ( .A(b[9]), .B(a[14]), .Z(n1408) );
  NANDN U1526 ( .A(n17739), .B(n1408), .Z(n1312) );
  NAND U1527 ( .A(n1313), .B(n1312), .Z(n1420) );
  XOR U1528 ( .A(n1421), .B(n1420), .Z(n1423) );
  XOR U1529 ( .A(n1422), .B(n1423), .Z(n1364) );
  NANDN U1530 ( .A(n1314), .B(n18084), .Z(n1316) );
  XNOR U1531 ( .A(b[11]), .B(a[12]), .Z(n1391) );
  NANDN U1532 ( .A(n1391), .B(n18085), .Z(n1315) );
  AND U1533 ( .A(n1316), .B(n1315), .Z(n1363) );
  XOR U1534 ( .A(n1364), .B(n1363), .Z(n1366) );
  XOR U1535 ( .A(n1365), .B(n1366), .Z(n1360) );
  NANDN U1536 ( .A(n1318), .B(n1317), .Z(n1322) );
  NANDN U1537 ( .A(n1320), .B(n1319), .Z(n1321) );
  AND U1538 ( .A(n1322), .B(n1321), .Z(n1358) );
  NANDN U1539 ( .A(n1324), .B(n1323), .Z(n1328) );
  OR U1540 ( .A(n1326), .B(n1325), .Z(n1327) );
  NAND U1541 ( .A(n1328), .B(n1327), .Z(n1357) );
  XNOR U1542 ( .A(n1358), .B(n1357), .Z(n1359) );
  XOR U1543 ( .A(n1360), .B(n1359), .Z(n1348) );
  XOR U1544 ( .A(n1347), .B(n1348), .Z(n1342) );
  XNOR U1545 ( .A(n1341), .B(n1342), .Z(n1434) );
  XOR U1546 ( .A(n1435), .B(n1434), .Z(n1334) );
  XNOR U1547 ( .A(n1334), .B(n1333), .Z(n1335) );
  XNOR U1548 ( .A(n1336), .B(n1335), .Z(n1439) );
  XNOR U1549 ( .A(n1440), .B(n1439), .Z(c[118]) );
  NANDN U1550 ( .A(n1334), .B(n1333), .Z(n1338) );
  NANDN U1551 ( .A(n1336), .B(n1335), .Z(n1337) );
  AND U1552 ( .A(n1338), .B(n1337), .Z(n1451) );
  NANDN U1553 ( .A(n1340), .B(n1339), .Z(n1344) );
  NANDN U1554 ( .A(n1342), .B(n1341), .Z(n1343) );
  AND U1555 ( .A(n1344), .B(n1343), .Z(n1549) );
  NANDN U1556 ( .A(n1346), .B(n1345), .Z(n1350) );
  NANDN U1557 ( .A(n1348), .B(n1347), .Z(n1349) );
  AND U1558 ( .A(n1350), .B(n1349), .Z(n1457) );
  NANDN U1559 ( .A(n1352), .B(n1351), .Z(n1356) );
  OR U1560 ( .A(n1354), .B(n1353), .Z(n1355) );
  AND U1561 ( .A(n1356), .B(n1355), .Z(n1455) );
  NANDN U1562 ( .A(n1358), .B(n1357), .Z(n1362) );
  NANDN U1563 ( .A(n1360), .B(n1359), .Z(n1361) );
  AND U1564 ( .A(n1362), .B(n1361), .Z(n1454) );
  XNOR U1565 ( .A(n1455), .B(n1454), .Z(n1456) );
  XOR U1566 ( .A(n1457), .B(n1456), .Z(n1548) );
  NANDN U1567 ( .A(n1364), .B(n1363), .Z(n1368) );
  OR U1568 ( .A(n1366), .B(n1365), .Z(n1367) );
  AND U1569 ( .A(n1368), .B(n1367), .Z(n1460) );
  NANDN U1570 ( .A(n1369), .B(n1381), .Z(n1373) );
  OR U1571 ( .A(n1371), .B(n1370), .Z(n1372) );
  AND U1572 ( .A(n1373), .B(n1372), .Z(n1544) );
  NANDN U1573 ( .A(n17067), .B(n1374), .Z(n1376) );
  XOR U1574 ( .A(b[3]), .B(a[21]), .Z(n1489) );
  NANDN U1575 ( .A(n17068), .B(n1489), .Z(n1375) );
  AND U1576 ( .A(n1376), .B(n1375), .Z(n1495) );
  NANDN U1577 ( .A(n18487), .B(n1377), .Z(n1379) );
  XOR U1578 ( .A(b[15]), .B(a[9]), .Z(n1519) );
  NANDN U1579 ( .A(n18311), .B(n1519), .Z(n1378) );
  AND U1580 ( .A(n1379), .B(n1378), .Z(n1493) );
  NAND U1581 ( .A(b[21]), .B(b[22]), .Z(n1380) );
  AND U1582 ( .A(b[23]), .B(n1380), .Z(n19228) );
  ANDN U1583 ( .B(n19228), .A(n1381), .Z(n1492) );
  XNOR U1584 ( .A(n1493), .B(n1492), .Z(n1494) );
  XNOR U1585 ( .A(n1495), .B(n1494), .Z(n1541) );
  NANDN U1586 ( .A(n18514), .B(n1382), .Z(n1384) );
  XOR U1587 ( .A(b[17]), .B(a[7]), .Z(n1516) );
  NANDN U1588 ( .A(n18585), .B(n1516), .Z(n1383) );
  AND U1589 ( .A(n1384), .B(n1383), .Z(n1481) );
  NANDN U1590 ( .A(n18673), .B(n1385), .Z(n1387) );
  XOR U1591 ( .A(b[19]), .B(a[5]), .Z(n1525) );
  NANDN U1592 ( .A(n18758), .B(n1525), .Z(n1386) );
  AND U1593 ( .A(n1387), .B(n1386), .Z(n1479) );
  NANDN U1594 ( .A(n18113), .B(n1388), .Z(n1390) );
  XOR U1595 ( .A(b[13]), .B(a[11]), .Z(n1486) );
  NANDN U1596 ( .A(n18229), .B(n1486), .Z(n1389) );
  NAND U1597 ( .A(n1390), .B(n1389), .Z(n1478) );
  XNOR U1598 ( .A(n1479), .B(n1478), .Z(n1480) );
  XOR U1599 ( .A(n1481), .B(n1480), .Z(n1542) );
  XNOR U1600 ( .A(n1541), .B(n1542), .Z(n1543) );
  XOR U1601 ( .A(n1544), .B(n1543), .Z(n1461) );
  XNOR U1602 ( .A(n1460), .B(n1461), .Z(n1462) );
  NANDN U1603 ( .A(n1391), .B(n18084), .Z(n1393) );
  XOR U1604 ( .A(b[11]), .B(a[13]), .Z(n1522) );
  NANDN U1605 ( .A(n18025), .B(n1522), .Z(n1392) );
  NAND U1606 ( .A(n1393), .B(n1392), .Z(n1472) );
  NAND U1607 ( .A(b[0]), .B(a[23]), .Z(n1394) );
  XNOR U1608 ( .A(b[1]), .B(n1394), .Z(n1396) );
  NANDN U1609 ( .A(b[0]), .B(a[22]), .Z(n1395) );
  NAND U1610 ( .A(n1396), .B(n1395), .Z(n1473) );
  XNOR U1611 ( .A(n1472), .B(n1473), .Z(n1474) );
  XOR U1612 ( .A(b[23]), .B(a[0]), .Z(n1399) );
  XOR U1613 ( .A(b[23]), .B(b[21]), .Z(n1397) );
  XOR U1614 ( .A(b[23]), .B(b[22]), .Z(n1528) );
  AND U1615 ( .A(n1397), .B(n1528), .Z(n1398) );
  NAND U1616 ( .A(n1399), .B(n1398), .Z(n1401) );
  XOR U1617 ( .A(b[23]), .B(a[1]), .Z(n1529) );
  NANDN U1618 ( .A(n19055), .B(n1529), .Z(n1400) );
  AND U1619 ( .A(n1401), .B(n1400), .Z(n1484) );
  NANDN U1620 ( .A(n18853), .B(n1402), .Z(n1404) );
  XOR U1621 ( .A(b[21]), .B(a[3]), .Z(n1507) );
  NANDN U1622 ( .A(n18926), .B(n1507), .Z(n1403) );
  NAND U1623 ( .A(n1404), .B(n1403), .Z(n1485) );
  XOR U1624 ( .A(n1484), .B(n1485), .Z(n1475) );
  XNOR U1625 ( .A(n1474), .B(n1475), .Z(n1536) );
  NANDN U1626 ( .A(n17362), .B(n1405), .Z(n1407) );
  XOR U1627 ( .A(b[7]), .B(a[17]), .Z(n1510) );
  NANDN U1628 ( .A(n17522), .B(n1510), .Z(n1406) );
  AND U1629 ( .A(n1407), .B(n1406), .Z(n1500) );
  NANDN U1630 ( .A(n17613), .B(n1408), .Z(n1410) );
  XOR U1631 ( .A(b[9]), .B(a[15]), .Z(n1532) );
  NANDN U1632 ( .A(n17739), .B(n1532), .Z(n1409) );
  AND U1633 ( .A(n1410), .B(n1409), .Z(n1499) );
  NANDN U1634 ( .A(n17072), .B(n1411), .Z(n1413) );
  XOR U1635 ( .A(b[5]), .B(a[19]), .Z(n1513) );
  NANDN U1636 ( .A(n17223), .B(n1513), .Z(n1412) );
  NAND U1637 ( .A(n1413), .B(n1412), .Z(n1498) );
  XOR U1638 ( .A(n1499), .B(n1498), .Z(n1501) );
  XOR U1639 ( .A(n1500), .B(n1501), .Z(n1535) );
  XOR U1640 ( .A(n1536), .B(n1535), .Z(n1538) );
  NANDN U1641 ( .A(n1415), .B(n1414), .Z(n1419) );
  NAND U1642 ( .A(n1417), .B(n1416), .Z(n1418) );
  NAND U1643 ( .A(n1419), .B(n1418), .Z(n1537) );
  XOR U1644 ( .A(n1538), .B(n1537), .Z(n1468) );
  NANDN U1645 ( .A(n1421), .B(n1420), .Z(n1425) );
  OR U1646 ( .A(n1423), .B(n1422), .Z(n1424) );
  AND U1647 ( .A(n1425), .B(n1424), .Z(n1467) );
  NANDN U1648 ( .A(n1427), .B(n1426), .Z(n1431) );
  OR U1649 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U1650 ( .A(n1431), .B(n1430), .Z(n1466) );
  XOR U1651 ( .A(n1467), .B(n1466), .Z(n1469) );
  XOR U1652 ( .A(n1468), .B(n1469), .Z(n1463) );
  XNOR U1653 ( .A(n1462), .B(n1463), .Z(n1547) );
  XOR U1654 ( .A(n1548), .B(n1547), .Z(n1550) );
  XOR U1655 ( .A(n1549), .B(n1550), .Z(n1449) );
  NANDN U1656 ( .A(n1433), .B(n1432), .Z(n1437) );
  NAND U1657 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U1658 ( .A(n1437), .B(n1436), .Z(n1448) );
  XNOR U1659 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U1660 ( .A(n1451), .B(n1450), .Z(n1443) );
  XNOR U1661 ( .A(sreg[119]), .B(n1443), .Z(n1445) );
  OR U1662 ( .A(sreg[118]), .B(n1438), .Z(n1442) );
  NAND U1663 ( .A(n1440), .B(n1439), .Z(n1441) );
  NAND U1664 ( .A(n1442), .B(n1441), .Z(n1444) );
  XNOR U1665 ( .A(n1445), .B(n1444), .Z(c[119]) );
  NANDN U1666 ( .A(sreg[119]), .B(n1443), .Z(n1447) );
  NAND U1667 ( .A(n1445), .B(n1444), .Z(n1446) );
  NAND U1668 ( .A(n1447), .B(n1446), .Z(n1662) );
  XNOR U1669 ( .A(sreg[120]), .B(n1662), .Z(n1664) );
  NANDN U1670 ( .A(n1449), .B(n1448), .Z(n1453) );
  NANDN U1671 ( .A(n1451), .B(n1450), .Z(n1452) );
  AND U1672 ( .A(n1453), .B(n1452), .Z(n1556) );
  NANDN U1673 ( .A(n1455), .B(n1454), .Z(n1459) );
  NAND U1674 ( .A(n1457), .B(n1456), .Z(n1458) );
  AND U1675 ( .A(n1459), .B(n1458), .Z(n1562) );
  NANDN U1676 ( .A(n1461), .B(n1460), .Z(n1465) );
  NANDN U1677 ( .A(n1463), .B(n1462), .Z(n1464) );
  AND U1678 ( .A(n1465), .B(n1464), .Z(n1559) );
  NANDN U1679 ( .A(n1467), .B(n1466), .Z(n1471) );
  NANDN U1680 ( .A(n1469), .B(n1468), .Z(n1470) );
  AND U1681 ( .A(n1471), .B(n1470), .Z(n1658) );
  NANDN U1682 ( .A(n1473), .B(n1472), .Z(n1477) );
  NANDN U1683 ( .A(n1475), .B(n1474), .Z(n1476) );
  AND U1684 ( .A(n1477), .B(n1476), .Z(n1578) );
  NANDN U1685 ( .A(n1479), .B(n1478), .Z(n1483) );
  NANDN U1686 ( .A(n1481), .B(n1480), .Z(n1482) );
  AND U1687 ( .A(n1483), .B(n1482), .Z(n1575) );
  ANDN U1688 ( .B(n1485), .A(n1484), .Z(n1616) );
  NAND U1689 ( .A(n18347), .B(n1486), .Z(n1488) );
  XNOR U1690 ( .A(b[13]), .B(a[12]), .Z(n1602) );
  NANDN U1691 ( .A(n1602), .B(n18345), .Z(n1487) );
  AND U1692 ( .A(n1488), .B(n1487), .Z(n1613) );
  NAND U1693 ( .A(n2664), .B(n1489), .Z(n1491) );
  XNOR U1694 ( .A(b[3]), .B(a[22]), .Z(n1605) );
  NANDN U1695 ( .A(n1605), .B(n2512), .Z(n1490) );
  NAND U1696 ( .A(n1491), .B(n1490), .Z(n1614) );
  XNOR U1697 ( .A(n1613), .B(n1614), .Z(n1615) );
  XOR U1698 ( .A(n1616), .B(n1615), .Z(n1576) );
  XNOR U1699 ( .A(n1575), .B(n1576), .Z(n1577) );
  XOR U1700 ( .A(n1578), .B(n1577), .Z(n1657) );
  NANDN U1701 ( .A(n1493), .B(n1492), .Z(n1497) );
  NANDN U1702 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U1703 ( .A(n1497), .B(n1496), .Z(n1572) );
  NANDN U1704 ( .A(n1499), .B(n1498), .Z(n1503) );
  OR U1705 ( .A(n1501), .B(n1500), .Z(n1502) );
  NAND U1706 ( .A(n1503), .B(n1502), .Z(n1571) );
  XNOR U1707 ( .A(n1572), .B(n1571), .Z(n1574) );
  NAND U1708 ( .A(b[0]), .B(a[24]), .Z(n1504) );
  XNOR U1709 ( .A(b[1]), .B(n1504), .Z(n1506) );
  NANDN U1710 ( .A(b[0]), .B(a[23]), .Z(n1505) );
  NAND U1711 ( .A(n1506), .B(n1505), .Z(n1589) );
  XOR U1712 ( .A(b[24]), .B(b[23]), .Z(n19224) );
  IV U1713 ( .A(n19224), .Z(n19179) );
  ANDN U1714 ( .B(a[0]), .A(n19179), .Z(n1612) );
  NANDN U1715 ( .A(n18853), .B(n1507), .Z(n1509) );
  XOR U1716 ( .A(b[21]), .B(a[4]), .Z(n1647) );
  NANDN U1717 ( .A(n18926), .B(n1647), .Z(n1508) );
  AND U1718 ( .A(n1509), .B(n1508), .Z(n1587) );
  XNOR U1719 ( .A(n1612), .B(n1587), .Z(n1588) );
  XNOR U1720 ( .A(n1589), .B(n1588), .Z(n1581) );
  NANDN U1721 ( .A(n17362), .B(n1510), .Z(n1512) );
  XOR U1722 ( .A(b[7]), .B(a[18]), .Z(n1635) );
  NANDN U1723 ( .A(n17522), .B(n1635), .Z(n1511) );
  AND U1724 ( .A(n1512), .B(n1511), .Z(n1632) );
  NANDN U1725 ( .A(n17072), .B(n1513), .Z(n1515) );
  XOR U1726 ( .A(b[5]), .B(a[20]), .Z(n1638) );
  NANDN U1727 ( .A(n17223), .B(n1638), .Z(n1514) );
  AND U1728 ( .A(n1515), .B(n1514), .Z(n1630) );
  NANDN U1729 ( .A(n18514), .B(n1516), .Z(n1518) );
  XOR U1730 ( .A(b[17]), .B(a[8]), .Z(n1641) );
  NANDN U1731 ( .A(n18585), .B(n1641), .Z(n1517) );
  NAND U1732 ( .A(n1518), .B(n1517), .Z(n1629) );
  XNOR U1733 ( .A(n1630), .B(n1629), .Z(n1631) );
  XOR U1734 ( .A(n1632), .B(n1631), .Z(n1582) );
  XNOR U1735 ( .A(n1581), .B(n1582), .Z(n1583) );
  NANDN U1736 ( .A(n18487), .B(n1519), .Z(n1521) );
  XOR U1737 ( .A(b[15]), .B(a[10]), .Z(n1608) );
  NANDN U1738 ( .A(n18311), .B(n1608), .Z(n1520) );
  AND U1739 ( .A(n1521), .B(n1520), .Z(n1626) );
  NANDN U1740 ( .A(n17888), .B(n1522), .Z(n1524) );
  XOR U1741 ( .A(b[11]), .B(a[14]), .Z(n1653) );
  NANDN U1742 ( .A(n18025), .B(n1653), .Z(n1523) );
  NAND U1743 ( .A(n1524), .B(n1523), .Z(n1625) );
  XNOR U1744 ( .A(n1626), .B(n1625), .Z(n1628) );
  NAND U1745 ( .A(n18881), .B(n1525), .Z(n1527) );
  XNOR U1746 ( .A(b[19]), .B(a[6]), .Z(n1644) );
  NANDN U1747 ( .A(n1644), .B(n18882), .Z(n1526) );
  NAND U1748 ( .A(n1527), .B(n1526), .Z(n1621) );
  ANDN U1749 ( .B(n1528), .A(n19127), .Z(n19126) );
  NAND U1750 ( .A(n19126), .B(n1529), .Z(n1531) );
  XNOR U1751 ( .A(b[23]), .B(a[2]), .Z(n1592) );
  NANDN U1752 ( .A(n1592), .B(n19127), .Z(n1530) );
  NAND U1753 ( .A(n1531), .B(n1530), .Z(n1620) );
  NANDN U1754 ( .A(n17613), .B(n1532), .Z(n1534) );
  XOR U1755 ( .A(b[9]), .B(a[16]), .Z(n1650) );
  NANDN U1756 ( .A(n17739), .B(n1650), .Z(n1533) );
  NAND U1757 ( .A(n1534), .B(n1533), .Z(n1619) );
  XOR U1758 ( .A(n1620), .B(n1619), .Z(n1622) );
  XOR U1759 ( .A(n1621), .B(n1622), .Z(n1627) );
  XNOR U1760 ( .A(n1628), .B(n1627), .Z(n1584) );
  XNOR U1761 ( .A(n1583), .B(n1584), .Z(n1573) );
  XOR U1762 ( .A(n1574), .B(n1573), .Z(n1656) );
  XOR U1763 ( .A(n1657), .B(n1656), .Z(n1659) );
  XOR U1764 ( .A(n1658), .B(n1659), .Z(n1568) );
  NAND U1765 ( .A(n1536), .B(n1535), .Z(n1540) );
  NAND U1766 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1767 ( .A(n1540), .B(n1539), .Z(n1565) );
  NANDN U1768 ( .A(n1542), .B(n1541), .Z(n1546) );
  NANDN U1769 ( .A(n1544), .B(n1543), .Z(n1545) );
  NAND U1770 ( .A(n1546), .B(n1545), .Z(n1566) );
  XNOR U1771 ( .A(n1565), .B(n1566), .Z(n1567) );
  XOR U1772 ( .A(n1568), .B(n1567), .Z(n1560) );
  XNOR U1773 ( .A(n1559), .B(n1560), .Z(n1561) );
  XNOR U1774 ( .A(n1562), .B(n1561), .Z(n1553) );
  NANDN U1775 ( .A(n1548), .B(n1547), .Z(n1552) );
  OR U1776 ( .A(n1550), .B(n1549), .Z(n1551) );
  NAND U1777 ( .A(n1552), .B(n1551), .Z(n1554) );
  XNOR U1778 ( .A(n1553), .B(n1554), .Z(n1555) );
  XNOR U1779 ( .A(n1556), .B(n1555), .Z(n1663) );
  XNOR U1780 ( .A(n1664), .B(n1663), .Z(c[120]) );
  NANDN U1781 ( .A(n1554), .B(n1553), .Z(n1558) );
  NANDN U1782 ( .A(n1556), .B(n1555), .Z(n1557) );
  AND U1783 ( .A(n1558), .B(n1557), .Z(n1675) );
  NANDN U1784 ( .A(n1560), .B(n1559), .Z(n1564) );
  NANDN U1785 ( .A(n1562), .B(n1561), .Z(n1563) );
  AND U1786 ( .A(n1564), .B(n1563), .Z(n1673) );
  NANDN U1787 ( .A(n1566), .B(n1565), .Z(n1570) );
  NANDN U1788 ( .A(n1568), .B(n1567), .Z(n1569) );
  AND U1789 ( .A(n1570), .B(n1569), .Z(n1681) );
  NANDN U1790 ( .A(n1576), .B(n1575), .Z(n1580) );
  NAND U1791 ( .A(n1578), .B(n1577), .Z(n1579) );
  AND U1792 ( .A(n1580), .B(n1579), .Z(n1690) );
  XNOR U1793 ( .A(n1691), .B(n1690), .Z(n1693) );
  NANDN U1794 ( .A(n1582), .B(n1581), .Z(n1586) );
  NANDN U1795 ( .A(n1584), .B(n1583), .Z(n1585) );
  AND U1796 ( .A(n1586), .B(n1585), .Z(n1685) );
  NANDN U1797 ( .A(n1587), .B(n1612), .Z(n1591) );
  NANDN U1798 ( .A(n1589), .B(n1588), .Z(n1590) );
  AND U1799 ( .A(n1591), .B(n1590), .Z(n1698) );
  NANDN U1800 ( .A(n1592), .B(n19126), .Z(n1594) );
  XOR U1801 ( .A(b[23]), .B(a[3]), .Z(n1733) );
  NANDN U1802 ( .A(n19055), .B(n1733), .Z(n1593) );
  AND U1803 ( .A(n1594), .B(n1593), .Z(n1751) );
  XOR U1804 ( .A(b[25]), .B(b[24]), .Z(n1711) );
  XOR U1805 ( .A(b[25]), .B(a[0]), .Z(n1595) );
  NAND U1806 ( .A(n1711), .B(n1595), .Z(n1596) );
  OR U1807 ( .A(n1596), .B(n19224), .Z(n1598) );
  XOR U1808 ( .A(b[25]), .B(a[1]), .Z(n1712) );
  NAND U1809 ( .A(n19224), .B(n1712), .Z(n1597) );
  AND U1810 ( .A(n1598), .B(n1597), .Z(n1752) );
  XOR U1811 ( .A(n1751), .B(n1752), .Z(n1704) );
  NAND U1812 ( .A(b[0]), .B(a[25]), .Z(n1599) );
  XNOR U1813 ( .A(b[1]), .B(n1599), .Z(n1601) );
  NANDN U1814 ( .A(b[0]), .B(a[24]), .Z(n1600) );
  NAND U1815 ( .A(n1601), .B(n1600), .Z(n1702) );
  NANDN U1816 ( .A(n1602), .B(n18347), .Z(n1604) );
  XNOR U1817 ( .A(b[13]), .B(a[13]), .Z(n1759) );
  NANDN U1818 ( .A(n1759), .B(n18345), .Z(n1603) );
  NAND U1819 ( .A(n1604), .B(n1603), .Z(n1703) );
  XOR U1820 ( .A(n1702), .B(n1703), .Z(n1705) );
  XOR U1821 ( .A(n1704), .B(n1705), .Z(n1697) );
  NANDN U1822 ( .A(n1605), .B(n2664), .Z(n1607) );
  XOR U1823 ( .A(b[3]), .B(a[23]), .Z(n1756) );
  NANDN U1824 ( .A(n17068), .B(n1756), .Z(n1606) );
  AND U1825 ( .A(n1607), .B(n1606), .Z(n1721) );
  NANDN U1826 ( .A(n18487), .B(n1608), .Z(n1610) );
  XOR U1827 ( .A(b[15]), .B(a[11]), .Z(n1753) );
  NANDN U1828 ( .A(n18311), .B(n1753), .Z(n1609) );
  AND U1829 ( .A(n1610), .B(n1609), .Z(n1719) );
  NAND U1830 ( .A(b[23]), .B(b[24]), .Z(n1611) );
  AND U1831 ( .A(b[25]), .B(n1611), .Z(n19314) );
  ANDN U1832 ( .B(n19314), .A(n1612), .Z(n1718) );
  XNOR U1833 ( .A(n1719), .B(n1718), .Z(n1720) );
  XNOR U1834 ( .A(n1721), .B(n1720), .Z(n1696) );
  XOR U1835 ( .A(n1697), .B(n1696), .Z(n1699) );
  XOR U1836 ( .A(n1698), .B(n1699), .Z(n1776) );
  NANDN U1837 ( .A(n1614), .B(n1613), .Z(n1618) );
  NANDN U1838 ( .A(n1616), .B(n1615), .Z(n1617) );
  AND U1839 ( .A(n1618), .B(n1617), .Z(n1775) );
  NAND U1840 ( .A(n1620), .B(n1619), .Z(n1624) );
  NAND U1841 ( .A(n1622), .B(n1621), .Z(n1623) );
  AND U1842 ( .A(n1624), .B(n1623), .Z(n1774) );
  XOR U1843 ( .A(n1775), .B(n1774), .Z(n1777) );
  XNOR U1844 ( .A(n1776), .B(n1777), .Z(n1684) );
  XNOR U1845 ( .A(n1685), .B(n1684), .Z(n1686) );
  NANDN U1846 ( .A(n1630), .B(n1629), .Z(n1634) );
  NANDN U1847 ( .A(n1632), .B(n1631), .Z(n1633) );
  AND U1848 ( .A(n1634), .B(n1633), .Z(n1781) );
  NANDN U1849 ( .A(n17362), .B(n1635), .Z(n1637) );
  XOR U1850 ( .A(b[7]), .B(a[19]), .Z(n1742) );
  NANDN U1851 ( .A(n17522), .B(n1742), .Z(n1636) );
  AND U1852 ( .A(n1637), .B(n1636), .Z(n1747) );
  NANDN U1853 ( .A(n17072), .B(n1638), .Z(n1640) );
  XOR U1854 ( .A(b[5]), .B(a[21]), .Z(n1765) );
  NANDN U1855 ( .A(n17223), .B(n1765), .Z(n1639) );
  AND U1856 ( .A(n1640), .B(n1639), .Z(n1746) );
  NANDN U1857 ( .A(n18514), .B(n1641), .Z(n1643) );
  XOR U1858 ( .A(b[17]), .B(a[9]), .Z(n1715) );
  NANDN U1859 ( .A(n18585), .B(n1715), .Z(n1642) );
  NAND U1860 ( .A(n1643), .B(n1642), .Z(n1745) );
  XOR U1861 ( .A(n1746), .B(n1745), .Z(n1748) );
  XOR U1862 ( .A(n1747), .B(n1748), .Z(n1770) );
  NANDN U1863 ( .A(n1644), .B(n18881), .Z(n1646) );
  XOR U1864 ( .A(b[19]), .B(a[7]), .Z(n1762) );
  NANDN U1865 ( .A(n18758), .B(n1762), .Z(n1645) );
  AND U1866 ( .A(n1646), .B(n1645), .Z(n1726) );
  NANDN U1867 ( .A(n18853), .B(n1647), .Z(n1649) );
  XOR U1868 ( .A(b[21]), .B(a[5]), .Z(n1708) );
  NANDN U1869 ( .A(n18926), .B(n1708), .Z(n1648) );
  AND U1870 ( .A(n1649), .B(n1648), .Z(n1725) );
  NANDN U1871 ( .A(n17613), .B(n1650), .Z(n1652) );
  XOR U1872 ( .A(b[9]), .B(a[17]), .Z(n1736) );
  NANDN U1873 ( .A(n17739), .B(n1736), .Z(n1651) );
  NAND U1874 ( .A(n1652), .B(n1651), .Z(n1724) );
  XOR U1875 ( .A(n1725), .B(n1724), .Z(n1727) );
  XOR U1876 ( .A(n1726), .B(n1727), .Z(n1769) );
  NAND U1877 ( .A(n18084), .B(n1653), .Z(n1655) );
  XNOR U1878 ( .A(b[11]), .B(a[15]), .Z(n1739) );
  NANDN U1879 ( .A(n1739), .B(n18085), .Z(n1654) );
  AND U1880 ( .A(n1655), .B(n1654), .Z(n1768) );
  XOR U1881 ( .A(n1769), .B(n1768), .Z(n1771) );
  XNOR U1882 ( .A(n1770), .B(n1771), .Z(n1780) );
  XNOR U1883 ( .A(n1781), .B(n1780), .Z(n1782) );
  XOR U1884 ( .A(n1783), .B(n1782), .Z(n1687) );
  XNOR U1885 ( .A(n1686), .B(n1687), .Z(n1692) );
  XOR U1886 ( .A(n1693), .B(n1692), .Z(n1679) );
  NANDN U1887 ( .A(n1657), .B(n1656), .Z(n1661) );
  OR U1888 ( .A(n1659), .B(n1658), .Z(n1660) );
  AND U1889 ( .A(n1661), .B(n1660), .Z(n1678) );
  XNOR U1890 ( .A(n1679), .B(n1678), .Z(n1680) );
  XNOR U1891 ( .A(n1681), .B(n1680), .Z(n1672) );
  XNOR U1892 ( .A(n1673), .B(n1672), .Z(n1674) );
  XNOR U1893 ( .A(n1675), .B(n1674), .Z(n1667) );
  XNOR U1894 ( .A(sreg[121]), .B(n1667), .Z(n1669) );
  NANDN U1895 ( .A(sreg[120]), .B(n1662), .Z(n1666) );
  NAND U1896 ( .A(n1664), .B(n1663), .Z(n1665) );
  NAND U1897 ( .A(n1666), .B(n1665), .Z(n1668) );
  XNOR U1898 ( .A(n1669), .B(n1668), .Z(c[121]) );
  NANDN U1899 ( .A(sreg[121]), .B(n1667), .Z(n1671) );
  NAND U1900 ( .A(n1669), .B(n1668), .Z(n1670) );
  AND U1901 ( .A(n1671), .B(n1670), .Z(n1787) );
  NANDN U1902 ( .A(n1673), .B(n1672), .Z(n1677) );
  NANDN U1903 ( .A(n1675), .B(n1674), .Z(n1676) );
  AND U1904 ( .A(n1677), .B(n1676), .Z(n1792) );
  NANDN U1905 ( .A(n1679), .B(n1678), .Z(n1683) );
  NANDN U1906 ( .A(n1681), .B(n1680), .Z(n1682) );
  AND U1907 ( .A(n1683), .B(n1682), .Z(n1790) );
  NANDN U1908 ( .A(n1685), .B(n1684), .Z(n1689) );
  NANDN U1909 ( .A(n1687), .B(n1686), .Z(n1688) );
  AND U1910 ( .A(n1689), .B(n1688), .Z(n1795) );
  NANDN U1911 ( .A(n1691), .B(n1690), .Z(n1695) );
  NAND U1912 ( .A(n1693), .B(n1692), .Z(n1694) );
  NAND U1913 ( .A(n1695), .B(n1694), .Z(n1796) );
  XNOR U1914 ( .A(n1795), .B(n1796), .Z(n1797) );
  NANDN U1915 ( .A(n1697), .B(n1696), .Z(n1701) );
  OR U1916 ( .A(n1699), .B(n1698), .Z(n1700) );
  AND U1917 ( .A(n1701), .B(n1700), .Z(n1814) );
  NANDN U1918 ( .A(n1703), .B(n1702), .Z(n1707) );
  OR U1919 ( .A(n1705), .B(n1704), .Z(n1706) );
  AND U1920 ( .A(n1707), .B(n1706), .Z(n1894) );
  NANDN U1921 ( .A(n18853), .B(n1708), .Z(n1710) );
  XOR U1922 ( .A(b[21]), .B(a[6]), .Z(n1878) );
  NANDN U1923 ( .A(n18926), .B(n1878), .Z(n1709) );
  AND U1924 ( .A(n1710), .B(n1709), .Z(n1849) );
  ANDN U1925 ( .B(n1711), .A(n19224), .Z(n19223) );
  IV U1926 ( .A(n19223), .Z(n19116) );
  NANDN U1927 ( .A(n19116), .B(n1712), .Z(n1714) );
  XOR U1928 ( .A(b[25]), .B(a[2]), .Z(n1829) );
  NANDN U1929 ( .A(n19179), .B(n1829), .Z(n1713) );
  AND U1930 ( .A(n1714), .B(n1713), .Z(n1848) );
  NANDN U1931 ( .A(n18514), .B(n1715), .Z(n1717) );
  XOR U1932 ( .A(b[17]), .B(a[10]), .Z(n1875) );
  NANDN U1933 ( .A(n18585), .B(n1875), .Z(n1716) );
  NAND U1934 ( .A(n1717), .B(n1716), .Z(n1847) );
  XOR U1935 ( .A(n1848), .B(n1847), .Z(n1850) );
  XNOR U1936 ( .A(n1849), .B(n1850), .Z(n1893) );
  XNOR U1937 ( .A(n1894), .B(n1893), .Z(n1896) );
  NANDN U1938 ( .A(n1719), .B(n1718), .Z(n1723) );
  NANDN U1939 ( .A(n1721), .B(n1720), .Z(n1722) );
  AND U1940 ( .A(n1723), .B(n1722), .Z(n1895) );
  XNOR U1941 ( .A(n1896), .B(n1895), .Z(n1813) );
  XNOR U1942 ( .A(n1814), .B(n1813), .Z(n1816) );
  NANDN U1943 ( .A(n1725), .B(n1724), .Z(n1729) );
  OR U1944 ( .A(n1727), .B(n1726), .Z(n1728) );
  AND U1945 ( .A(n1729), .B(n1728), .Z(n1902) );
  NAND U1946 ( .A(b[0]), .B(a[26]), .Z(n1730) );
  XNOR U1947 ( .A(b[1]), .B(n1730), .Z(n1732) );
  NANDN U1948 ( .A(b[0]), .B(a[25]), .Z(n1731) );
  NAND U1949 ( .A(n1732), .B(n1731), .Z(n1861) );
  XOR U1950 ( .A(b[26]), .B(b[25]), .Z(n19322) );
  IV U1951 ( .A(n19322), .Z(n19277) );
  ANDN U1952 ( .B(a[0]), .A(n19277), .Z(n1871) );
  IV U1953 ( .A(n19126), .Z(n19005) );
  NANDN U1954 ( .A(n19005), .B(n1733), .Z(n1735) );
  XOR U1955 ( .A(b[23]), .B(a[4]), .Z(n1881) );
  NANDN U1956 ( .A(n19055), .B(n1881), .Z(n1734) );
  AND U1957 ( .A(n1735), .B(n1734), .Z(n1859) );
  XNOR U1958 ( .A(n1871), .B(n1859), .Z(n1860) );
  XNOR U1959 ( .A(n1861), .B(n1860), .Z(n1899) );
  NANDN U1960 ( .A(n17613), .B(n1736), .Z(n1738) );
  XOR U1961 ( .A(b[9]), .B(a[18]), .Z(n1884) );
  NANDN U1962 ( .A(n17739), .B(n1884), .Z(n1737) );
  AND U1963 ( .A(n1738), .B(n1737), .Z(n1856) );
  NANDN U1964 ( .A(n1739), .B(n18084), .Z(n1741) );
  XOR U1965 ( .A(b[11]), .B(a[16]), .Z(n1872) );
  NANDN U1966 ( .A(n18025), .B(n1872), .Z(n1740) );
  AND U1967 ( .A(n1741), .B(n1740), .Z(n1854) );
  NANDN U1968 ( .A(n17362), .B(n1742), .Z(n1744) );
  XOR U1969 ( .A(b[7]), .B(a[20]), .Z(n1832) );
  NANDN U1970 ( .A(n17522), .B(n1832), .Z(n1743) );
  NAND U1971 ( .A(n1744), .B(n1743), .Z(n1853) );
  XNOR U1972 ( .A(n1854), .B(n1853), .Z(n1855) );
  XOR U1973 ( .A(n1856), .B(n1855), .Z(n1900) );
  XNOR U1974 ( .A(n1899), .B(n1900), .Z(n1901) );
  XNOR U1975 ( .A(n1902), .B(n1901), .Z(n1808) );
  NANDN U1976 ( .A(n1746), .B(n1745), .Z(n1750) );
  OR U1977 ( .A(n1748), .B(n1747), .Z(n1749) );
  AND U1978 ( .A(n1750), .B(n1749), .Z(n1907) );
  NOR U1979 ( .A(n1752), .B(n1751), .Z(n1843) );
  NAND U1980 ( .A(n18439), .B(n1753), .Z(n1755) );
  XNOR U1981 ( .A(b[15]), .B(a[12]), .Z(n1867) );
  NANDN U1982 ( .A(n1867), .B(n18486), .Z(n1754) );
  AND U1983 ( .A(n1755), .B(n1754), .Z(n1841) );
  NAND U1984 ( .A(n2664), .B(n1756), .Z(n1758) );
  XNOR U1985 ( .A(b[3]), .B(a[24]), .Z(n1864) );
  NANDN U1986 ( .A(n1864), .B(n2512), .Z(n1757) );
  NAND U1987 ( .A(n1758), .B(n1757), .Z(n1842) );
  XOR U1988 ( .A(n1841), .B(n1842), .Z(n1844) );
  XOR U1989 ( .A(n1843), .B(n1844), .Z(n1906) );
  NANDN U1990 ( .A(n1759), .B(n18347), .Z(n1761) );
  XOR U1991 ( .A(b[13]), .B(a[14]), .Z(n1822) );
  NANDN U1992 ( .A(n18229), .B(n1822), .Z(n1760) );
  AND U1993 ( .A(n1761), .B(n1760), .Z(n1890) );
  NANDN U1994 ( .A(n18673), .B(n1762), .Z(n1764) );
  XOR U1995 ( .A(b[19]), .B(a[8]), .Z(n1838) );
  NANDN U1996 ( .A(n18758), .B(n1838), .Z(n1763) );
  AND U1997 ( .A(n1764), .B(n1763), .Z(n1888) );
  NANDN U1998 ( .A(n17072), .B(n1765), .Z(n1767) );
  XOR U1999 ( .A(b[5]), .B(a[22]), .Z(n1835) );
  NANDN U2000 ( .A(n17223), .B(n1835), .Z(n1766) );
  NAND U2001 ( .A(n1767), .B(n1766), .Z(n1887) );
  XNOR U2002 ( .A(n1888), .B(n1887), .Z(n1889) );
  XNOR U2003 ( .A(n1890), .B(n1889), .Z(n1905) );
  XOR U2004 ( .A(n1906), .B(n1905), .Z(n1908) );
  XOR U2005 ( .A(n1907), .B(n1908), .Z(n1807) );
  XOR U2006 ( .A(n1808), .B(n1807), .Z(n1810) );
  NANDN U2007 ( .A(n1769), .B(n1768), .Z(n1773) );
  OR U2008 ( .A(n1771), .B(n1770), .Z(n1772) );
  AND U2009 ( .A(n1773), .B(n1772), .Z(n1809) );
  XOR U2010 ( .A(n1810), .B(n1809), .Z(n1815) );
  XOR U2011 ( .A(n1816), .B(n1815), .Z(n1804) );
  NANDN U2012 ( .A(n1775), .B(n1774), .Z(n1779) );
  OR U2013 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U2014 ( .A(n1779), .B(n1778), .Z(n1802) );
  NANDN U2015 ( .A(n1781), .B(n1780), .Z(n1785) );
  NANDN U2016 ( .A(n1783), .B(n1782), .Z(n1784) );
  AND U2017 ( .A(n1785), .B(n1784), .Z(n1801) );
  XNOR U2018 ( .A(n1802), .B(n1801), .Z(n1803) );
  XOR U2019 ( .A(n1804), .B(n1803), .Z(n1798) );
  XNOR U2020 ( .A(n1797), .B(n1798), .Z(n1789) );
  XNOR U2021 ( .A(n1790), .B(n1789), .Z(n1791) );
  XNOR U2022 ( .A(n1792), .B(n1791), .Z(n1788) );
  XNOR U2023 ( .A(sreg[122]), .B(n1788), .Z(n1786) );
  XOR U2024 ( .A(n1787), .B(n1786), .Z(c[122]) );
  NANDN U2025 ( .A(n1790), .B(n1789), .Z(n1794) );
  NANDN U2026 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U2027 ( .A(n1794), .B(n1793), .Z(n1919) );
  NANDN U2028 ( .A(n1796), .B(n1795), .Z(n1800) );
  NANDN U2029 ( .A(n1798), .B(n1797), .Z(n1799) );
  AND U2030 ( .A(n1800), .B(n1799), .Z(n1917) );
  NANDN U2031 ( .A(n1802), .B(n1801), .Z(n1806) );
  NANDN U2032 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U2033 ( .A(n1806), .B(n1805), .Z(n1925) );
  NAND U2034 ( .A(n1808), .B(n1807), .Z(n1812) );
  NAND U2035 ( .A(n1810), .B(n1809), .Z(n1811) );
  AND U2036 ( .A(n1812), .B(n1811), .Z(n1922) );
  NANDN U2037 ( .A(n1814), .B(n1813), .Z(n1818) );
  NAND U2038 ( .A(n1816), .B(n1815), .Z(n1817) );
  AND U2039 ( .A(n1818), .B(n1817), .Z(n2035) );
  NAND U2040 ( .A(b[0]), .B(a[27]), .Z(n1819) );
  XNOR U2041 ( .A(b[1]), .B(n1819), .Z(n1821) );
  NANDN U2042 ( .A(b[0]), .B(a[26]), .Z(n1820) );
  NAND U2043 ( .A(n1821), .B(n1820), .Z(n1983) );
  NANDN U2044 ( .A(n18113), .B(n1822), .Z(n1824) );
  XOR U2045 ( .A(b[13]), .B(a[15]), .Z(n1979) );
  NANDN U2046 ( .A(n18229), .B(n1979), .Z(n1823) );
  NAND U2047 ( .A(n1824), .B(n1823), .Z(n1982) );
  XNOR U2048 ( .A(n1983), .B(n1982), .Z(n1984) );
  XOR U2049 ( .A(b[27]), .B(b[26]), .Z(n2023) );
  XOR U2050 ( .A(b[27]), .B(a[0]), .Z(n1825) );
  NAND U2051 ( .A(n2023), .B(n1825), .Z(n1826) );
  OR U2052 ( .A(n1826), .B(n19322), .Z(n1828) );
  XOR U2053 ( .A(b[27]), .B(a[1]), .Z(n2024) );
  NAND U2054 ( .A(n19322), .B(n2024), .Z(n1827) );
  AND U2055 ( .A(n1828), .B(n1827), .Z(n2018) );
  NANDN U2056 ( .A(n19116), .B(n1829), .Z(n1831) );
  XOR U2057 ( .A(b[25]), .B(a[3]), .Z(n2015) );
  NANDN U2058 ( .A(n19179), .B(n2015), .Z(n1830) );
  NAND U2059 ( .A(n1831), .B(n1830), .Z(n2019) );
  XOR U2060 ( .A(n2018), .B(n2019), .Z(n1985) );
  XNOR U2061 ( .A(n1984), .B(n1985), .Z(n1946) );
  NANDN U2062 ( .A(n17362), .B(n1832), .Z(n1834) );
  XOR U2063 ( .A(b[7]), .B(a[21]), .Z(n1967) );
  NANDN U2064 ( .A(n17522), .B(n1967), .Z(n1833) );
  AND U2065 ( .A(n1834), .B(n1833), .Z(n2030) );
  NANDN U2066 ( .A(n17072), .B(n1835), .Z(n1837) );
  XOR U2067 ( .A(b[5]), .B(a[23]), .Z(n1958) );
  NANDN U2068 ( .A(n17223), .B(n1958), .Z(n1836) );
  AND U2069 ( .A(n1837), .B(n1836), .Z(n2028) );
  NANDN U2070 ( .A(n18673), .B(n1838), .Z(n1840) );
  XOR U2071 ( .A(b[19]), .B(a[9]), .Z(n1952) );
  NANDN U2072 ( .A(n18758), .B(n1952), .Z(n1839) );
  NAND U2073 ( .A(n1840), .B(n1839), .Z(n2027) );
  XNOR U2074 ( .A(n2028), .B(n2027), .Z(n2029) );
  XOR U2075 ( .A(n2030), .B(n2029), .Z(n1947) );
  XNOR U2076 ( .A(n1946), .B(n1947), .Z(n1948) );
  NANDN U2077 ( .A(n1842), .B(n1841), .Z(n1846) );
  OR U2078 ( .A(n1844), .B(n1843), .Z(n1845) );
  NAND U2079 ( .A(n1846), .B(n1845), .Z(n1949) );
  XNOR U2080 ( .A(n1948), .B(n1949), .Z(n1937) );
  NANDN U2081 ( .A(n1848), .B(n1847), .Z(n1852) );
  OR U2082 ( .A(n1850), .B(n1849), .Z(n1851) );
  NAND U2083 ( .A(n1852), .B(n1851), .Z(n1935) );
  NANDN U2084 ( .A(n1854), .B(n1853), .Z(n1858) );
  NANDN U2085 ( .A(n1856), .B(n1855), .Z(n1857) );
  NAND U2086 ( .A(n1858), .B(n1857), .Z(n1934) );
  XOR U2087 ( .A(n1935), .B(n1934), .Z(n1936) );
  XOR U2088 ( .A(n1937), .B(n1936), .Z(n1943) );
  NANDN U2089 ( .A(n1859), .B(n1871), .Z(n1863) );
  NANDN U2090 ( .A(n1861), .B(n1860), .Z(n1862) );
  AND U2091 ( .A(n1863), .B(n1862), .Z(n1995) );
  NANDN U2092 ( .A(n1864), .B(n2664), .Z(n1866) );
  XOR U2093 ( .A(b[3]), .B(a[25]), .Z(n1973) );
  NANDN U2094 ( .A(n17068), .B(n1973), .Z(n1865) );
  AND U2095 ( .A(n1866), .B(n1865), .Z(n2007) );
  NANDN U2096 ( .A(n1867), .B(n18439), .Z(n1869) );
  XOR U2097 ( .A(b[15]), .B(a[13]), .Z(n2020) );
  NANDN U2098 ( .A(n18311), .B(n2020), .Z(n1868) );
  NAND U2099 ( .A(n1869), .B(n1868), .Z(n2006) );
  XNOR U2100 ( .A(n2007), .B(n2006), .Z(n2008) );
  NAND U2101 ( .A(b[25]), .B(b[26]), .Z(n1870) );
  NAND U2102 ( .A(b[27]), .B(n1870), .Z(n19357) );
  NOR U2103 ( .A(n19357), .B(n1871), .Z(n2009) );
  XOR U2104 ( .A(n2008), .B(n2009), .Z(n1994) );
  XNOR U2105 ( .A(n1995), .B(n1994), .Z(n1997) );
  NANDN U2106 ( .A(n17888), .B(n1872), .Z(n1874) );
  XOR U2107 ( .A(b[11]), .B(a[17]), .Z(n1961) );
  NANDN U2108 ( .A(n18025), .B(n1961), .Z(n1873) );
  AND U2109 ( .A(n1874), .B(n1873), .Z(n2001) );
  NANDN U2110 ( .A(n18514), .B(n1875), .Z(n1877) );
  XOR U2111 ( .A(b[17]), .B(a[11]), .Z(n1964) );
  NANDN U2112 ( .A(n18585), .B(n1964), .Z(n1876) );
  NAND U2113 ( .A(n1877), .B(n1876), .Z(n2000) );
  XNOR U2114 ( .A(n2001), .B(n2000), .Z(n2002) );
  NANDN U2115 ( .A(n18853), .B(n1878), .Z(n1880) );
  XOR U2116 ( .A(b[21]), .B(a[7]), .Z(n1955) );
  NANDN U2117 ( .A(n18926), .B(n1955), .Z(n1879) );
  AND U2118 ( .A(n1880), .B(n1879), .Z(n1991) );
  NANDN U2119 ( .A(n19005), .B(n1881), .Z(n1883) );
  XOR U2120 ( .A(b[23]), .B(a[5]), .Z(n1976) );
  NANDN U2121 ( .A(n19055), .B(n1976), .Z(n1882) );
  AND U2122 ( .A(n1883), .B(n1882), .Z(n1989) );
  NANDN U2123 ( .A(n17613), .B(n1884), .Z(n1886) );
  XOR U2124 ( .A(b[9]), .B(a[19]), .Z(n1970) );
  NANDN U2125 ( .A(n17739), .B(n1970), .Z(n1885) );
  NAND U2126 ( .A(n1886), .B(n1885), .Z(n1988) );
  XNOR U2127 ( .A(n1989), .B(n1988), .Z(n1990) );
  XOR U2128 ( .A(n1991), .B(n1990), .Z(n2003) );
  XNOR U2129 ( .A(n2002), .B(n2003), .Z(n1996) );
  XOR U2130 ( .A(n1997), .B(n1996), .Z(n1941) );
  NANDN U2131 ( .A(n1888), .B(n1887), .Z(n1892) );
  NANDN U2132 ( .A(n1890), .B(n1889), .Z(n1891) );
  AND U2133 ( .A(n1892), .B(n1891), .Z(n1940) );
  XNOR U2134 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U2135 ( .A(n1943), .B(n1942), .Z(n2033) );
  NANDN U2136 ( .A(n1894), .B(n1893), .Z(n1898) );
  NAND U2137 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2138 ( .A(n1898), .B(n1897), .Z(n1931) );
  NANDN U2139 ( .A(n1900), .B(n1899), .Z(n1904) );
  NANDN U2140 ( .A(n1902), .B(n1901), .Z(n1903) );
  AND U2141 ( .A(n1904), .B(n1903), .Z(n1928) );
  NANDN U2142 ( .A(n1906), .B(n1905), .Z(n1910) );
  OR U2143 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U2144 ( .A(n1910), .B(n1909), .Z(n1929) );
  XNOR U2145 ( .A(n1928), .B(n1929), .Z(n1930) );
  XOR U2146 ( .A(n1931), .B(n1930), .Z(n2034) );
  XOR U2147 ( .A(n2033), .B(n2034), .Z(n2036) );
  XOR U2148 ( .A(n2035), .B(n2036), .Z(n1923) );
  XNOR U2149 ( .A(n1922), .B(n1923), .Z(n1924) );
  XNOR U2150 ( .A(n1925), .B(n1924), .Z(n1916) );
  XNOR U2151 ( .A(n1917), .B(n1916), .Z(n1918) );
  XNOR U2152 ( .A(n1919), .B(n1918), .Z(n1911) );
  XNOR U2153 ( .A(sreg[123]), .B(n1911), .Z(n1912) );
  XNOR U2154 ( .A(n1913), .B(n1912), .Z(c[123]) );
  NANDN U2155 ( .A(sreg[123]), .B(n1911), .Z(n1915) );
  NAND U2156 ( .A(n1913), .B(n1912), .Z(n1914) );
  NAND U2157 ( .A(n1915), .B(n1914), .Z(n2039) );
  XNOR U2158 ( .A(sreg[124]), .B(n2039), .Z(n2041) );
  NANDN U2159 ( .A(n1917), .B(n1916), .Z(n1921) );
  NANDN U2160 ( .A(n1919), .B(n1918), .Z(n1920) );
  AND U2161 ( .A(n1921), .B(n1920), .Z(n2046) );
  NANDN U2162 ( .A(n1923), .B(n1922), .Z(n1927) );
  NANDN U2163 ( .A(n1925), .B(n1924), .Z(n1926) );
  AND U2164 ( .A(n1927), .B(n1926), .Z(n2045) );
  NANDN U2165 ( .A(n1929), .B(n1928), .Z(n1933) );
  NANDN U2166 ( .A(n1931), .B(n1930), .Z(n1932) );
  AND U2167 ( .A(n1933), .B(n1932), .Z(n2053) );
  NAND U2168 ( .A(n1935), .B(n1934), .Z(n1939) );
  NAND U2169 ( .A(n1937), .B(n1936), .Z(n1938) );
  AND U2170 ( .A(n1939), .B(n1938), .Z(n2051) );
  NANDN U2171 ( .A(n1941), .B(n1940), .Z(n1945) );
  NANDN U2172 ( .A(n1943), .B(n1942), .Z(n1944) );
  AND U2173 ( .A(n1945), .B(n1944), .Z(n2050) );
  XNOR U2174 ( .A(n2051), .B(n2050), .Z(n2052) );
  XOR U2175 ( .A(n2053), .B(n2052), .Z(n2172) );
  NANDN U2176 ( .A(n1947), .B(n1946), .Z(n1951) );
  NANDN U2177 ( .A(n1949), .B(n1948), .Z(n1950) );
  AND U2178 ( .A(n1951), .B(n1950), .Z(n2142) );
  NANDN U2179 ( .A(n18673), .B(n1952), .Z(n1954) );
  XOR U2180 ( .A(b[19]), .B(a[10]), .Z(n2072) );
  NANDN U2181 ( .A(n18758), .B(n2072), .Z(n1953) );
  AND U2182 ( .A(n1954), .B(n1953), .Z(n2092) );
  NANDN U2183 ( .A(n18853), .B(n1955), .Z(n1957) );
  XOR U2184 ( .A(b[21]), .B(a[8]), .Z(n2099) );
  NANDN U2185 ( .A(n18926), .B(n2099), .Z(n1956) );
  AND U2186 ( .A(n1957), .B(n1956), .Z(n2091) );
  NANDN U2187 ( .A(n17072), .B(n1958), .Z(n1960) );
  XOR U2188 ( .A(b[5]), .B(a[24]), .Z(n2103) );
  NANDN U2189 ( .A(n17223), .B(n2103), .Z(n1959) );
  NAND U2190 ( .A(n1960), .B(n1959), .Z(n2090) );
  XOR U2191 ( .A(n2091), .B(n2090), .Z(n2093) );
  XOR U2192 ( .A(n2092), .B(n2093), .Z(n2160) );
  NANDN U2193 ( .A(n17888), .B(n1961), .Z(n1963) );
  XOR U2194 ( .A(b[11]), .B(a[18]), .Z(n2075) );
  NANDN U2195 ( .A(n18025), .B(n2075), .Z(n1962) );
  AND U2196 ( .A(n1963), .B(n1962), .Z(n2129) );
  NANDN U2197 ( .A(n18514), .B(n1964), .Z(n1966) );
  XOR U2198 ( .A(b[17]), .B(a[12]), .Z(n2109) );
  NANDN U2199 ( .A(n18585), .B(n2109), .Z(n1965) );
  AND U2200 ( .A(n1966), .B(n1965), .Z(n2128) );
  NANDN U2201 ( .A(n17362), .B(n1967), .Z(n1969) );
  XOR U2202 ( .A(b[7]), .B(a[22]), .Z(n2096) );
  NANDN U2203 ( .A(n17522), .B(n2096), .Z(n1968) );
  NAND U2204 ( .A(n1969), .B(n1968), .Z(n2127) );
  XOR U2205 ( .A(n2128), .B(n2127), .Z(n2130) );
  XOR U2206 ( .A(n2129), .B(n2130), .Z(n2158) );
  NAND U2207 ( .A(n17881), .B(n1970), .Z(n1972) );
  XNOR U2208 ( .A(b[9]), .B(a[20]), .Z(n2118) );
  NANDN U2209 ( .A(n2118), .B(n17879), .Z(n1971) );
  AND U2210 ( .A(n1972), .B(n1971), .Z(n2157) );
  XNOR U2211 ( .A(n2158), .B(n2157), .Z(n2159) );
  XNOR U2212 ( .A(n2160), .B(n2159), .Z(n2139) );
  NANDN U2213 ( .A(n17067), .B(n1973), .Z(n1975) );
  XOR U2214 ( .A(b[3]), .B(a[26]), .Z(n2106) );
  NANDN U2215 ( .A(n17068), .B(n2106), .Z(n1974) );
  AND U2216 ( .A(n1975), .B(n1974), .Z(n2086) );
  NANDN U2217 ( .A(n19005), .B(n1976), .Z(n1978) );
  XOR U2218 ( .A(b[23]), .B(a[6]), .Z(n2112) );
  NANDN U2219 ( .A(n19055), .B(n2112), .Z(n1977) );
  AND U2220 ( .A(n1978), .B(n1977), .Z(n2085) );
  NANDN U2221 ( .A(n18113), .B(n1979), .Z(n1981) );
  XOR U2222 ( .A(b[13]), .B(a[16]), .Z(n2069) );
  NANDN U2223 ( .A(n18229), .B(n2069), .Z(n1980) );
  NAND U2224 ( .A(n1981), .B(n1980), .Z(n2084) );
  XOR U2225 ( .A(n2085), .B(n2084), .Z(n2087) );
  XOR U2226 ( .A(n2086), .B(n2087), .Z(n2146) );
  NANDN U2227 ( .A(n1983), .B(n1982), .Z(n1987) );
  NANDN U2228 ( .A(n1985), .B(n1984), .Z(n1986) );
  AND U2229 ( .A(n1987), .B(n1986), .Z(n2145) );
  XNOR U2230 ( .A(n2146), .B(n2145), .Z(n2147) );
  NANDN U2231 ( .A(n1989), .B(n1988), .Z(n1993) );
  NANDN U2232 ( .A(n1991), .B(n1990), .Z(n1992) );
  NAND U2233 ( .A(n1993), .B(n1992), .Z(n2148) );
  XOR U2234 ( .A(n2147), .B(n2148), .Z(n2140) );
  XNOR U2235 ( .A(n2139), .B(n2140), .Z(n2141) );
  XOR U2236 ( .A(n2142), .B(n2141), .Z(n2165) );
  NANDN U2237 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U2238 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U2239 ( .A(n1999), .B(n1998), .Z(n2164) );
  NANDN U2240 ( .A(n2001), .B(n2000), .Z(n2005) );
  NANDN U2241 ( .A(n2003), .B(n2002), .Z(n2004) );
  AND U2242 ( .A(n2005), .B(n2004), .Z(n2136) );
  NANDN U2243 ( .A(n2007), .B(n2006), .Z(n2011) );
  NAND U2244 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U2245 ( .A(n2011), .B(n2010), .Z(n2134) );
  NAND U2246 ( .A(b[0]), .B(a[28]), .Z(n2012) );
  XNOR U2247 ( .A(b[1]), .B(n2012), .Z(n2014) );
  NANDN U2248 ( .A(b[0]), .B(a[27]), .Z(n2013) );
  NAND U2249 ( .A(n2014), .B(n2013), .Z(n2124) );
  XOR U2250 ( .A(b[27]), .B(b[28]), .Z(n19012) );
  IV U2251 ( .A(n19012), .Z(n19395) );
  ANDN U2252 ( .B(a[0]), .A(n19395), .Z(n2121) );
  NANDN U2253 ( .A(n19116), .B(n2015), .Z(n2017) );
  XOR U2254 ( .A(b[25]), .B(a[4]), .Z(n2115) );
  NANDN U2255 ( .A(n19179), .B(n2115), .Z(n2016) );
  AND U2256 ( .A(n2017), .B(n2016), .Z(n2122) );
  XOR U2257 ( .A(n2121), .B(n2122), .Z(n2123) );
  XOR U2258 ( .A(n2124), .B(n2123), .Z(n2152) );
  ANDN U2259 ( .B(n2019), .A(n2018), .Z(n2081) );
  NAND U2260 ( .A(n18439), .B(n2020), .Z(n2022) );
  XNOR U2261 ( .A(b[15]), .B(a[14]), .Z(n2066) );
  NANDN U2262 ( .A(n2066), .B(n18486), .Z(n2021) );
  AND U2263 ( .A(n2022), .B(n2021), .Z(n2078) );
  ANDN U2264 ( .B(n2023), .A(n19322), .Z(n19321) );
  NAND U2265 ( .A(n19321), .B(n2024), .Z(n2026) );
  XNOR U2266 ( .A(b[27]), .B(a[2]), .Z(n2060) );
  NANDN U2267 ( .A(n2060), .B(n19322), .Z(n2025) );
  NAND U2268 ( .A(n2026), .B(n2025), .Z(n2079) );
  XNOR U2269 ( .A(n2078), .B(n2079), .Z(n2080) );
  XNOR U2270 ( .A(n2081), .B(n2080), .Z(n2151) );
  XNOR U2271 ( .A(n2152), .B(n2151), .Z(n2154) );
  NANDN U2272 ( .A(n2028), .B(n2027), .Z(n2032) );
  NANDN U2273 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U2274 ( .A(n2032), .B(n2031), .Z(n2153) );
  XNOR U2275 ( .A(n2154), .B(n2153), .Z(n2133) );
  XNOR U2276 ( .A(n2134), .B(n2133), .Z(n2135) );
  XNOR U2277 ( .A(n2136), .B(n2135), .Z(n2163) );
  XOR U2278 ( .A(n2164), .B(n2163), .Z(n2166) );
  XOR U2279 ( .A(n2165), .B(n2166), .Z(n2170) );
  NANDN U2280 ( .A(n2034), .B(n2033), .Z(n2038) );
  NANDN U2281 ( .A(n2036), .B(n2035), .Z(n2037) );
  NAND U2282 ( .A(n2038), .B(n2037), .Z(n2169) );
  XNOR U2283 ( .A(n2170), .B(n2169), .Z(n2171) );
  XNOR U2284 ( .A(n2172), .B(n2171), .Z(n2044) );
  XOR U2285 ( .A(n2045), .B(n2044), .Z(n2047) );
  XNOR U2286 ( .A(n2046), .B(n2047), .Z(n2040) );
  XOR U2287 ( .A(n2041), .B(n2040), .Z(c[124]) );
  NANDN U2288 ( .A(n2039), .B(sreg[124]), .Z(n2043) );
  NAND U2289 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U2290 ( .A(n2043), .B(n2042), .Z(n2177) );
  NANDN U2291 ( .A(n2045), .B(n2044), .Z(n2049) );
  OR U2292 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U2293 ( .A(n2049), .B(n2048), .Z(n2180) );
  NANDN U2294 ( .A(n2051), .B(n2050), .Z(n2055) );
  NAND U2295 ( .A(n2053), .B(n2052), .Z(n2054) );
  AND U2296 ( .A(n2055), .B(n2054), .Z(n2306) );
  XOR U2297 ( .A(b[29]), .B(b[28]), .Z(n2255) );
  XOR U2298 ( .A(b[29]), .B(a[0]), .Z(n2056) );
  NAND U2299 ( .A(n2255), .B(n2056), .Z(n2057) );
  OR U2300 ( .A(n2057), .B(n19012), .Z(n2059) );
  XOR U2301 ( .A(b[29]), .B(a[1]), .Z(n2256) );
  NAND U2302 ( .A(n19012), .B(n2256), .Z(n2058) );
  AND U2303 ( .A(n2059), .B(n2058), .Z(n2254) );
  NANDN U2304 ( .A(n2060), .B(n19321), .Z(n2062) );
  XOR U2305 ( .A(b[27]), .B(a[3]), .Z(n2220) );
  NANDN U2306 ( .A(n19277), .B(n2220), .Z(n2061) );
  AND U2307 ( .A(n2062), .B(n2061), .Z(n2253) );
  XOR U2308 ( .A(n2254), .B(n2253), .Z(n2288) );
  NAND U2309 ( .A(b[0]), .B(a[29]), .Z(n2063) );
  XNOR U2310 ( .A(b[1]), .B(n2063), .Z(n2065) );
  NANDN U2311 ( .A(b[0]), .B(a[28]), .Z(n2064) );
  NAND U2312 ( .A(n2065), .B(n2064), .Z(n2286) );
  NANDN U2313 ( .A(n2066), .B(n18439), .Z(n2068) );
  XNOR U2314 ( .A(b[15]), .B(a[15]), .Z(n2268) );
  NANDN U2315 ( .A(n2268), .B(n18486), .Z(n2067) );
  NAND U2316 ( .A(n2068), .B(n2067), .Z(n2287) );
  XOR U2317 ( .A(n2286), .B(n2287), .Z(n2289) );
  XOR U2318 ( .A(n2288), .B(n2289), .Z(n2248) );
  NANDN U2319 ( .A(n18113), .B(n2069), .Z(n2071) );
  XOR U2320 ( .A(b[13]), .B(a[17]), .Z(n2277) );
  NANDN U2321 ( .A(n18229), .B(n2277), .Z(n2070) );
  AND U2322 ( .A(n2071), .B(n2070), .Z(n2295) );
  NANDN U2323 ( .A(n18673), .B(n2072), .Z(n2074) );
  XOR U2324 ( .A(b[19]), .B(a[11]), .Z(n2280) );
  NANDN U2325 ( .A(n18758), .B(n2280), .Z(n2073) );
  AND U2326 ( .A(n2074), .B(n2073), .Z(n2293) );
  NANDN U2327 ( .A(n17888), .B(n2075), .Z(n2077) );
  XOR U2328 ( .A(b[11]), .B(a[19]), .Z(n2271) );
  NANDN U2329 ( .A(n18025), .B(n2271), .Z(n2076) );
  NAND U2330 ( .A(n2077), .B(n2076), .Z(n2292) );
  XNOR U2331 ( .A(n2293), .B(n2292), .Z(n2294) );
  XNOR U2332 ( .A(n2295), .B(n2294), .Z(n2247) );
  XNOR U2333 ( .A(n2248), .B(n2247), .Z(n2249) );
  NANDN U2334 ( .A(n2079), .B(n2078), .Z(n2083) );
  NANDN U2335 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U2336 ( .A(n2083), .B(n2082), .Z(n2250) );
  XNOR U2337 ( .A(n2249), .B(n2250), .Z(n2193) );
  NANDN U2338 ( .A(n2085), .B(n2084), .Z(n2089) );
  OR U2339 ( .A(n2087), .B(n2086), .Z(n2088) );
  AND U2340 ( .A(n2089), .B(n2088), .Z(n2191) );
  NANDN U2341 ( .A(n2091), .B(n2090), .Z(n2095) );
  OR U2342 ( .A(n2093), .B(n2092), .Z(n2094) );
  AND U2343 ( .A(n2095), .B(n2094), .Z(n2199) );
  NANDN U2344 ( .A(n17362), .B(n2096), .Z(n2098) );
  XOR U2345 ( .A(b[7]), .B(a[23]), .Z(n2283) );
  NANDN U2346 ( .A(n17522), .B(n2283), .Z(n2097) );
  AND U2347 ( .A(n2098), .B(n2097), .Z(n2209) );
  NANDN U2348 ( .A(n18853), .B(n2099), .Z(n2101) );
  XOR U2349 ( .A(b[21]), .B(a[9]), .Z(n2232) );
  NANDN U2350 ( .A(n18926), .B(n2232), .Z(n2100) );
  NAND U2351 ( .A(n2101), .B(n2100), .Z(n2208) );
  XNOR U2352 ( .A(n2209), .B(n2208), .Z(n2210) );
  NAND U2353 ( .A(b[27]), .B(b[28]), .Z(n2102) );
  NAND U2354 ( .A(b[29]), .B(n2102), .Z(n19420) );
  NOR U2355 ( .A(n19420), .B(n2121), .Z(n2211) );
  XOR U2356 ( .A(n2210), .B(n2211), .Z(n2196) );
  NANDN U2357 ( .A(n17072), .B(n2103), .Z(n2105) );
  XOR U2358 ( .A(b[5]), .B(a[25]), .Z(n2262) );
  NANDN U2359 ( .A(n17223), .B(n2262), .Z(n2104) );
  AND U2360 ( .A(n2105), .B(n2104), .Z(n2217) );
  NANDN U2361 ( .A(n17067), .B(n2106), .Z(n2108) );
  XOR U2362 ( .A(b[3]), .B(a[27]), .Z(n2265) );
  NANDN U2363 ( .A(n17068), .B(n2265), .Z(n2107) );
  AND U2364 ( .A(n2108), .B(n2107), .Z(n2215) );
  NANDN U2365 ( .A(n18514), .B(n2109), .Z(n2111) );
  XOR U2366 ( .A(b[17]), .B(a[13]), .Z(n2259) );
  NANDN U2367 ( .A(n18585), .B(n2259), .Z(n2110) );
  NAND U2368 ( .A(n2111), .B(n2110), .Z(n2214) );
  XNOR U2369 ( .A(n2215), .B(n2214), .Z(n2216) );
  XOR U2370 ( .A(n2217), .B(n2216), .Z(n2197) );
  XNOR U2371 ( .A(n2196), .B(n2197), .Z(n2198) );
  XNOR U2372 ( .A(n2199), .B(n2198), .Z(n2190) );
  XNOR U2373 ( .A(n2191), .B(n2190), .Z(n2192) );
  XOR U2374 ( .A(n2193), .B(n2192), .Z(n2299) );
  NANDN U2375 ( .A(n19005), .B(n2112), .Z(n2114) );
  XOR U2376 ( .A(b[23]), .B(a[7]), .Z(n2226) );
  NANDN U2377 ( .A(n19055), .B(n2226), .Z(n2113) );
  AND U2378 ( .A(n2114), .B(n2113), .Z(n2204) );
  NANDN U2379 ( .A(n19116), .B(n2115), .Z(n2117) );
  XOR U2380 ( .A(b[25]), .B(a[5]), .Z(n2229) );
  NANDN U2381 ( .A(n19179), .B(n2229), .Z(n2116) );
  AND U2382 ( .A(n2117), .B(n2116), .Z(n2203) );
  NANDN U2383 ( .A(n2118), .B(n17881), .Z(n2120) );
  XOR U2384 ( .A(b[9]), .B(a[21]), .Z(n2274) );
  NANDN U2385 ( .A(n17739), .B(n2274), .Z(n2119) );
  NAND U2386 ( .A(n2120), .B(n2119), .Z(n2202) );
  XOR U2387 ( .A(n2203), .B(n2202), .Z(n2205) );
  XOR U2388 ( .A(n2204), .B(n2205), .Z(n2242) );
  NANDN U2389 ( .A(n2122), .B(n2121), .Z(n2126) );
  OR U2390 ( .A(n2124), .B(n2123), .Z(n2125) );
  AND U2391 ( .A(n2126), .B(n2125), .Z(n2241) );
  XNOR U2392 ( .A(n2242), .B(n2241), .Z(n2243) );
  NANDN U2393 ( .A(n2128), .B(n2127), .Z(n2132) );
  OR U2394 ( .A(n2130), .B(n2129), .Z(n2131) );
  NAND U2395 ( .A(n2132), .B(n2131), .Z(n2244) );
  XNOR U2396 ( .A(n2243), .B(n2244), .Z(n2298) );
  XNOR U2397 ( .A(n2299), .B(n2298), .Z(n2300) );
  NANDN U2398 ( .A(n2134), .B(n2133), .Z(n2138) );
  NANDN U2399 ( .A(n2136), .B(n2135), .Z(n2137) );
  NAND U2400 ( .A(n2138), .B(n2137), .Z(n2301) );
  XNOR U2401 ( .A(n2300), .B(n2301), .Z(n2187) );
  NANDN U2402 ( .A(n2140), .B(n2139), .Z(n2144) );
  NAND U2403 ( .A(n2142), .B(n2141), .Z(n2143) );
  AND U2404 ( .A(n2144), .B(n2143), .Z(n2185) );
  NANDN U2405 ( .A(n2146), .B(n2145), .Z(n2150) );
  NANDN U2406 ( .A(n2148), .B(n2147), .Z(n2149) );
  AND U2407 ( .A(n2150), .B(n2149), .Z(n2238) );
  NANDN U2408 ( .A(n2152), .B(n2151), .Z(n2156) );
  NAND U2409 ( .A(n2154), .B(n2153), .Z(n2155) );
  AND U2410 ( .A(n2156), .B(n2155), .Z(n2236) );
  NANDN U2411 ( .A(n2158), .B(n2157), .Z(n2162) );
  NANDN U2412 ( .A(n2160), .B(n2159), .Z(n2161) );
  NAND U2413 ( .A(n2162), .B(n2161), .Z(n2235) );
  XNOR U2414 ( .A(n2236), .B(n2235), .Z(n2237) );
  XNOR U2415 ( .A(n2238), .B(n2237), .Z(n2184) );
  XNOR U2416 ( .A(n2185), .B(n2184), .Z(n2186) );
  XOR U2417 ( .A(n2187), .B(n2186), .Z(n2305) );
  NANDN U2418 ( .A(n2164), .B(n2163), .Z(n2168) );
  OR U2419 ( .A(n2166), .B(n2165), .Z(n2167) );
  NAND U2420 ( .A(n2168), .B(n2167), .Z(n2304) );
  XOR U2421 ( .A(n2305), .B(n2304), .Z(n2307) );
  XOR U2422 ( .A(n2306), .B(n2307), .Z(n2179) );
  NANDN U2423 ( .A(n2170), .B(n2169), .Z(n2174) );
  NANDN U2424 ( .A(n2172), .B(n2171), .Z(n2173) );
  NAND U2425 ( .A(n2174), .B(n2173), .Z(n2178) );
  XOR U2426 ( .A(n2179), .B(n2178), .Z(n2181) );
  XOR U2427 ( .A(n2180), .B(n2181), .Z(n2176) );
  XOR U2428 ( .A(sreg[125]), .B(n2176), .Z(n2175) );
  XNOR U2429 ( .A(n2177), .B(n2175), .Z(c[125]) );
  XOR U2430 ( .A(sreg[126]), .B(n2310), .Z(n2312) );
  NANDN U2431 ( .A(n2179), .B(n2178), .Z(n2183) );
  OR U2432 ( .A(n2181), .B(n2180), .Z(n2182) );
  AND U2433 ( .A(n2183), .B(n2182), .Z(n2318) );
  NANDN U2434 ( .A(n2185), .B(n2184), .Z(n2189) );
  NAND U2435 ( .A(n2187), .B(n2186), .Z(n2188) );
  AND U2436 ( .A(n2189), .B(n2188), .Z(n2452) );
  NANDN U2437 ( .A(n2191), .B(n2190), .Z(n2195) );
  NAND U2438 ( .A(n2193), .B(n2192), .Z(n2194) );
  AND U2439 ( .A(n2195), .B(n2194), .Z(n2329) );
  NANDN U2440 ( .A(n2197), .B(n2196), .Z(n2201) );
  NANDN U2441 ( .A(n2199), .B(n2198), .Z(n2200) );
  AND U2442 ( .A(n2201), .B(n2200), .Z(n2328) );
  NANDN U2443 ( .A(n2203), .B(n2202), .Z(n2207) );
  OR U2444 ( .A(n2205), .B(n2204), .Z(n2206) );
  AND U2445 ( .A(n2207), .B(n2206), .Z(n2334) );
  NANDN U2446 ( .A(n2209), .B(n2208), .Z(n2213) );
  NAND U2447 ( .A(n2211), .B(n2210), .Z(n2212) );
  NAND U2448 ( .A(n2213), .B(n2212), .Z(n2333) );
  XNOR U2449 ( .A(n2334), .B(n2333), .Z(n2335) );
  NANDN U2450 ( .A(n2215), .B(n2214), .Z(n2219) );
  NANDN U2451 ( .A(n2217), .B(n2216), .Z(n2218) );
  AND U2452 ( .A(n2219), .B(n2218), .Z(n2378) );
  XOR U2453 ( .A(b[29]), .B(b[30]), .Z(n19411) );
  IV U2454 ( .A(n19411), .Z(n19426) );
  ANDN U2455 ( .B(a[0]), .A(n19426), .Z(n2423) );
  IV U2456 ( .A(n19321), .Z(n19237) );
  NANDN U2457 ( .A(n19237), .B(n2220), .Z(n2222) );
  XOR U2458 ( .A(b[27]), .B(a[4]), .Z(n2393) );
  NANDN U2459 ( .A(n19277), .B(n2393), .Z(n2221) );
  AND U2460 ( .A(n2222), .B(n2221), .Z(n2364) );
  XNOR U2461 ( .A(n2423), .B(n2364), .Z(n2365) );
  NAND U2462 ( .A(b[0]), .B(a[30]), .Z(n2223) );
  XNOR U2463 ( .A(b[1]), .B(n2223), .Z(n2225) );
  NANDN U2464 ( .A(b[0]), .B(a[29]), .Z(n2224) );
  NAND U2465 ( .A(n2225), .B(n2224), .Z(n2366) );
  XNOR U2466 ( .A(n2365), .B(n2366), .Z(n2375) );
  NANDN U2467 ( .A(n19005), .B(n2226), .Z(n2228) );
  XOR U2468 ( .A(b[23]), .B(a[8]), .Z(n2387) );
  NANDN U2469 ( .A(n19055), .B(n2387), .Z(n2227) );
  AND U2470 ( .A(n2228), .B(n2227), .Z(n2440) );
  NANDN U2471 ( .A(n19116), .B(n2229), .Z(n2231) );
  XOR U2472 ( .A(b[25]), .B(a[6]), .Z(n2390) );
  NANDN U2473 ( .A(n19179), .B(n2390), .Z(n2230) );
  AND U2474 ( .A(n2231), .B(n2230), .Z(n2438) );
  NANDN U2475 ( .A(n18853), .B(n2232), .Z(n2234) );
  XOR U2476 ( .A(b[21]), .B(a[10]), .Z(n2399) );
  NANDN U2477 ( .A(n18926), .B(n2399), .Z(n2233) );
  NAND U2478 ( .A(n2234), .B(n2233), .Z(n2437) );
  XNOR U2479 ( .A(n2438), .B(n2437), .Z(n2439) );
  XOR U2480 ( .A(n2440), .B(n2439), .Z(n2376) );
  XNOR U2481 ( .A(n2375), .B(n2376), .Z(n2377) );
  XOR U2482 ( .A(n2378), .B(n2377), .Z(n2336) );
  XNOR U2483 ( .A(n2335), .B(n2336), .Z(n2327) );
  XOR U2484 ( .A(n2328), .B(n2327), .Z(n2330) );
  XOR U2485 ( .A(n2329), .B(n2330), .Z(n2323) );
  NANDN U2486 ( .A(n2236), .B(n2235), .Z(n2240) );
  NANDN U2487 ( .A(n2238), .B(n2237), .Z(n2239) );
  AND U2488 ( .A(n2240), .B(n2239), .Z(n2322) );
  NANDN U2489 ( .A(n2242), .B(n2241), .Z(n2246) );
  NANDN U2490 ( .A(n2244), .B(n2243), .Z(n2245) );
  AND U2491 ( .A(n2246), .B(n2245), .Z(n2372) );
  NANDN U2492 ( .A(n2248), .B(n2247), .Z(n2252) );
  NANDN U2493 ( .A(n2250), .B(n2249), .Z(n2251) );
  AND U2494 ( .A(n2252), .B(n2251), .Z(n2369) );
  NOR U2495 ( .A(n2254), .B(n2253), .Z(n2427) );
  ANDN U2496 ( .B(n2255), .A(n19012), .Z(n19065) );
  NAND U2497 ( .A(n19065), .B(n2256), .Z(n2258) );
  XNOR U2498 ( .A(b[29]), .B(a[2]), .Z(n2351) );
  NANDN U2499 ( .A(n2351), .B(n19012), .Z(n2257) );
  AND U2500 ( .A(n2258), .B(n2257), .Z(n2425) );
  NAND U2501 ( .A(n18683), .B(n2259), .Z(n2261) );
  XNOR U2502 ( .A(b[17]), .B(a[14]), .Z(n2420) );
  NANDN U2503 ( .A(n2420), .B(n18684), .Z(n2260) );
  NAND U2504 ( .A(n2261), .B(n2260), .Z(n2426) );
  XOR U2505 ( .A(n2425), .B(n2426), .Z(n2428) );
  XOR U2506 ( .A(n2427), .B(n2428), .Z(n2382) );
  NANDN U2507 ( .A(n17072), .B(n2262), .Z(n2264) );
  XOR U2508 ( .A(b[5]), .B(a[26]), .Z(n2411) );
  NANDN U2509 ( .A(n17223), .B(n2411), .Z(n2263) );
  AND U2510 ( .A(n2264), .B(n2263), .Z(n2446) );
  NANDN U2511 ( .A(n17067), .B(n2265), .Z(n2267) );
  XOR U2512 ( .A(b[3]), .B(a[28]), .Z(n2417) );
  NANDN U2513 ( .A(n17068), .B(n2417), .Z(n2266) );
  AND U2514 ( .A(n2267), .B(n2266), .Z(n2444) );
  NANDN U2515 ( .A(n2268), .B(n18439), .Z(n2270) );
  XOR U2516 ( .A(b[15]), .B(a[16]), .Z(n2361) );
  NANDN U2517 ( .A(n18311), .B(n2361), .Z(n2269) );
  NAND U2518 ( .A(n2270), .B(n2269), .Z(n2443) );
  XNOR U2519 ( .A(n2444), .B(n2443), .Z(n2445) );
  XNOR U2520 ( .A(n2446), .B(n2445), .Z(n2381) );
  XNOR U2521 ( .A(n2382), .B(n2381), .Z(n2384) );
  NANDN U2522 ( .A(n17888), .B(n2271), .Z(n2273) );
  XOR U2523 ( .A(b[11]), .B(a[20]), .Z(n2405) );
  NANDN U2524 ( .A(n18025), .B(n2405), .Z(n2272) );
  AND U2525 ( .A(n2273), .B(n2272), .Z(n2432) );
  NANDN U2526 ( .A(n17613), .B(n2274), .Z(n2276) );
  XOR U2527 ( .A(b[9]), .B(a[22]), .Z(n2402) );
  NANDN U2528 ( .A(n17739), .B(n2402), .Z(n2275) );
  NAND U2529 ( .A(n2276), .B(n2275), .Z(n2431) );
  XNOR U2530 ( .A(n2432), .B(n2431), .Z(n2433) );
  NANDN U2531 ( .A(n18113), .B(n2277), .Z(n2279) );
  XOR U2532 ( .A(b[13]), .B(a[18]), .Z(n2396) );
  NANDN U2533 ( .A(n18229), .B(n2396), .Z(n2278) );
  AND U2534 ( .A(n2279), .B(n2278), .Z(n2348) );
  NANDN U2535 ( .A(n18673), .B(n2280), .Z(n2282) );
  XOR U2536 ( .A(b[19]), .B(a[12]), .Z(n2414) );
  NANDN U2537 ( .A(n18758), .B(n2414), .Z(n2281) );
  AND U2538 ( .A(n2282), .B(n2281), .Z(n2346) );
  NANDN U2539 ( .A(n17362), .B(n2283), .Z(n2285) );
  XOR U2540 ( .A(b[7]), .B(a[24]), .Z(n2408) );
  NANDN U2541 ( .A(n17522), .B(n2408), .Z(n2284) );
  NAND U2542 ( .A(n2285), .B(n2284), .Z(n2345) );
  XNOR U2543 ( .A(n2346), .B(n2345), .Z(n2347) );
  XOR U2544 ( .A(n2348), .B(n2347), .Z(n2434) );
  XNOR U2545 ( .A(n2433), .B(n2434), .Z(n2383) );
  XOR U2546 ( .A(n2384), .B(n2383), .Z(n2342) );
  NANDN U2547 ( .A(n2287), .B(n2286), .Z(n2291) );
  OR U2548 ( .A(n2289), .B(n2288), .Z(n2290) );
  AND U2549 ( .A(n2291), .B(n2290), .Z(n2340) );
  NANDN U2550 ( .A(n2293), .B(n2292), .Z(n2297) );
  NANDN U2551 ( .A(n2295), .B(n2294), .Z(n2296) );
  AND U2552 ( .A(n2297), .B(n2296), .Z(n2339) );
  XNOR U2553 ( .A(n2340), .B(n2339), .Z(n2341) );
  XOR U2554 ( .A(n2342), .B(n2341), .Z(n2370) );
  XNOR U2555 ( .A(n2369), .B(n2370), .Z(n2371) );
  XNOR U2556 ( .A(n2372), .B(n2371), .Z(n2321) );
  XOR U2557 ( .A(n2322), .B(n2321), .Z(n2324) );
  XOR U2558 ( .A(n2323), .B(n2324), .Z(n2450) );
  NANDN U2559 ( .A(n2299), .B(n2298), .Z(n2303) );
  NANDN U2560 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U2561 ( .A(n2303), .B(n2302), .Z(n2449) );
  XNOR U2562 ( .A(n2450), .B(n2449), .Z(n2451) );
  XOR U2563 ( .A(n2452), .B(n2451), .Z(n2316) );
  NANDN U2564 ( .A(n2305), .B(n2304), .Z(n2309) );
  OR U2565 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U2566 ( .A(n2309), .B(n2308), .Z(n2315) );
  XNOR U2567 ( .A(n2316), .B(n2315), .Z(n2317) );
  XNOR U2568 ( .A(n2318), .B(n2317), .Z(n2311) );
  XNOR U2569 ( .A(n2312), .B(n2311), .Z(c[126]) );
  OR U2570 ( .A(sreg[126]), .B(n2310), .Z(n2314) );
  NAND U2571 ( .A(n2312), .B(n2311), .Z(n2313) );
  AND U2572 ( .A(n2314), .B(n2313), .Z(n2598) );
  NANDN U2573 ( .A(n2316), .B(n2315), .Z(n2320) );
  NANDN U2574 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U2575 ( .A(n2320), .B(n2319), .Z(n2457) );
  NANDN U2576 ( .A(n2322), .B(n2321), .Z(n2326) );
  OR U2577 ( .A(n2324), .B(n2323), .Z(n2325) );
  AND U2578 ( .A(n2326), .B(n2325), .Z(n2593) );
  NANDN U2579 ( .A(n2328), .B(n2327), .Z(n2332) );
  OR U2580 ( .A(n2330), .B(n2329), .Z(n2331) );
  AND U2581 ( .A(n2332), .B(n2331), .Z(n2590) );
  NANDN U2582 ( .A(n2334), .B(n2333), .Z(n2338) );
  NANDN U2583 ( .A(n2336), .B(n2335), .Z(n2337) );
  AND U2584 ( .A(n2338), .B(n2337), .Z(n2469) );
  NANDN U2585 ( .A(n2340), .B(n2339), .Z(n2344) );
  NANDN U2586 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U2587 ( .A(n2344), .B(n2343), .Z(n2467) );
  NANDN U2588 ( .A(n2346), .B(n2345), .Z(n2350) );
  NANDN U2589 ( .A(n2348), .B(n2347), .Z(n2349) );
  AND U2590 ( .A(n2350), .B(n2349), .Z(n2575) );
  NANDN U2591 ( .A(n2351), .B(n19065), .Z(n2353) );
  XOR U2592 ( .A(b[29]), .B(a[3]), .Z(n2557) );
  NANDN U2593 ( .A(n19395), .B(n2557), .Z(n2352) );
  AND U2594 ( .A(n2353), .B(n2352), .Z(n2510) );
  XOR U2595 ( .A(b[30]), .B(b[31]), .Z(n2354) );
  ANDN U2596 ( .B(n2354), .A(n19411), .Z(n19409) );
  IV U2597 ( .A(n19409), .Z(n19425) );
  XOR U2598 ( .A(a[0]), .B(b[31]), .Z(n2355) );
  NANDN U2599 ( .A(n19425), .B(n2355), .Z(n2357) );
  XOR U2600 ( .A(b[31]), .B(a[1]), .Z(n2521) );
  ANDN U2601 ( .B(n2521), .A(n19426), .Z(n2356) );
  ANDN U2602 ( .B(n2357), .A(n2356), .Z(n2509) );
  XOR U2603 ( .A(n2510), .B(n2509), .Z(n2541) );
  NAND U2604 ( .A(b[0]), .B(a[31]), .Z(n2358) );
  XNOR U2605 ( .A(b[1]), .B(n2358), .Z(n2360) );
  NANDN U2606 ( .A(b[0]), .B(a[30]), .Z(n2359) );
  NAND U2607 ( .A(n2360), .B(n2359), .Z(n2539) );
  NAND U2608 ( .A(n18439), .B(n2361), .Z(n2363) );
  XNOR U2609 ( .A(b[15]), .B(a[17]), .Z(n2548) );
  NANDN U2610 ( .A(n2548), .B(n18486), .Z(n2362) );
  NAND U2611 ( .A(n2363), .B(n2362), .Z(n2540) );
  XOR U2612 ( .A(n2539), .B(n2540), .Z(n2542) );
  XOR U2613 ( .A(n2541), .B(n2542), .Z(n2573) );
  NANDN U2614 ( .A(n2364), .B(n2423), .Z(n2368) );
  NANDN U2615 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U2616 ( .A(n2368), .B(n2367), .Z(n2572) );
  XNOR U2617 ( .A(n2573), .B(n2572), .Z(n2574) );
  XOR U2618 ( .A(n2575), .B(n2574), .Z(n2468) );
  XOR U2619 ( .A(n2467), .B(n2468), .Z(n2470) );
  XOR U2620 ( .A(n2469), .B(n2470), .Z(n2464) );
  NANDN U2621 ( .A(n2370), .B(n2369), .Z(n2374) );
  NANDN U2622 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U2623 ( .A(n2374), .B(n2373), .Z(n2462) );
  NANDN U2624 ( .A(n2376), .B(n2375), .Z(n2380) );
  NANDN U2625 ( .A(n2378), .B(n2377), .Z(n2379) );
  AND U2626 ( .A(n2380), .B(n2379), .Z(n2585) );
  NANDN U2627 ( .A(n2382), .B(n2381), .Z(n2386) );
  NAND U2628 ( .A(n2384), .B(n2383), .Z(n2385) );
  NAND U2629 ( .A(n2386), .B(n2385), .Z(n2584) );
  XNOR U2630 ( .A(n2585), .B(n2584), .Z(n2587) );
  NANDN U2631 ( .A(n19005), .B(n2387), .Z(n2389) );
  XOR U2632 ( .A(b[23]), .B(a[9]), .Z(n2524) );
  NANDN U2633 ( .A(n19055), .B(n2524), .Z(n2388) );
  AND U2634 ( .A(n2389), .B(n2388), .Z(n2499) );
  NANDN U2635 ( .A(n19116), .B(n2390), .Z(n2392) );
  XOR U2636 ( .A(b[25]), .B(a[7]), .Z(n2479) );
  NANDN U2637 ( .A(n19179), .B(n2479), .Z(n2391) );
  AND U2638 ( .A(n2392), .B(n2391), .Z(n2498) );
  NANDN U2639 ( .A(n19237), .B(n2393), .Z(n2395) );
  XOR U2640 ( .A(b[27]), .B(a[5]), .Z(n2482) );
  NANDN U2641 ( .A(n19277), .B(n2482), .Z(n2394) );
  NAND U2642 ( .A(n2395), .B(n2394), .Z(n2497) );
  XOR U2643 ( .A(n2498), .B(n2497), .Z(n2500) );
  XOR U2644 ( .A(n2499), .B(n2500), .Z(n2475) );
  NANDN U2645 ( .A(n18113), .B(n2396), .Z(n2398) );
  XOR U2646 ( .A(b[13]), .B(a[19]), .Z(n2551) );
  NANDN U2647 ( .A(n18229), .B(n2551), .Z(n2397) );
  AND U2648 ( .A(n2398), .B(n2397), .Z(n2562) );
  NANDN U2649 ( .A(n18853), .B(n2399), .Z(n2401) );
  XOR U2650 ( .A(b[21]), .B(a[11]), .Z(n2545) );
  NANDN U2651 ( .A(n18926), .B(n2545), .Z(n2400) );
  AND U2652 ( .A(n2401), .B(n2400), .Z(n2561) );
  NANDN U2653 ( .A(n17613), .B(n2402), .Z(n2404) );
  XOR U2654 ( .A(b[9]), .B(a[23]), .Z(n2518) );
  NANDN U2655 ( .A(n17739), .B(n2518), .Z(n2403) );
  NAND U2656 ( .A(n2404), .B(n2403), .Z(n2560) );
  XOR U2657 ( .A(n2561), .B(n2560), .Z(n2563) );
  XOR U2658 ( .A(n2562), .B(n2563), .Z(n2474) );
  NAND U2659 ( .A(n18084), .B(n2405), .Z(n2407) );
  XNOR U2660 ( .A(b[11]), .B(a[21]), .Z(n2485) );
  NANDN U2661 ( .A(n2485), .B(n18085), .Z(n2406) );
  AND U2662 ( .A(n2407), .B(n2406), .Z(n2473) );
  XOR U2663 ( .A(n2474), .B(n2473), .Z(n2476) );
  XOR U2664 ( .A(n2475), .B(n2476), .Z(n2579) );
  NANDN U2665 ( .A(n17362), .B(n2408), .Z(n2410) );
  XOR U2666 ( .A(b[7]), .B(a[25]), .Z(n2488) );
  NANDN U2667 ( .A(n17522), .B(n2488), .Z(n2409) );
  AND U2668 ( .A(n2410), .B(n2409), .Z(n2506) );
  NANDN U2669 ( .A(n17072), .B(n2411), .Z(n2413) );
  XOR U2670 ( .A(b[5]), .B(a[27]), .Z(n2491) );
  NANDN U2671 ( .A(n17223), .B(n2491), .Z(n2412) );
  AND U2672 ( .A(n2413), .B(n2412), .Z(n2504) );
  NANDN U2673 ( .A(n18673), .B(n2414), .Z(n2416) );
  XOR U2674 ( .A(b[19]), .B(a[13]), .Z(n2494) );
  NANDN U2675 ( .A(n18758), .B(n2494), .Z(n2415) );
  NAND U2676 ( .A(n2416), .B(n2415), .Z(n2503) );
  XNOR U2677 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U2678 ( .A(n2506), .B(n2505), .Z(n2566) );
  NANDN U2679 ( .A(n17067), .B(n2417), .Z(n2419) );
  XOR U2680 ( .A(b[3]), .B(a[29]), .Z(n2511) );
  NANDN U2681 ( .A(n17068), .B(n2511), .Z(n2418) );
  AND U2682 ( .A(n2419), .B(n2418), .Z(n2536) );
  NANDN U2683 ( .A(n2420), .B(n18683), .Z(n2422) );
  XOR U2684 ( .A(b[17]), .B(a[15]), .Z(n2515) );
  NANDN U2685 ( .A(n18585), .B(n2515), .Z(n2421) );
  AND U2686 ( .A(n2422), .B(n2421), .Z(n2534) );
  NAND U2687 ( .A(b[29]), .B(b[30]), .Z(n19443) );
  ANDN U2688 ( .B(n19443), .A(n2423), .Z(n2424) );
  AND U2689 ( .A(b[31]), .B(n2424), .Z(n2533) );
  XNOR U2690 ( .A(n2534), .B(n2533), .Z(n2535) );
  XOR U2691 ( .A(n2536), .B(n2535), .Z(n2567) );
  XNOR U2692 ( .A(n2566), .B(n2567), .Z(n2568) );
  NANDN U2693 ( .A(n2426), .B(n2425), .Z(n2430) );
  OR U2694 ( .A(n2428), .B(n2427), .Z(n2429) );
  NAND U2695 ( .A(n2430), .B(n2429), .Z(n2569) );
  XNOR U2696 ( .A(n2568), .B(n2569), .Z(n2578) );
  XNOR U2697 ( .A(n2579), .B(n2578), .Z(n2580) );
  NANDN U2698 ( .A(n2432), .B(n2431), .Z(n2436) );
  NANDN U2699 ( .A(n2434), .B(n2433), .Z(n2435) );
  AND U2700 ( .A(n2436), .B(n2435), .Z(n2530) );
  NANDN U2701 ( .A(n2438), .B(n2437), .Z(n2442) );
  NANDN U2702 ( .A(n2440), .B(n2439), .Z(n2441) );
  AND U2703 ( .A(n2442), .B(n2441), .Z(n2528) );
  NANDN U2704 ( .A(n2444), .B(n2443), .Z(n2448) );
  NANDN U2705 ( .A(n2446), .B(n2445), .Z(n2447) );
  NAND U2706 ( .A(n2448), .B(n2447), .Z(n2527) );
  XNOR U2707 ( .A(n2528), .B(n2527), .Z(n2529) );
  XOR U2708 ( .A(n2530), .B(n2529), .Z(n2581) );
  XNOR U2709 ( .A(n2580), .B(n2581), .Z(n2586) );
  XNOR U2710 ( .A(n2587), .B(n2586), .Z(n2461) );
  XNOR U2711 ( .A(n2462), .B(n2461), .Z(n2463) );
  XOR U2712 ( .A(n2464), .B(n2463), .Z(n2591) );
  XNOR U2713 ( .A(n2590), .B(n2591), .Z(n2592) );
  XNOR U2714 ( .A(n2593), .B(n2592), .Z(n2455) );
  NANDN U2715 ( .A(n2450), .B(n2449), .Z(n2454) );
  NAND U2716 ( .A(n2452), .B(n2451), .Z(n2453) );
  NAND U2717 ( .A(n2454), .B(n2453), .Z(n2456) );
  XOR U2718 ( .A(n2455), .B(n2456), .Z(n2458) );
  XOR U2719 ( .A(n2457), .B(n2458), .Z(n2596) );
  XNOR U2720 ( .A(n2596), .B(sreg[127]), .Z(n2597) );
  XOR U2721 ( .A(n2598), .B(n2597), .Z(c[127]) );
  NANDN U2722 ( .A(n2456), .B(n2455), .Z(n2460) );
  OR U2723 ( .A(n2458), .B(n2457), .Z(n2459) );
  AND U2724 ( .A(n2460), .B(n2459), .Z(n2607) );
  NANDN U2725 ( .A(n2462), .B(n2461), .Z(n2466) );
  NANDN U2726 ( .A(n2464), .B(n2463), .Z(n2465) );
  AND U2727 ( .A(n2466), .B(n2465), .Z(n2746) );
  NANDN U2728 ( .A(n2468), .B(n2467), .Z(n2472) );
  OR U2729 ( .A(n2470), .B(n2469), .Z(n2471) );
  AND U2730 ( .A(n2472), .B(n2471), .Z(n2744) );
  NANDN U2731 ( .A(n2474), .B(n2473), .Z(n2478) );
  OR U2732 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U2733 ( .A(n2478), .B(n2477), .Z(n2643) );
  NANDN U2734 ( .A(n19116), .B(n2479), .Z(n2481) );
  XOR U2735 ( .A(b[25]), .B(a[8]), .Z(n2668) );
  NANDN U2736 ( .A(n19179), .B(n2668), .Z(n2480) );
  AND U2737 ( .A(n2481), .B(n2480), .Z(n2688) );
  NANDN U2738 ( .A(n19237), .B(n2482), .Z(n2484) );
  XOR U2739 ( .A(b[27]), .B(a[6]), .Z(n2677) );
  NANDN U2740 ( .A(n19277), .B(n2677), .Z(n2483) );
  AND U2741 ( .A(n2484), .B(n2483), .Z(n2687) );
  NANDN U2742 ( .A(n2485), .B(n18084), .Z(n2487) );
  XOR U2743 ( .A(b[11]), .B(a[22]), .Z(n2661) );
  NANDN U2744 ( .A(n18025), .B(n2661), .Z(n2486) );
  NAND U2745 ( .A(n2487), .B(n2486), .Z(n2686) );
  XOR U2746 ( .A(n2687), .B(n2686), .Z(n2689) );
  XOR U2747 ( .A(n2688), .B(n2689), .Z(n2629) );
  NANDN U2748 ( .A(n17362), .B(n2488), .Z(n2490) );
  XOR U2749 ( .A(b[7]), .B(a[26]), .Z(n2652) );
  NANDN U2750 ( .A(n17522), .B(n2652), .Z(n2489) );
  AND U2751 ( .A(n2490), .B(n2489), .Z(n2715) );
  NANDN U2752 ( .A(n17072), .B(n2491), .Z(n2493) );
  XOR U2753 ( .A(b[5]), .B(a[28]), .Z(n2655) );
  NANDN U2754 ( .A(n17223), .B(n2655), .Z(n2492) );
  AND U2755 ( .A(n2493), .B(n2492), .Z(n2714) );
  NANDN U2756 ( .A(n18673), .B(n2494), .Z(n2496) );
  XOR U2757 ( .A(b[19]), .B(a[14]), .Z(n2704) );
  NANDN U2758 ( .A(n18758), .B(n2704), .Z(n2495) );
  NAND U2759 ( .A(n2496), .B(n2495), .Z(n2713) );
  XOR U2760 ( .A(n2714), .B(n2713), .Z(n2716) );
  XNOR U2761 ( .A(n2715), .B(n2716), .Z(n2628) );
  XNOR U2762 ( .A(n2629), .B(n2628), .Z(n2631) );
  NANDN U2763 ( .A(n2498), .B(n2497), .Z(n2502) );
  OR U2764 ( .A(n2500), .B(n2499), .Z(n2501) );
  AND U2765 ( .A(n2502), .B(n2501), .Z(n2630) );
  XOR U2766 ( .A(n2631), .B(n2630), .Z(n2641) );
  NANDN U2767 ( .A(n2504), .B(n2503), .Z(n2508) );
  NANDN U2768 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U2769 ( .A(n2508), .B(n2507), .Z(n2625) );
  NOR U2770 ( .A(n2510), .B(n2509), .Z(n2648) );
  NAND U2771 ( .A(n2664), .B(n2511), .Z(n2514) );
  XNOR U2772 ( .A(b[3]), .B(a[30]), .Z(n2665) );
  NANDN U2773 ( .A(n2665), .B(n2512), .Z(n2513) );
  AND U2774 ( .A(n2514), .B(n2513), .Z(n2646) );
  NAND U2775 ( .A(n18683), .B(n2515), .Z(n2517) );
  XNOR U2776 ( .A(b[17]), .B(a[16]), .Z(n2683) );
  NANDN U2777 ( .A(n2683), .B(n18684), .Z(n2516) );
  NAND U2778 ( .A(n2517), .B(n2516), .Z(n2647) );
  XOR U2779 ( .A(n2646), .B(n2647), .Z(n2649) );
  XOR U2780 ( .A(n2648), .B(n2649), .Z(n2623) );
  NANDN U2781 ( .A(n17613), .B(n2518), .Z(n2520) );
  XOR U2782 ( .A(b[9]), .B(a[24]), .Z(n2658) );
  NANDN U2783 ( .A(n17739), .B(n2658), .Z(n2519) );
  AND U2784 ( .A(n2520), .B(n2519), .Z(n2728) );
  NANDN U2785 ( .A(n19425), .B(n2521), .Z(n2523) );
  XOR U2786 ( .A(b[31]), .B(a[2]), .Z(n2680) );
  NANDN U2787 ( .A(n19426), .B(n2680), .Z(n2522) );
  AND U2788 ( .A(n2523), .B(n2522), .Z(n2726) );
  NANDN U2789 ( .A(n19005), .B(n2524), .Z(n2526) );
  XOR U2790 ( .A(b[23]), .B(a[10]), .Z(n2701) );
  NANDN U2791 ( .A(n19055), .B(n2701), .Z(n2525) );
  NAND U2792 ( .A(n2526), .B(n2525), .Z(n2725) );
  XNOR U2793 ( .A(n2726), .B(n2725), .Z(n2727) );
  XNOR U2794 ( .A(n2728), .B(n2727), .Z(n2622) );
  XNOR U2795 ( .A(n2623), .B(n2622), .Z(n2624) );
  XNOR U2796 ( .A(n2625), .B(n2624), .Z(n2640) );
  XNOR U2797 ( .A(n2641), .B(n2640), .Z(n2642) );
  XOR U2798 ( .A(n2643), .B(n2642), .Z(n2611) );
  NANDN U2799 ( .A(n2528), .B(n2527), .Z(n2532) );
  NANDN U2800 ( .A(n2530), .B(n2529), .Z(n2531) );
  AND U2801 ( .A(n2532), .B(n2531), .Z(n2610) );
  XNOR U2802 ( .A(n2611), .B(n2610), .Z(n2613) );
  NANDN U2803 ( .A(n2534), .B(n2533), .Z(n2538) );
  NANDN U2804 ( .A(n2536), .B(n2535), .Z(n2537) );
  AND U2805 ( .A(n2538), .B(n2537), .Z(n2617) );
  NANDN U2806 ( .A(n2540), .B(n2539), .Z(n2544) );
  OR U2807 ( .A(n2542), .B(n2541), .Z(n2543) );
  AND U2808 ( .A(n2544), .B(n2543), .Z(n2616) );
  XNOR U2809 ( .A(n2617), .B(n2616), .Z(n2619) );
  NANDN U2810 ( .A(n18853), .B(n2545), .Z(n2547) );
  XOR U2811 ( .A(b[21]), .B(a[12]), .Z(n2698) );
  NANDN U2812 ( .A(n18926), .B(n2698), .Z(n2546) );
  AND U2813 ( .A(n2547), .B(n2546), .Z(n2695) );
  NANDN U2814 ( .A(n2548), .B(n18439), .Z(n2550) );
  XOR U2815 ( .A(b[15]), .B(a[18]), .Z(n2707) );
  NANDN U2816 ( .A(n18311), .B(n2707), .Z(n2549) );
  AND U2817 ( .A(n2550), .B(n2549), .Z(n2693) );
  NANDN U2818 ( .A(n18113), .B(n2551), .Z(n2553) );
  XOR U2819 ( .A(b[13]), .B(a[20]), .Z(n2674) );
  NANDN U2820 ( .A(n18229), .B(n2674), .Z(n2552) );
  NAND U2821 ( .A(n2553), .B(n2552), .Z(n2692) );
  XNOR U2822 ( .A(n2693), .B(n2692), .Z(n2694) );
  XNOR U2823 ( .A(n2695), .B(n2694), .Z(n2732) );
  NAND U2824 ( .A(b[0]), .B(a[32]), .Z(n2554) );
  XNOR U2825 ( .A(b[1]), .B(n2554), .Z(n2556) );
  NANDN U2826 ( .A(b[0]), .B(a[31]), .Z(n2555) );
  NAND U2827 ( .A(n2556), .B(n2555), .Z(n2722) );
  IV U2828 ( .A(n19065), .Z(n19394) );
  NANDN U2829 ( .A(n19394), .B(n2557), .Z(n2559) );
  XOR U2830 ( .A(b[29]), .B(a[4]), .Z(n2710) );
  NANDN U2831 ( .A(n19395), .B(n2710), .Z(n2558) );
  AND U2832 ( .A(n2559), .B(n2558), .Z(n2720) );
  AND U2833 ( .A(b[31]), .B(a[0]), .Z(n2719) );
  XOR U2834 ( .A(n2720), .B(n2719), .Z(n2721) );
  XOR U2835 ( .A(n2722), .B(n2721), .Z(n2731) );
  XOR U2836 ( .A(n2732), .B(n2731), .Z(n2734) );
  NANDN U2837 ( .A(n2561), .B(n2560), .Z(n2565) );
  OR U2838 ( .A(n2563), .B(n2562), .Z(n2564) );
  NAND U2839 ( .A(n2565), .B(n2564), .Z(n2733) );
  XOR U2840 ( .A(n2734), .B(n2733), .Z(n2618) );
  XOR U2841 ( .A(n2619), .B(n2618), .Z(n2635) );
  NANDN U2842 ( .A(n2567), .B(n2566), .Z(n2571) );
  NANDN U2843 ( .A(n2569), .B(n2568), .Z(n2570) );
  AND U2844 ( .A(n2571), .B(n2570), .Z(n2634) );
  XNOR U2845 ( .A(n2635), .B(n2634), .Z(n2636) );
  NANDN U2846 ( .A(n2573), .B(n2572), .Z(n2577) );
  NANDN U2847 ( .A(n2575), .B(n2574), .Z(n2576) );
  NAND U2848 ( .A(n2577), .B(n2576), .Z(n2637) );
  XNOR U2849 ( .A(n2636), .B(n2637), .Z(n2612) );
  XOR U2850 ( .A(n2613), .B(n2612), .Z(n2740) );
  NANDN U2851 ( .A(n2579), .B(n2578), .Z(n2583) );
  NANDN U2852 ( .A(n2581), .B(n2580), .Z(n2582) );
  AND U2853 ( .A(n2583), .B(n2582), .Z(n2738) );
  NANDN U2854 ( .A(n2585), .B(n2584), .Z(n2589) );
  NAND U2855 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U2856 ( .A(n2589), .B(n2588), .Z(n2737) );
  XNOR U2857 ( .A(n2738), .B(n2737), .Z(n2739) );
  XNOR U2858 ( .A(n2740), .B(n2739), .Z(n2743) );
  XNOR U2859 ( .A(n2744), .B(n2743), .Z(n2745) );
  XOR U2860 ( .A(n2746), .B(n2745), .Z(n2605) );
  NANDN U2861 ( .A(n2591), .B(n2590), .Z(n2595) );
  NANDN U2862 ( .A(n2593), .B(n2592), .Z(n2594) );
  NAND U2863 ( .A(n2595), .B(n2594), .Z(n2604) );
  XNOR U2864 ( .A(n2605), .B(n2604), .Z(n2606) );
  XNOR U2865 ( .A(n2607), .B(n2606), .Z(n2603) );
  NANDN U2866 ( .A(n2596), .B(sreg[127]), .Z(n2600) );
  NAND U2867 ( .A(n2598), .B(n2597), .Z(n2599) );
  NAND U2868 ( .A(n2600), .B(n2599), .Z(n2602) );
  XOR U2869 ( .A(n2602), .B(sreg[128]), .Z(n2601) );
  XNOR U2870 ( .A(n2603), .B(n2601), .Z(c[128]) );
  NANDN U2871 ( .A(n2605), .B(n2604), .Z(n2609) );
  NANDN U2872 ( .A(n2607), .B(n2606), .Z(n2608) );
  AND U2873 ( .A(n2609), .B(n2608), .Z(n2752) );
  NANDN U2874 ( .A(n2611), .B(n2610), .Z(n2615) );
  NAND U2875 ( .A(n2613), .B(n2612), .Z(n2614) );
  AND U2876 ( .A(n2615), .B(n2614), .Z(n2764) );
  NANDN U2877 ( .A(n2617), .B(n2616), .Z(n2621) );
  NAND U2878 ( .A(n2619), .B(n2618), .Z(n2620) );
  AND U2879 ( .A(n2621), .B(n2620), .Z(n2775) );
  NANDN U2880 ( .A(n2623), .B(n2622), .Z(n2627) );
  NANDN U2881 ( .A(n2625), .B(n2624), .Z(n2626) );
  AND U2882 ( .A(n2627), .B(n2626), .Z(n2774) );
  NANDN U2883 ( .A(n2629), .B(n2628), .Z(n2633) );
  NAND U2884 ( .A(n2631), .B(n2630), .Z(n2632) );
  AND U2885 ( .A(n2633), .B(n2632), .Z(n2773) );
  XOR U2886 ( .A(n2774), .B(n2773), .Z(n2776) );
  XOR U2887 ( .A(n2775), .B(n2776), .Z(n2762) );
  NANDN U2888 ( .A(n2635), .B(n2634), .Z(n2639) );
  NANDN U2889 ( .A(n2637), .B(n2636), .Z(n2638) );
  NAND U2890 ( .A(n2639), .B(n2638), .Z(n2761) );
  XNOR U2891 ( .A(n2762), .B(n2761), .Z(n2763) );
  XNOR U2892 ( .A(n2764), .B(n2763), .Z(n2755) );
  NANDN U2893 ( .A(n2641), .B(n2640), .Z(n2645) );
  NAND U2894 ( .A(n2643), .B(n2642), .Z(n2644) );
  AND U2895 ( .A(n2645), .B(n2644), .Z(n2889) );
  NANDN U2896 ( .A(n2647), .B(n2646), .Z(n2651) );
  OR U2897 ( .A(n2649), .B(n2648), .Z(n2650) );
  AND U2898 ( .A(n2651), .B(n2650), .Z(n2767) );
  NANDN U2899 ( .A(n17362), .B(n2652), .Z(n2654) );
  XOR U2900 ( .A(b[7]), .B(a[27]), .Z(n2866) );
  NANDN U2901 ( .A(n17522), .B(n2866), .Z(n2653) );
  AND U2902 ( .A(n2654), .B(n2653), .Z(n2798) );
  NANDN U2903 ( .A(n17072), .B(n2655), .Z(n2657) );
  XOR U2904 ( .A(b[5]), .B(a[29]), .Z(n2815) );
  NANDN U2905 ( .A(n17223), .B(n2815), .Z(n2656) );
  NAND U2906 ( .A(n2657), .B(n2656), .Z(n2797) );
  XNOR U2907 ( .A(n2798), .B(n2797), .Z(n2800) );
  NANDN U2908 ( .A(n17613), .B(n2658), .Z(n2660) );
  XOR U2909 ( .A(b[9]), .B(a[25]), .Z(n2884) );
  NANDN U2910 ( .A(n17739), .B(n2884), .Z(n2659) );
  AND U2911 ( .A(n2660), .B(n2659), .Z(n2794) );
  NANDN U2912 ( .A(n17888), .B(n2661), .Z(n2663) );
  XOR U2913 ( .A(b[11]), .B(a[23]), .Z(n2875) );
  NANDN U2914 ( .A(n18025), .B(n2875), .Z(n2662) );
  AND U2915 ( .A(n2663), .B(n2662), .Z(n2792) );
  NANDN U2916 ( .A(n2665), .B(n2664), .Z(n2667) );
  XOR U2917 ( .A(b[3]), .B(a[31]), .Z(n2806) );
  NANDN U2918 ( .A(n17068), .B(n2806), .Z(n2666) );
  NAND U2919 ( .A(n2667), .B(n2666), .Z(n2791) );
  XNOR U2920 ( .A(n2792), .B(n2791), .Z(n2793) );
  XNOR U2921 ( .A(n2794), .B(n2793), .Z(n2799) );
  XOR U2922 ( .A(n2800), .B(n2799), .Z(n2841) );
  NANDN U2923 ( .A(n19116), .B(n2668), .Z(n2670) );
  XOR U2924 ( .A(b[25]), .B(a[9]), .Z(n2869) );
  NANDN U2925 ( .A(n19179), .B(n2869), .Z(n2669) );
  AND U2926 ( .A(n2670), .B(n2669), .Z(n2847) );
  NAND U2927 ( .A(b[0]), .B(a[33]), .Z(n2671) );
  XNOR U2928 ( .A(b[1]), .B(n2671), .Z(n2673) );
  NANDN U2929 ( .A(b[0]), .B(a[32]), .Z(n2672) );
  NAND U2930 ( .A(n2673), .B(n2672), .Z(n2846) );
  NANDN U2931 ( .A(n18113), .B(n2674), .Z(n2676) );
  XOR U2932 ( .A(b[13]), .B(a[21]), .Z(n2872) );
  NANDN U2933 ( .A(n18229), .B(n2872), .Z(n2675) );
  NAND U2934 ( .A(n2676), .B(n2675), .Z(n2845) );
  XOR U2935 ( .A(n2846), .B(n2845), .Z(n2848) );
  XOR U2936 ( .A(n2847), .B(n2848), .Z(n2840) );
  NANDN U2937 ( .A(n19237), .B(n2677), .Z(n2679) );
  XOR U2938 ( .A(b[27]), .B(a[7]), .Z(n2812) );
  NANDN U2939 ( .A(n19277), .B(n2812), .Z(n2678) );
  AND U2940 ( .A(n2679), .B(n2678), .Z(n2787) );
  NANDN U2941 ( .A(n19425), .B(n2680), .Z(n2682) );
  XOR U2942 ( .A(b[31]), .B(a[3]), .Z(n2803) );
  NANDN U2943 ( .A(n19426), .B(n2803), .Z(n2681) );
  AND U2944 ( .A(n2682), .B(n2681), .Z(n2786) );
  NANDN U2945 ( .A(n2683), .B(n18683), .Z(n2685) );
  XOR U2946 ( .A(b[17]), .B(a[17]), .Z(n2809) );
  NANDN U2947 ( .A(n18585), .B(n2809), .Z(n2684) );
  NAND U2948 ( .A(n2685), .B(n2684), .Z(n2785) );
  XOR U2949 ( .A(n2786), .B(n2785), .Z(n2788) );
  XNOR U2950 ( .A(n2787), .B(n2788), .Z(n2839) );
  XOR U2951 ( .A(n2840), .B(n2839), .Z(n2842) );
  XOR U2952 ( .A(n2841), .B(n2842), .Z(n2830) );
  NANDN U2953 ( .A(n2687), .B(n2686), .Z(n2691) );
  OR U2954 ( .A(n2689), .B(n2688), .Z(n2690) );
  AND U2955 ( .A(n2691), .B(n2690), .Z(n2828) );
  NANDN U2956 ( .A(n2693), .B(n2692), .Z(n2697) );
  NANDN U2957 ( .A(n2695), .B(n2694), .Z(n2696) );
  NAND U2958 ( .A(n2697), .B(n2696), .Z(n2827) );
  XNOR U2959 ( .A(n2828), .B(n2827), .Z(n2829) );
  XOR U2960 ( .A(n2830), .B(n2829), .Z(n2768) );
  XNOR U2961 ( .A(n2767), .B(n2768), .Z(n2770) );
  NANDN U2962 ( .A(n18853), .B(n2698), .Z(n2700) );
  XOR U2963 ( .A(b[21]), .B(a[13]), .Z(n2881) );
  NANDN U2964 ( .A(n18926), .B(n2881), .Z(n2699) );
  AND U2965 ( .A(n2700), .B(n2699), .Z(n2853) );
  NANDN U2966 ( .A(n19005), .B(n2701), .Z(n2703) );
  XOR U2967 ( .A(b[23]), .B(a[11]), .Z(n2863) );
  NANDN U2968 ( .A(n19055), .B(n2863), .Z(n2702) );
  AND U2969 ( .A(n2703), .B(n2702), .Z(n2852) );
  NANDN U2970 ( .A(n18673), .B(n2704), .Z(n2706) );
  XOR U2971 ( .A(b[19]), .B(a[15]), .Z(n2818) );
  NANDN U2972 ( .A(n18758), .B(n2818), .Z(n2705) );
  NAND U2973 ( .A(n2706), .B(n2705), .Z(n2851) );
  XOR U2974 ( .A(n2852), .B(n2851), .Z(n2854) );
  XOR U2975 ( .A(n2853), .B(n2854), .Z(n2780) );
  NANDN U2976 ( .A(n18487), .B(n2707), .Z(n2709) );
  XOR U2977 ( .A(b[15]), .B(a[19]), .Z(n2878) );
  NANDN U2978 ( .A(n18311), .B(n2878), .Z(n2708) );
  AND U2979 ( .A(n2709), .B(n2708), .Z(n2823) );
  NANDN U2980 ( .A(n19394), .B(n2710), .Z(n2712) );
  XOR U2981 ( .A(b[29]), .B(a[5]), .Z(n2860) );
  NANDN U2982 ( .A(n19395), .B(n2860), .Z(n2711) );
  AND U2983 ( .A(n2712), .B(n2711), .Z(n2822) );
  AND U2984 ( .A(b[31]), .B(a[1]), .Z(n2821) );
  XOR U2985 ( .A(n2822), .B(n2821), .Z(n2824) );
  XNOR U2986 ( .A(n2823), .B(n2824), .Z(n2779) );
  XNOR U2987 ( .A(n2780), .B(n2779), .Z(n2782) );
  NANDN U2988 ( .A(n2714), .B(n2713), .Z(n2718) );
  OR U2989 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U2990 ( .A(n2718), .B(n2717), .Z(n2781) );
  XOR U2991 ( .A(n2782), .B(n2781), .Z(n2836) );
  NANDN U2992 ( .A(n2720), .B(n2719), .Z(n2724) );
  OR U2993 ( .A(n2722), .B(n2721), .Z(n2723) );
  AND U2994 ( .A(n2724), .B(n2723), .Z(n2834) );
  NANDN U2995 ( .A(n2726), .B(n2725), .Z(n2730) );
  NANDN U2996 ( .A(n2728), .B(n2727), .Z(n2729) );
  NAND U2997 ( .A(n2730), .B(n2729), .Z(n2833) );
  XNOR U2998 ( .A(n2834), .B(n2833), .Z(n2835) );
  XNOR U2999 ( .A(n2836), .B(n2835), .Z(n2769) );
  XOR U3000 ( .A(n2770), .B(n2769), .Z(n2888) );
  NAND U3001 ( .A(n2732), .B(n2731), .Z(n2736) );
  NAND U3002 ( .A(n2734), .B(n2733), .Z(n2735) );
  AND U3003 ( .A(n2736), .B(n2735), .Z(n2887) );
  XOR U3004 ( .A(n2888), .B(n2887), .Z(n2890) );
  XOR U3005 ( .A(n2889), .B(n2890), .Z(n2756) );
  XNOR U3006 ( .A(n2755), .B(n2756), .Z(n2757) );
  NANDN U3007 ( .A(n2738), .B(n2737), .Z(n2742) );
  NANDN U3008 ( .A(n2740), .B(n2739), .Z(n2741) );
  NAND U3009 ( .A(n2742), .B(n2741), .Z(n2758) );
  XNOR U3010 ( .A(n2757), .B(n2758), .Z(n2749) );
  NANDN U3011 ( .A(n2744), .B(n2743), .Z(n2748) );
  NAND U3012 ( .A(n2746), .B(n2745), .Z(n2747) );
  NAND U3013 ( .A(n2748), .B(n2747), .Z(n2750) );
  XNOR U3014 ( .A(n2749), .B(n2750), .Z(n2751) );
  XNOR U3015 ( .A(n2752), .B(n2751), .Z(n2893) );
  XNOR U3016 ( .A(sreg[129]), .B(n2893), .Z(n2894) );
  XNOR U3017 ( .A(n2895), .B(n2894), .Z(c[129]) );
  NANDN U3018 ( .A(n2750), .B(n2749), .Z(n2754) );
  NANDN U3019 ( .A(n2752), .B(n2751), .Z(n2753) );
  AND U3020 ( .A(n2754), .B(n2753), .Z(n2901) );
  NANDN U3021 ( .A(n2756), .B(n2755), .Z(n2760) );
  NANDN U3022 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U3023 ( .A(n2760), .B(n2759), .Z(n2899) );
  NANDN U3024 ( .A(n2762), .B(n2761), .Z(n2766) );
  NANDN U3025 ( .A(n2764), .B(n2763), .Z(n2765) );
  AND U3026 ( .A(n2766), .B(n2765), .Z(n2907) );
  NANDN U3027 ( .A(n2768), .B(n2767), .Z(n2772) );
  NAND U3028 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U3029 ( .A(n2772), .B(n2771), .Z(n3037) );
  NANDN U3030 ( .A(n2774), .B(n2773), .Z(n2778) );
  OR U3031 ( .A(n2776), .B(n2775), .Z(n2777) );
  NAND U3032 ( .A(n2778), .B(n2777), .Z(n3036) );
  XNOR U3033 ( .A(n3037), .B(n3036), .Z(n3039) );
  NANDN U3034 ( .A(n2780), .B(n2779), .Z(n2784) );
  NAND U3035 ( .A(n2782), .B(n2781), .Z(n2783) );
  AND U3036 ( .A(n2784), .B(n2783), .Z(n2918) );
  NANDN U3037 ( .A(n2786), .B(n2785), .Z(n2790) );
  OR U3038 ( .A(n2788), .B(n2787), .Z(n2789) );
  AND U3039 ( .A(n2790), .B(n2789), .Z(n3024) );
  NANDN U3040 ( .A(n2792), .B(n2791), .Z(n2796) );
  NANDN U3041 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U3042 ( .A(n2796), .B(n2795), .Z(n3025) );
  XNOR U3043 ( .A(n3024), .B(n3025), .Z(n3026) );
  NANDN U3044 ( .A(n2798), .B(n2797), .Z(n2802) );
  NAND U3045 ( .A(n2800), .B(n2799), .Z(n2801) );
  NAND U3046 ( .A(n2802), .B(n2801), .Z(n3027) );
  XNOR U3047 ( .A(n3026), .B(n3027), .Z(n2916) );
  NANDN U3048 ( .A(n19425), .B(n2803), .Z(n2805) );
  XOR U3049 ( .A(b[31]), .B(a[4]), .Z(n2937) );
  NANDN U3050 ( .A(n19426), .B(n2937), .Z(n2804) );
  AND U3051 ( .A(n2805), .B(n2804), .Z(n2948) );
  NANDN U3052 ( .A(n17067), .B(n2806), .Z(n2808) );
  XOR U3053 ( .A(b[3]), .B(a[32]), .Z(n2940) );
  NANDN U3054 ( .A(n17068), .B(n2940), .Z(n2807) );
  AND U3055 ( .A(n2808), .B(n2807), .Z(n2947) );
  NANDN U3056 ( .A(n18514), .B(n2809), .Z(n2811) );
  XOR U3057 ( .A(b[17]), .B(a[18]), .Z(n2943) );
  NANDN U3058 ( .A(n18585), .B(n2943), .Z(n2810) );
  NAND U3059 ( .A(n2811), .B(n2810), .Z(n2946) );
  XOR U3060 ( .A(n2947), .B(n2946), .Z(n2949) );
  XOR U3061 ( .A(n2948), .B(n2949), .Z(n3013) );
  NANDN U3062 ( .A(n19237), .B(n2812), .Z(n2814) );
  XOR U3063 ( .A(b[27]), .B(a[8]), .Z(n2928) );
  NANDN U3064 ( .A(n19277), .B(n2928), .Z(n2813) );
  AND U3065 ( .A(n2814), .B(n2813), .Z(n2972) );
  NANDN U3066 ( .A(n17072), .B(n2815), .Z(n2817) );
  XOR U3067 ( .A(b[5]), .B(a[30]), .Z(n2931) );
  NANDN U3068 ( .A(n17223), .B(n2931), .Z(n2816) );
  AND U3069 ( .A(n2817), .B(n2816), .Z(n2971) );
  NANDN U3070 ( .A(n18673), .B(n2818), .Z(n2820) );
  XOR U3071 ( .A(b[19]), .B(a[16]), .Z(n2934) );
  NANDN U3072 ( .A(n18758), .B(n2934), .Z(n2819) );
  NAND U3073 ( .A(n2820), .B(n2819), .Z(n2970) );
  XOR U3074 ( .A(n2971), .B(n2970), .Z(n2973) );
  XNOR U3075 ( .A(n2972), .B(n2973), .Z(n3012) );
  XNOR U3076 ( .A(n3013), .B(n3012), .Z(n3014) );
  NANDN U3077 ( .A(n2822), .B(n2821), .Z(n2826) );
  OR U3078 ( .A(n2824), .B(n2823), .Z(n2825) );
  NAND U3079 ( .A(n2826), .B(n2825), .Z(n3015) );
  XOR U3080 ( .A(n3014), .B(n3015), .Z(n2917) );
  XOR U3081 ( .A(n2916), .B(n2917), .Z(n2919) );
  XOR U3082 ( .A(n2918), .B(n2919), .Z(n3033) );
  NANDN U3083 ( .A(n2828), .B(n2827), .Z(n2832) );
  NANDN U3084 ( .A(n2830), .B(n2829), .Z(n2831) );
  AND U3085 ( .A(n2832), .B(n2831), .Z(n3031) );
  NANDN U3086 ( .A(n2834), .B(n2833), .Z(n2838) );
  NANDN U3087 ( .A(n2836), .B(n2835), .Z(n2837) );
  AND U3088 ( .A(n2838), .B(n2837), .Z(n2913) );
  NANDN U3089 ( .A(n2840), .B(n2839), .Z(n2844) );
  OR U3090 ( .A(n2842), .B(n2841), .Z(n2843) );
  AND U3091 ( .A(n2844), .B(n2843), .Z(n2910) );
  NANDN U3092 ( .A(n2846), .B(n2845), .Z(n2850) );
  OR U3093 ( .A(n2848), .B(n2847), .Z(n2849) );
  AND U3094 ( .A(n2850), .B(n2849), .Z(n3019) );
  NANDN U3095 ( .A(n2852), .B(n2851), .Z(n2856) );
  OR U3096 ( .A(n2854), .B(n2853), .Z(n2855) );
  NAND U3097 ( .A(n2856), .B(n2855), .Z(n3018) );
  XNOR U3098 ( .A(n3019), .B(n3018), .Z(n3020) );
  NAND U3099 ( .A(b[0]), .B(a[34]), .Z(n2857) );
  XNOR U3100 ( .A(b[1]), .B(n2857), .Z(n2859) );
  NANDN U3101 ( .A(b[0]), .B(a[33]), .Z(n2858) );
  NAND U3102 ( .A(n2859), .B(n2858), .Z(n2925) );
  NANDN U3103 ( .A(n19394), .B(n2860), .Z(n2862) );
  XOR U3104 ( .A(b[29]), .B(a[6]), .Z(n2982) );
  NANDN U3105 ( .A(n19395), .B(n2982), .Z(n2861) );
  AND U3106 ( .A(n2862), .B(n2861), .Z(n2923) );
  AND U3107 ( .A(b[31]), .B(a[2]), .Z(n2922) );
  XNOR U3108 ( .A(n2923), .B(n2922), .Z(n2924) );
  XNOR U3109 ( .A(n2925), .B(n2924), .Z(n2964) );
  NANDN U3110 ( .A(n19005), .B(n2863), .Z(n2865) );
  XOR U3111 ( .A(b[23]), .B(a[12]), .Z(n2988) );
  NANDN U3112 ( .A(n19055), .B(n2988), .Z(n2864) );
  AND U3113 ( .A(n2865), .B(n2864), .Z(n2979) );
  NANDN U3114 ( .A(n17362), .B(n2866), .Z(n2868) );
  XOR U3115 ( .A(b[7]), .B(a[28]), .Z(n2991) );
  NANDN U3116 ( .A(n17522), .B(n2991), .Z(n2867) );
  AND U3117 ( .A(n2868), .B(n2867), .Z(n2977) );
  NANDN U3118 ( .A(n19116), .B(n2869), .Z(n2871) );
  XOR U3119 ( .A(b[25]), .B(a[10]), .Z(n2994) );
  NANDN U3120 ( .A(n19179), .B(n2994), .Z(n2870) );
  NAND U3121 ( .A(n2871), .B(n2870), .Z(n2976) );
  XNOR U3122 ( .A(n2977), .B(n2976), .Z(n2978) );
  XOR U3123 ( .A(n2979), .B(n2978), .Z(n2965) );
  XNOR U3124 ( .A(n2964), .B(n2965), .Z(n2966) );
  NANDN U3125 ( .A(n18113), .B(n2872), .Z(n2874) );
  XOR U3126 ( .A(b[13]), .B(a[22]), .Z(n2997) );
  NANDN U3127 ( .A(n18229), .B(n2997), .Z(n2873) );
  AND U3128 ( .A(n2874), .B(n2873), .Z(n2959) );
  NANDN U3129 ( .A(n17888), .B(n2875), .Z(n2877) );
  XOR U3130 ( .A(b[11]), .B(a[24]), .Z(n3000) );
  NANDN U3131 ( .A(n18025), .B(n3000), .Z(n2876) );
  NAND U3132 ( .A(n2877), .B(n2876), .Z(n2958) );
  XNOR U3133 ( .A(n2959), .B(n2958), .Z(n2960) );
  NANDN U3134 ( .A(n18487), .B(n2878), .Z(n2880) );
  XOR U3135 ( .A(b[15]), .B(a[20]), .Z(n3003) );
  NANDN U3136 ( .A(n18311), .B(n3003), .Z(n2879) );
  AND U3137 ( .A(n2880), .B(n2879), .Z(n2955) );
  NANDN U3138 ( .A(n18853), .B(n2881), .Z(n2883) );
  XOR U3139 ( .A(b[21]), .B(a[14]), .Z(n3006) );
  NANDN U3140 ( .A(n18926), .B(n3006), .Z(n2882) );
  AND U3141 ( .A(n2883), .B(n2882), .Z(n2953) );
  NANDN U3142 ( .A(n17613), .B(n2884), .Z(n2886) );
  XOR U3143 ( .A(b[9]), .B(a[26]), .Z(n3009) );
  NANDN U3144 ( .A(n17739), .B(n3009), .Z(n2885) );
  NAND U3145 ( .A(n2886), .B(n2885), .Z(n2952) );
  XNOR U3146 ( .A(n2953), .B(n2952), .Z(n2954) );
  XOR U3147 ( .A(n2955), .B(n2954), .Z(n2961) );
  XOR U3148 ( .A(n2960), .B(n2961), .Z(n2967) );
  XOR U3149 ( .A(n2966), .B(n2967), .Z(n3021) );
  XOR U3150 ( .A(n3020), .B(n3021), .Z(n2911) );
  XNOR U3151 ( .A(n2910), .B(n2911), .Z(n2912) );
  XNOR U3152 ( .A(n2913), .B(n2912), .Z(n3030) );
  XNOR U3153 ( .A(n3031), .B(n3030), .Z(n3032) );
  XNOR U3154 ( .A(n3033), .B(n3032), .Z(n3038) );
  XOR U3155 ( .A(n3039), .B(n3038), .Z(n2905) );
  NANDN U3156 ( .A(n2888), .B(n2887), .Z(n2892) );
  NANDN U3157 ( .A(n2890), .B(n2889), .Z(n2891) );
  NAND U3158 ( .A(n2892), .B(n2891), .Z(n2904) );
  XNOR U3159 ( .A(n2905), .B(n2904), .Z(n2906) );
  XNOR U3160 ( .A(n2907), .B(n2906), .Z(n2898) );
  XNOR U3161 ( .A(n2899), .B(n2898), .Z(n2900) );
  XNOR U3162 ( .A(n2901), .B(n2900), .Z(n3042) );
  XNOR U3163 ( .A(sreg[130]), .B(n3042), .Z(n3044) );
  NANDN U3164 ( .A(sreg[129]), .B(n2893), .Z(n2897) );
  NAND U3165 ( .A(n2895), .B(n2894), .Z(n2896) );
  NAND U3166 ( .A(n2897), .B(n2896), .Z(n3043) );
  XNOR U3167 ( .A(n3044), .B(n3043), .Z(c[130]) );
  NANDN U3168 ( .A(n2899), .B(n2898), .Z(n2903) );
  NANDN U3169 ( .A(n2901), .B(n2900), .Z(n2902) );
  AND U3170 ( .A(n2903), .B(n2902), .Z(n3052) );
  NANDN U3171 ( .A(n2905), .B(n2904), .Z(n2909) );
  NANDN U3172 ( .A(n2907), .B(n2906), .Z(n2908) );
  AND U3173 ( .A(n2909), .B(n2908), .Z(n3051) );
  NANDN U3174 ( .A(n2911), .B(n2910), .Z(n2915) );
  NANDN U3175 ( .A(n2913), .B(n2912), .Z(n2914) );
  AND U3176 ( .A(n2915), .B(n2914), .Z(n3189) );
  NANDN U3177 ( .A(n2917), .B(n2916), .Z(n2921) );
  OR U3178 ( .A(n2919), .B(n2918), .Z(n2920) );
  AND U3179 ( .A(n2921), .B(n2920), .Z(n3188) );
  XNOR U3180 ( .A(n3189), .B(n3188), .Z(n3191) );
  NANDN U3181 ( .A(n2923), .B(n2922), .Z(n2927) );
  NANDN U3182 ( .A(n2925), .B(n2924), .Z(n2926) );
  AND U3183 ( .A(n2927), .B(n2926), .Z(n3136) );
  NANDN U3184 ( .A(n19237), .B(n2928), .Z(n2930) );
  XOR U3185 ( .A(b[27]), .B(a[9]), .Z(n3080) );
  NANDN U3186 ( .A(n19277), .B(n3080), .Z(n2929) );
  AND U3187 ( .A(n2930), .B(n2929), .Z(n3143) );
  NANDN U3188 ( .A(n17072), .B(n2931), .Z(n2933) );
  XOR U3189 ( .A(b[5]), .B(a[31]), .Z(n3083) );
  NANDN U3190 ( .A(n17223), .B(n3083), .Z(n2932) );
  AND U3191 ( .A(n2933), .B(n2932), .Z(n3141) );
  NANDN U3192 ( .A(n18673), .B(n2934), .Z(n2936) );
  XOR U3193 ( .A(b[19]), .B(a[17]), .Z(n3086) );
  NANDN U3194 ( .A(n18758), .B(n3086), .Z(n2935) );
  NAND U3195 ( .A(n2936), .B(n2935), .Z(n3140) );
  XNOR U3196 ( .A(n3141), .B(n3140), .Z(n3142) );
  XNOR U3197 ( .A(n3143), .B(n3142), .Z(n3134) );
  NANDN U3198 ( .A(n19425), .B(n2937), .Z(n2939) );
  XOR U3199 ( .A(b[31]), .B(a[5]), .Z(n3089) );
  NANDN U3200 ( .A(n19426), .B(n3089), .Z(n2938) );
  AND U3201 ( .A(n2939), .B(n2938), .Z(n3101) );
  NANDN U3202 ( .A(n17067), .B(n2940), .Z(n2942) );
  XOR U3203 ( .A(b[3]), .B(a[33]), .Z(n3092) );
  NANDN U3204 ( .A(n17068), .B(n3092), .Z(n2941) );
  AND U3205 ( .A(n2942), .B(n2941), .Z(n3099) );
  NANDN U3206 ( .A(n18514), .B(n2943), .Z(n2945) );
  XOR U3207 ( .A(b[17]), .B(a[19]), .Z(n3095) );
  NANDN U3208 ( .A(n18585), .B(n3095), .Z(n2944) );
  NAND U3209 ( .A(n2945), .B(n2944), .Z(n3098) );
  XNOR U3210 ( .A(n3099), .B(n3098), .Z(n3100) );
  XOR U3211 ( .A(n3101), .B(n3100), .Z(n3135) );
  XOR U3212 ( .A(n3134), .B(n3135), .Z(n3137) );
  XOR U3213 ( .A(n3136), .B(n3137), .Z(n3063) );
  NANDN U3214 ( .A(n2947), .B(n2946), .Z(n2951) );
  OR U3215 ( .A(n2949), .B(n2948), .Z(n2950) );
  AND U3216 ( .A(n2951), .B(n2950), .Z(n3122) );
  NANDN U3217 ( .A(n2953), .B(n2952), .Z(n2957) );
  NANDN U3218 ( .A(n2955), .B(n2954), .Z(n2956) );
  NAND U3219 ( .A(n2957), .B(n2956), .Z(n3123) );
  XNOR U3220 ( .A(n3122), .B(n3123), .Z(n3124) );
  NANDN U3221 ( .A(n2959), .B(n2958), .Z(n2963) );
  NANDN U3222 ( .A(n2961), .B(n2960), .Z(n2962) );
  NAND U3223 ( .A(n2963), .B(n2962), .Z(n3125) );
  XNOR U3224 ( .A(n3124), .B(n3125), .Z(n3062) );
  XNOR U3225 ( .A(n3063), .B(n3062), .Z(n3065) );
  NANDN U3226 ( .A(n2965), .B(n2964), .Z(n2969) );
  NANDN U3227 ( .A(n2967), .B(n2966), .Z(n2968) );
  AND U3228 ( .A(n2969), .B(n2968), .Z(n3064) );
  XOR U3229 ( .A(n3065), .B(n3064), .Z(n3185) );
  NANDN U3230 ( .A(n2971), .B(n2970), .Z(n2975) );
  OR U3231 ( .A(n2973), .B(n2972), .Z(n2974) );
  AND U3232 ( .A(n2975), .B(n2974), .Z(n3129) );
  NANDN U3233 ( .A(n2977), .B(n2976), .Z(n2981) );
  NANDN U3234 ( .A(n2979), .B(n2978), .Z(n2980) );
  NAND U3235 ( .A(n2981), .B(n2980), .Z(n3128) );
  XNOR U3236 ( .A(n3129), .B(n3128), .Z(n3131) );
  NANDN U3237 ( .A(n19394), .B(n2982), .Z(n2984) );
  XOR U3238 ( .A(b[29]), .B(a[7]), .Z(n3155) );
  NANDN U3239 ( .A(n19395), .B(n3155), .Z(n2983) );
  AND U3240 ( .A(n2984), .B(n2983), .Z(n3075) );
  AND U3241 ( .A(b[31]), .B(a[3]), .Z(n3074) );
  XNOR U3242 ( .A(n3075), .B(n3074), .Z(n3076) );
  NAND U3243 ( .A(b[0]), .B(a[35]), .Z(n2985) );
  XNOR U3244 ( .A(b[1]), .B(n2985), .Z(n2987) );
  NANDN U3245 ( .A(b[0]), .B(a[34]), .Z(n2986) );
  NAND U3246 ( .A(n2987), .B(n2986), .Z(n3077) );
  XNOR U3247 ( .A(n3076), .B(n3077), .Z(n3116) );
  NANDN U3248 ( .A(n19005), .B(n2988), .Z(n2990) );
  XOR U3249 ( .A(b[23]), .B(a[13]), .Z(n3158) );
  NANDN U3250 ( .A(n19055), .B(n3158), .Z(n2989) );
  AND U3251 ( .A(n2990), .B(n2989), .Z(n3149) );
  NANDN U3252 ( .A(n17362), .B(n2991), .Z(n2993) );
  XOR U3253 ( .A(b[7]), .B(a[29]), .Z(n3161) );
  NANDN U3254 ( .A(n17522), .B(n3161), .Z(n2992) );
  AND U3255 ( .A(n2993), .B(n2992), .Z(n3147) );
  NANDN U3256 ( .A(n19116), .B(n2994), .Z(n2996) );
  XOR U3257 ( .A(b[25]), .B(a[11]), .Z(n3164) );
  NANDN U3258 ( .A(n19179), .B(n3164), .Z(n2995) );
  NAND U3259 ( .A(n2996), .B(n2995), .Z(n3146) );
  XNOR U3260 ( .A(n3147), .B(n3146), .Z(n3148) );
  XOR U3261 ( .A(n3149), .B(n3148), .Z(n3117) );
  XNOR U3262 ( .A(n3116), .B(n3117), .Z(n3118) );
  NANDN U3263 ( .A(n18113), .B(n2997), .Z(n2999) );
  XOR U3264 ( .A(b[13]), .B(a[23]), .Z(n3167) );
  NANDN U3265 ( .A(n18229), .B(n3167), .Z(n2998) );
  AND U3266 ( .A(n2999), .B(n2998), .Z(n3111) );
  NANDN U3267 ( .A(n17888), .B(n3000), .Z(n3002) );
  XOR U3268 ( .A(b[11]), .B(a[25]), .Z(n3170) );
  NANDN U3269 ( .A(n18025), .B(n3170), .Z(n3001) );
  NAND U3270 ( .A(n3002), .B(n3001), .Z(n3110) );
  XNOR U3271 ( .A(n3111), .B(n3110), .Z(n3112) );
  NANDN U3272 ( .A(n18487), .B(n3003), .Z(n3005) );
  XOR U3273 ( .A(b[15]), .B(a[21]), .Z(n3173) );
  NANDN U3274 ( .A(n18311), .B(n3173), .Z(n3004) );
  AND U3275 ( .A(n3005), .B(n3004), .Z(n3107) );
  NANDN U3276 ( .A(n18853), .B(n3006), .Z(n3008) );
  XOR U3277 ( .A(b[21]), .B(a[15]), .Z(n3176) );
  NANDN U3278 ( .A(n18926), .B(n3176), .Z(n3007) );
  AND U3279 ( .A(n3008), .B(n3007), .Z(n3105) );
  NANDN U3280 ( .A(n17613), .B(n3009), .Z(n3011) );
  XOR U3281 ( .A(b[9]), .B(a[27]), .Z(n3179) );
  NANDN U3282 ( .A(n17739), .B(n3179), .Z(n3010) );
  NAND U3283 ( .A(n3011), .B(n3010), .Z(n3104) );
  XNOR U3284 ( .A(n3105), .B(n3104), .Z(n3106) );
  XOR U3285 ( .A(n3107), .B(n3106), .Z(n3113) );
  XOR U3286 ( .A(n3112), .B(n3113), .Z(n3119) );
  XNOR U3287 ( .A(n3118), .B(n3119), .Z(n3130) );
  XOR U3288 ( .A(n3131), .B(n3130), .Z(n3069) );
  NANDN U3289 ( .A(n3013), .B(n3012), .Z(n3017) );
  NANDN U3290 ( .A(n3015), .B(n3014), .Z(n3016) );
  NAND U3291 ( .A(n3017), .B(n3016), .Z(n3068) );
  XNOR U3292 ( .A(n3069), .B(n3068), .Z(n3071) );
  NANDN U3293 ( .A(n3019), .B(n3018), .Z(n3023) );
  NANDN U3294 ( .A(n3021), .B(n3020), .Z(n3022) );
  AND U3295 ( .A(n3023), .B(n3022), .Z(n3070) );
  XOR U3296 ( .A(n3071), .B(n3070), .Z(n3183) );
  NANDN U3297 ( .A(n3025), .B(n3024), .Z(n3029) );
  NANDN U3298 ( .A(n3027), .B(n3026), .Z(n3028) );
  AND U3299 ( .A(n3029), .B(n3028), .Z(n3182) );
  XNOR U3300 ( .A(n3183), .B(n3182), .Z(n3184) );
  XNOR U3301 ( .A(n3185), .B(n3184), .Z(n3190) );
  XOR U3302 ( .A(n3191), .B(n3190), .Z(n3057) );
  NANDN U3303 ( .A(n3031), .B(n3030), .Z(n3035) );
  NANDN U3304 ( .A(n3033), .B(n3032), .Z(n3034) );
  AND U3305 ( .A(n3035), .B(n3034), .Z(n3056) );
  XNOR U3306 ( .A(n3057), .B(n3056), .Z(n3058) );
  NANDN U3307 ( .A(n3037), .B(n3036), .Z(n3041) );
  NAND U3308 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U3309 ( .A(n3041), .B(n3040), .Z(n3059) );
  XNOR U3310 ( .A(n3058), .B(n3059), .Z(n3050) );
  XOR U3311 ( .A(n3051), .B(n3050), .Z(n3053) );
  XOR U3312 ( .A(n3052), .B(n3053), .Z(n3048) );
  NANDN U3313 ( .A(sreg[130]), .B(n3042), .Z(n3046) );
  NAND U3314 ( .A(n3044), .B(n3043), .Z(n3045) );
  AND U3315 ( .A(n3046), .B(n3045), .Z(n3049) );
  XNOR U3316 ( .A(sreg[131]), .B(n3049), .Z(n3047) );
  XOR U3317 ( .A(n3048), .B(n3047), .Z(c[131]) );
  NANDN U3318 ( .A(n3051), .B(n3050), .Z(n3055) );
  OR U3319 ( .A(n3053), .B(n3052), .Z(n3054) );
  AND U3320 ( .A(n3055), .B(n3054), .Z(n3197) );
  NANDN U3321 ( .A(n3057), .B(n3056), .Z(n3061) );
  NANDN U3322 ( .A(n3059), .B(n3058), .Z(n3060) );
  AND U3323 ( .A(n3061), .B(n3060), .Z(n3195) );
  NANDN U3324 ( .A(n3063), .B(n3062), .Z(n3067) );
  NAND U3325 ( .A(n3065), .B(n3064), .Z(n3066) );
  AND U3326 ( .A(n3067), .B(n3066), .Z(n3332) );
  NANDN U3327 ( .A(n3069), .B(n3068), .Z(n3073) );
  NAND U3328 ( .A(n3071), .B(n3070), .Z(n3072) );
  NAND U3329 ( .A(n3073), .B(n3072), .Z(n3333) );
  XNOR U3330 ( .A(n3332), .B(n3333), .Z(n3335) );
  NANDN U3331 ( .A(n3075), .B(n3074), .Z(n3079) );
  NANDN U3332 ( .A(n3077), .B(n3076), .Z(n3078) );
  AND U3333 ( .A(n3079), .B(n3078), .Z(n3280) );
  NANDN U3334 ( .A(n19237), .B(n3080), .Z(n3082) );
  XOR U3335 ( .A(b[27]), .B(a[10]), .Z(n3224) );
  NANDN U3336 ( .A(n19277), .B(n3224), .Z(n3081) );
  AND U3337 ( .A(n3082), .B(n3081), .Z(n3287) );
  NANDN U3338 ( .A(n17072), .B(n3083), .Z(n3085) );
  XOR U3339 ( .A(b[5]), .B(a[32]), .Z(n3227) );
  NANDN U3340 ( .A(n17223), .B(n3227), .Z(n3084) );
  AND U3341 ( .A(n3085), .B(n3084), .Z(n3285) );
  NANDN U3342 ( .A(n18673), .B(n3086), .Z(n3088) );
  XOR U3343 ( .A(b[19]), .B(a[18]), .Z(n3230) );
  NANDN U3344 ( .A(n18758), .B(n3230), .Z(n3087) );
  NAND U3345 ( .A(n3088), .B(n3087), .Z(n3284) );
  XNOR U3346 ( .A(n3285), .B(n3284), .Z(n3286) );
  XNOR U3347 ( .A(n3287), .B(n3286), .Z(n3278) );
  NANDN U3348 ( .A(n19425), .B(n3089), .Z(n3091) );
  XOR U3349 ( .A(b[31]), .B(a[6]), .Z(n3233) );
  NANDN U3350 ( .A(n19426), .B(n3233), .Z(n3090) );
  AND U3351 ( .A(n3091), .B(n3090), .Z(n3245) );
  NANDN U3352 ( .A(n17067), .B(n3092), .Z(n3094) );
  XOR U3353 ( .A(b[3]), .B(a[34]), .Z(n3236) );
  NANDN U3354 ( .A(n17068), .B(n3236), .Z(n3093) );
  AND U3355 ( .A(n3094), .B(n3093), .Z(n3243) );
  NANDN U3356 ( .A(n18514), .B(n3095), .Z(n3097) );
  XOR U3357 ( .A(b[17]), .B(a[20]), .Z(n3239) );
  NANDN U3358 ( .A(n18585), .B(n3239), .Z(n3096) );
  NAND U3359 ( .A(n3097), .B(n3096), .Z(n3242) );
  XNOR U3360 ( .A(n3243), .B(n3242), .Z(n3244) );
  XOR U3361 ( .A(n3245), .B(n3244), .Z(n3279) );
  XOR U3362 ( .A(n3278), .B(n3279), .Z(n3281) );
  XOR U3363 ( .A(n3280), .B(n3281), .Z(n3213) );
  NANDN U3364 ( .A(n3099), .B(n3098), .Z(n3103) );
  NANDN U3365 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3366 ( .A(n3103), .B(n3102), .Z(n3266) );
  NANDN U3367 ( .A(n3105), .B(n3104), .Z(n3109) );
  NANDN U3368 ( .A(n3107), .B(n3106), .Z(n3108) );
  NAND U3369 ( .A(n3109), .B(n3108), .Z(n3267) );
  XNOR U3370 ( .A(n3266), .B(n3267), .Z(n3268) );
  NANDN U3371 ( .A(n3111), .B(n3110), .Z(n3115) );
  NANDN U3372 ( .A(n3113), .B(n3112), .Z(n3114) );
  NAND U3373 ( .A(n3115), .B(n3114), .Z(n3269) );
  XNOR U3374 ( .A(n3268), .B(n3269), .Z(n3212) );
  XNOR U3375 ( .A(n3213), .B(n3212), .Z(n3215) );
  NANDN U3376 ( .A(n3117), .B(n3116), .Z(n3121) );
  NANDN U3377 ( .A(n3119), .B(n3118), .Z(n3120) );
  AND U3378 ( .A(n3121), .B(n3120), .Z(n3214) );
  XOR U3379 ( .A(n3215), .B(n3214), .Z(n3329) );
  NANDN U3380 ( .A(n3123), .B(n3122), .Z(n3127) );
  NANDN U3381 ( .A(n3125), .B(n3124), .Z(n3126) );
  AND U3382 ( .A(n3127), .B(n3126), .Z(n3326) );
  NANDN U3383 ( .A(n3129), .B(n3128), .Z(n3133) );
  NAND U3384 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U3385 ( .A(n3133), .B(n3132), .Z(n3209) );
  NANDN U3386 ( .A(n3135), .B(n3134), .Z(n3139) );
  OR U3387 ( .A(n3137), .B(n3136), .Z(n3138) );
  AND U3388 ( .A(n3139), .B(n3138), .Z(n3207) );
  NANDN U3389 ( .A(n3141), .B(n3140), .Z(n3145) );
  NANDN U3390 ( .A(n3143), .B(n3142), .Z(n3144) );
  AND U3391 ( .A(n3145), .B(n3144), .Z(n3273) );
  NANDN U3392 ( .A(n3147), .B(n3146), .Z(n3151) );
  NANDN U3393 ( .A(n3149), .B(n3148), .Z(n3150) );
  NAND U3394 ( .A(n3151), .B(n3150), .Z(n3272) );
  XNOR U3395 ( .A(n3273), .B(n3272), .Z(n3274) );
  NAND U3396 ( .A(b[0]), .B(a[36]), .Z(n3152) );
  XNOR U3397 ( .A(b[1]), .B(n3152), .Z(n3154) );
  NANDN U3398 ( .A(b[0]), .B(a[35]), .Z(n3153) );
  NAND U3399 ( .A(n3154), .B(n3153), .Z(n3221) );
  NANDN U3400 ( .A(n19394), .B(n3155), .Z(n3157) );
  XOR U3401 ( .A(b[29]), .B(a[8]), .Z(n3299) );
  NANDN U3402 ( .A(n19395), .B(n3299), .Z(n3156) );
  AND U3403 ( .A(n3157), .B(n3156), .Z(n3219) );
  AND U3404 ( .A(b[31]), .B(a[4]), .Z(n3218) );
  XNOR U3405 ( .A(n3219), .B(n3218), .Z(n3220) );
  XNOR U3406 ( .A(n3221), .B(n3220), .Z(n3260) );
  NANDN U3407 ( .A(n19005), .B(n3158), .Z(n3160) );
  XOR U3408 ( .A(b[23]), .B(a[14]), .Z(n3302) );
  NANDN U3409 ( .A(n19055), .B(n3302), .Z(n3159) );
  AND U3410 ( .A(n3160), .B(n3159), .Z(n3293) );
  NANDN U3411 ( .A(n17362), .B(n3161), .Z(n3163) );
  XOR U3412 ( .A(b[7]), .B(a[30]), .Z(n3305) );
  NANDN U3413 ( .A(n17522), .B(n3305), .Z(n3162) );
  AND U3414 ( .A(n3163), .B(n3162), .Z(n3291) );
  NANDN U3415 ( .A(n19116), .B(n3164), .Z(n3166) );
  XOR U3416 ( .A(b[25]), .B(a[12]), .Z(n3308) );
  NANDN U3417 ( .A(n19179), .B(n3308), .Z(n3165) );
  NAND U3418 ( .A(n3166), .B(n3165), .Z(n3290) );
  XNOR U3419 ( .A(n3291), .B(n3290), .Z(n3292) );
  XOR U3420 ( .A(n3293), .B(n3292), .Z(n3261) );
  XNOR U3421 ( .A(n3260), .B(n3261), .Z(n3262) );
  NANDN U3422 ( .A(n18113), .B(n3167), .Z(n3169) );
  XOR U3423 ( .A(b[13]), .B(a[24]), .Z(n3311) );
  NANDN U3424 ( .A(n18229), .B(n3311), .Z(n3168) );
  AND U3425 ( .A(n3169), .B(n3168), .Z(n3255) );
  NANDN U3426 ( .A(n17888), .B(n3170), .Z(n3172) );
  XOR U3427 ( .A(b[11]), .B(a[26]), .Z(n3314) );
  NANDN U3428 ( .A(n18025), .B(n3314), .Z(n3171) );
  NAND U3429 ( .A(n3172), .B(n3171), .Z(n3254) );
  XNOR U3430 ( .A(n3255), .B(n3254), .Z(n3256) );
  NANDN U3431 ( .A(n18487), .B(n3173), .Z(n3175) );
  XOR U3432 ( .A(b[15]), .B(a[22]), .Z(n3317) );
  NANDN U3433 ( .A(n18311), .B(n3317), .Z(n3174) );
  AND U3434 ( .A(n3175), .B(n3174), .Z(n3251) );
  NANDN U3435 ( .A(n18853), .B(n3176), .Z(n3178) );
  XOR U3436 ( .A(b[21]), .B(a[16]), .Z(n3320) );
  NANDN U3437 ( .A(n18926), .B(n3320), .Z(n3177) );
  AND U3438 ( .A(n3178), .B(n3177), .Z(n3249) );
  NANDN U3439 ( .A(n17613), .B(n3179), .Z(n3181) );
  XOR U3440 ( .A(b[9]), .B(a[28]), .Z(n3323) );
  NANDN U3441 ( .A(n17739), .B(n3323), .Z(n3180) );
  NAND U3442 ( .A(n3181), .B(n3180), .Z(n3248) );
  XNOR U3443 ( .A(n3249), .B(n3248), .Z(n3250) );
  XOR U3444 ( .A(n3251), .B(n3250), .Z(n3257) );
  XOR U3445 ( .A(n3256), .B(n3257), .Z(n3263) );
  XOR U3446 ( .A(n3262), .B(n3263), .Z(n3275) );
  XNOR U3447 ( .A(n3274), .B(n3275), .Z(n3206) );
  XNOR U3448 ( .A(n3207), .B(n3206), .Z(n3208) );
  XOR U3449 ( .A(n3209), .B(n3208), .Z(n3327) );
  XNOR U3450 ( .A(n3326), .B(n3327), .Z(n3328) );
  XNOR U3451 ( .A(n3329), .B(n3328), .Z(n3334) );
  XOR U3452 ( .A(n3335), .B(n3334), .Z(n3201) );
  NANDN U3453 ( .A(n3183), .B(n3182), .Z(n3187) );
  NANDN U3454 ( .A(n3185), .B(n3184), .Z(n3186) );
  AND U3455 ( .A(n3187), .B(n3186), .Z(n3200) );
  XNOR U3456 ( .A(n3201), .B(n3200), .Z(n3202) );
  NANDN U3457 ( .A(n3189), .B(n3188), .Z(n3193) );
  NAND U3458 ( .A(n3191), .B(n3190), .Z(n3192) );
  NAND U3459 ( .A(n3193), .B(n3192), .Z(n3203) );
  XNOR U3460 ( .A(n3202), .B(n3203), .Z(n3194) );
  XNOR U3461 ( .A(n3195), .B(n3194), .Z(n3196) );
  XNOR U3462 ( .A(n3197), .B(n3196), .Z(n3338) );
  XNOR U3463 ( .A(sreg[132]), .B(n3338), .Z(n3339) );
  XOR U3464 ( .A(n3340), .B(n3339), .Z(c[132]) );
  NANDN U3465 ( .A(n3195), .B(n3194), .Z(n3199) );
  NANDN U3466 ( .A(n3197), .B(n3196), .Z(n3198) );
  AND U3467 ( .A(n3199), .B(n3198), .Z(n3346) );
  NANDN U3468 ( .A(n3201), .B(n3200), .Z(n3205) );
  NANDN U3469 ( .A(n3203), .B(n3202), .Z(n3204) );
  AND U3470 ( .A(n3205), .B(n3204), .Z(n3344) );
  NANDN U3471 ( .A(n3207), .B(n3206), .Z(n3211) );
  NANDN U3472 ( .A(n3209), .B(n3208), .Z(n3210) );
  AND U3473 ( .A(n3211), .B(n3210), .Z(n3356) );
  NANDN U3474 ( .A(n3213), .B(n3212), .Z(n3217) );
  NAND U3475 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U3476 ( .A(n3217), .B(n3216), .Z(n3355) );
  XNOR U3477 ( .A(n3356), .B(n3355), .Z(n3358) );
  NANDN U3478 ( .A(n3219), .B(n3218), .Z(n3223) );
  NANDN U3479 ( .A(n3221), .B(n3220), .Z(n3222) );
  AND U3480 ( .A(n3223), .B(n3222), .Z(n3435) );
  NANDN U3481 ( .A(n19237), .B(n3224), .Z(n3226) );
  XOR U3482 ( .A(b[27]), .B(a[11]), .Z(n3379) );
  NANDN U3483 ( .A(n19277), .B(n3379), .Z(n3225) );
  AND U3484 ( .A(n3226), .B(n3225), .Z(n3442) );
  NANDN U3485 ( .A(n17072), .B(n3227), .Z(n3229) );
  XOR U3486 ( .A(b[5]), .B(a[33]), .Z(n3382) );
  NANDN U3487 ( .A(n17223), .B(n3382), .Z(n3228) );
  AND U3488 ( .A(n3229), .B(n3228), .Z(n3440) );
  NANDN U3489 ( .A(n18673), .B(n3230), .Z(n3232) );
  XOR U3490 ( .A(b[19]), .B(a[19]), .Z(n3385) );
  NANDN U3491 ( .A(n18758), .B(n3385), .Z(n3231) );
  NAND U3492 ( .A(n3232), .B(n3231), .Z(n3439) );
  XNOR U3493 ( .A(n3440), .B(n3439), .Z(n3441) );
  XNOR U3494 ( .A(n3442), .B(n3441), .Z(n3433) );
  NANDN U3495 ( .A(n19425), .B(n3233), .Z(n3235) );
  XOR U3496 ( .A(b[31]), .B(a[7]), .Z(n3388) );
  NANDN U3497 ( .A(n19426), .B(n3388), .Z(n3234) );
  AND U3498 ( .A(n3235), .B(n3234), .Z(n3400) );
  NANDN U3499 ( .A(n17067), .B(n3236), .Z(n3238) );
  XOR U3500 ( .A(b[3]), .B(a[35]), .Z(n3391) );
  NANDN U3501 ( .A(n17068), .B(n3391), .Z(n3237) );
  AND U3502 ( .A(n3238), .B(n3237), .Z(n3398) );
  NANDN U3503 ( .A(n18514), .B(n3239), .Z(n3241) );
  XOR U3504 ( .A(b[17]), .B(a[21]), .Z(n3394) );
  NANDN U3505 ( .A(n18585), .B(n3394), .Z(n3240) );
  NAND U3506 ( .A(n3241), .B(n3240), .Z(n3397) );
  XNOR U3507 ( .A(n3398), .B(n3397), .Z(n3399) );
  XOR U3508 ( .A(n3400), .B(n3399), .Z(n3434) );
  XOR U3509 ( .A(n3433), .B(n3434), .Z(n3436) );
  XOR U3510 ( .A(n3435), .B(n3436), .Z(n3368) );
  NANDN U3511 ( .A(n3243), .B(n3242), .Z(n3247) );
  NANDN U3512 ( .A(n3245), .B(n3244), .Z(n3246) );
  AND U3513 ( .A(n3247), .B(n3246), .Z(n3421) );
  NANDN U3514 ( .A(n3249), .B(n3248), .Z(n3253) );
  NANDN U3515 ( .A(n3251), .B(n3250), .Z(n3252) );
  NAND U3516 ( .A(n3253), .B(n3252), .Z(n3422) );
  XNOR U3517 ( .A(n3421), .B(n3422), .Z(n3423) );
  NANDN U3518 ( .A(n3255), .B(n3254), .Z(n3259) );
  NANDN U3519 ( .A(n3257), .B(n3256), .Z(n3258) );
  NAND U3520 ( .A(n3259), .B(n3258), .Z(n3424) );
  XNOR U3521 ( .A(n3423), .B(n3424), .Z(n3367) );
  XNOR U3522 ( .A(n3368), .B(n3367), .Z(n3370) );
  NANDN U3523 ( .A(n3261), .B(n3260), .Z(n3265) );
  NANDN U3524 ( .A(n3263), .B(n3262), .Z(n3264) );
  AND U3525 ( .A(n3265), .B(n3264), .Z(n3369) );
  XOR U3526 ( .A(n3370), .B(n3369), .Z(n3484) );
  NANDN U3527 ( .A(n3267), .B(n3266), .Z(n3271) );
  NANDN U3528 ( .A(n3269), .B(n3268), .Z(n3270) );
  AND U3529 ( .A(n3271), .B(n3270), .Z(n3481) );
  NANDN U3530 ( .A(n3273), .B(n3272), .Z(n3277) );
  NANDN U3531 ( .A(n3275), .B(n3274), .Z(n3276) );
  AND U3532 ( .A(n3277), .B(n3276), .Z(n3364) );
  NANDN U3533 ( .A(n3279), .B(n3278), .Z(n3283) );
  OR U3534 ( .A(n3281), .B(n3280), .Z(n3282) );
  AND U3535 ( .A(n3283), .B(n3282), .Z(n3362) );
  NANDN U3536 ( .A(n3285), .B(n3284), .Z(n3289) );
  NANDN U3537 ( .A(n3287), .B(n3286), .Z(n3288) );
  AND U3538 ( .A(n3289), .B(n3288), .Z(n3428) );
  NANDN U3539 ( .A(n3291), .B(n3290), .Z(n3295) );
  NANDN U3540 ( .A(n3293), .B(n3292), .Z(n3294) );
  NAND U3541 ( .A(n3295), .B(n3294), .Z(n3427) );
  XNOR U3542 ( .A(n3428), .B(n3427), .Z(n3429) );
  NAND U3543 ( .A(b[0]), .B(a[37]), .Z(n3296) );
  XNOR U3544 ( .A(b[1]), .B(n3296), .Z(n3298) );
  NANDN U3545 ( .A(b[0]), .B(a[36]), .Z(n3297) );
  NAND U3546 ( .A(n3298), .B(n3297), .Z(n3376) );
  NANDN U3547 ( .A(n19394), .B(n3299), .Z(n3301) );
  XOR U3548 ( .A(b[29]), .B(a[9]), .Z(n3454) );
  NANDN U3549 ( .A(n19395), .B(n3454), .Z(n3300) );
  AND U3550 ( .A(n3301), .B(n3300), .Z(n3374) );
  AND U3551 ( .A(b[31]), .B(a[5]), .Z(n3373) );
  XNOR U3552 ( .A(n3374), .B(n3373), .Z(n3375) );
  XNOR U3553 ( .A(n3376), .B(n3375), .Z(n3415) );
  NANDN U3554 ( .A(n19005), .B(n3302), .Z(n3304) );
  XOR U3555 ( .A(b[23]), .B(a[15]), .Z(n3457) );
  NANDN U3556 ( .A(n19055), .B(n3457), .Z(n3303) );
  AND U3557 ( .A(n3304), .B(n3303), .Z(n3448) );
  NANDN U3558 ( .A(n17362), .B(n3305), .Z(n3307) );
  XOR U3559 ( .A(b[7]), .B(a[31]), .Z(n3460) );
  NANDN U3560 ( .A(n17522), .B(n3460), .Z(n3306) );
  AND U3561 ( .A(n3307), .B(n3306), .Z(n3446) );
  NANDN U3562 ( .A(n19116), .B(n3308), .Z(n3310) );
  XOR U3563 ( .A(b[25]), .B(a[13]), .Z(n3463) );
  NANDN U3564 ( .A(n19179), .B(n3463), .Z(n3309) );
  NAND U3565 ( .A(n3310), .B(n3309), .Z(n3445) );
  XNOR U3566 ( .A(n3446), .B(n3445), .Z(n3447) );
  XOR U3567 ( .A(n3448), .B(n3447), .Z(n3416) );
  XNOR U3568 ( .A(n3415), .B(n3416), .Z(n3417) );
  NANDN U3569 ( .A(n18113), .B(n3311), .Z(n3313) );
  XOR U3570 ( .A(b[13]), .B(a[25]), .Z(n3466) );
  NANDN U3571 ( .A(n18229), .B(n3466), .Z(n3312) );
  AND U3572 ( .A(n3313), .B(n3312), .Z(n3410) );
  NANDN U3573 ( .A(n17888), .B(n3314), .Z(n3316) );
  XOR U3574 ( .A(b[11]), .B(a[27]), .Z(n3469) );
  NANDN U3575 ( .A(n18025), .B(n3469), .Z(n3315) );
  NAND U3576 ( .A(n3316), .B(n3315), .Z(n3409) );
  XNOR U3577 ( .A(n3410), .B(n3409), .Z(n3411) );
  NANDN U3578 ( .A(n18487), .B(n3317), .Z(n3319) );
  XOR U3579 ( .A(b[15]), .B(a[23]), .Z(n3472) );
  NANDN U3580 ( .A(n18311), .B(n3472), .Z(n3318) );
  AND U3581 ( .A(n3319), .B(n3318), .Z(n3406) );
  NANDN U3582 ( .A(n18853), .B(n3320), .Z(n3322) );
  XOR U3583 ( .A(b[21]), .B(a[17]), .Z(n3475) );
  NANDN U3584 ( .A(n18926), .B(n3475), .Z(n3321) );
  AND U3585 ( .A(n3322), .B(n3321), .Z(n3404) );
  NANDN U3586 ( .A(n17613), .B(n3323), .Z(n3325) );
  XOR U3587 ( .A(b[9]), .B(a[29]), .Z(n3478) );
  NANDN U3588 ( .A(n17739), .B(n3478), .Z(n3324) );
  NAND U3589 ( .A(n3325), .B(n3324), .Z(n3403) );
  XNOR U3590 ( .A(n3404), .B(n3403), .Z(n3405) );
  XOR U3591 ( .A(n3406), .B(n3405), .Z(n3412) );
  XOR U3592 ( .A(n3411), .B(n3412), .Z(n3418) );
  XOR U3593 ( .A(n3417), .B(n3418), .Z(n3430) );
  XNOR U3594 ( .A(n3429), .B(n3430), .Z(n3361) );
  XNOR U3595 ( .A(n3362), .B(n3361), .Z(n3363) );
  XOR U3596 ( .A(n3364), .B(n3363), .Z(n3482) );
  XNOR U3597 ( .A(n3481), .B(n3482), .Z(n3483) );
  XNOR U3598 ( .A(n3484), .B(n3483), .Z(n3357) );
  XOR U3599 ( .A(n3358), .B(n3357), .Z(n3350) );
  NANDN U3600 ( .A(n3327), .B(n3326), .Z(n3331) );
  NANDN U3601 ( .A(n3329), .B(n3328), .Z(n3330) );
  AND U3602 ( .A(n3331), .B(n3330), .Z(n3349) );
  XNOR U3603 ( .A(n3350), .B(n3349), .Z(n3351) );
  NANDN U3604 ( .A(n3333), .B(n3332), .Z(n3337) );
  NAND U3605 ( .A(n3335), .B(n3334), .Z(n3336) );
  NAND U3606 ( .A(n3337), .B(n3336), .Z(n3352) );
  XNOR U3607 ( .A(n3351), .B(n3352), .Z(n3343) );
  XNOR U3608 ( .A(n3344), .B(n3343), .Z(n3345) );
  XNOR U3609 ( .A(n3346), .B(n3345), .Z(n3487) );
  XNOR U3610 ( .A(sreg[133]), .B(n3487), .Z(n3489) );
  NANDN U3611 ( .A(sreg[132]), .B(n3338), .Z(n3342) );
  NANDN U3612 ( .A(n3340), .B(n3339), .Z(n3341) );
  NAND U3613 ( .A(n3342), .B(n3341), .Z(n3488) );
  XNOR U3614 ( .A(n3489), .B(n3488), .Z(c[133]) );
  NANDN U3615 ( .A(n3344), .B(n3343), .Z(n3348) );
  NANDN U3616 ( .A(n3346), .B(n3345), .Z(n3347) );
  AND U3617 ( .A(n3348), .B(n3347), .Z(n3495) );
  NANDN U3618 ( .A(n3350), .B(n3349), .Z(n3354) );
  NANDN U3619 ( .A(n3352), .B(n3351), .Z(n3353) );
  AND U3620 ( .A(n3354), .B(n3353), .Z(n3493) );
  NANDN U3621 ( .A(n3356), .B(n3355), .Z(n3360) );
  NAND U3622 ( .A(n3358), .B(n3357), .Z(n3359) );
  AND U3623 ( .A(n3360), .B(n3359), .Z(n3500) );
  NANDN U3624 ( .A(n3362), .B(n3361), .Z(n3366) );
  NANDN U3625 ( .A(n3364), .B(n3363), .Z(n3365) );
  AND U3626 ( .A(n3366), .B(n3365), .Z(n3629) );
  NANDN U3627 ( .A(n3368), .B(n3367), .Z(n3372) );
  NAND U3628 ( .A(n3370), .B(n3369), .Z(n3371) );
  AND U3629 ( .A(n3372), .B(n3371), .Z(n3628) );
  XNOR U3630 ( .A(n3629), .B(n3628), .Z(n3631) );
  NANDN U3631 ( .A(n3374), .B(n3373), .Z(n3378) );
  NANDN U3632 ( .A(n3376), .B(n3375), .Z(n3377) );
  AND U3633 ( .A(n3378), .B(n3377), .Z(n3576) );
  NANDN U3634 ( .A(n19237), .B(n3379), .Z(n3381) );
  XOR U3635 ( .A(b[27]), .B(a[12]), .Z(n3522) );
  NANDN U3636 ( .A(n19277), .B(n3522), .Z(n3380) );
  AND U3637 ( .A(n3381), .B(n3380), .Z(n3583) );
  NANDN U3638 ( .A(n17072), .B(n3382), .Z(n3384) );
  XOR U3639 ( .A(b[5]), .B(a[34]), .Z(n3525) );
  NANDN U3640 ( .A(n17223), .B(n3525), .Z(n3383) );
  AND U3641 ( .A(n3384), .B(n3383), .Z(n3581) );
  NANDN U3642 ( .A(n18673), .B(n3385), .Z(n3387) );
  XOR U3643 ( .A(b[19]), .B(a[20]), .Z(n3528) );
  NANDN U3644 ( .A(n18758), .B(n3528), .Z(n3386) );
  NAND U3645 ( .A(n3387), .B(n3386), .Z(n3580) );
  XNOR U3646 ( .A(n3581), .B(n3580), .Z(n3582) );
  XNOR U3647 ( .A(n3583), .B(n3582), .Z(n3574) );
  NANDN U3648 ( .A(n19425), .B(n3388), .Z(n3390) );
  XOR U3649 ( .A(b[31]), .B(a[8]), .Z(n3531) );
  NANDN U3650 ( .A(n19426), .B(n3531), .Z(n3389) );
  AND U3651 ( .A(n3390), .B(n3389), .Z(n3543) );
  NANDN U3652 ( .A(n17067), .B(n3391), .Z(n3393) );
  XOR U3653 ( .A(b[3]), .B(a[36]), .Z(n3534) );
  NANDN U3654 ( .A(n17068), .B(n3534), .Z(n3392) );
  AND U3655 ( .A(n3393), .B(n3392), .Z(n3541) );
  NANDN U3656 ( .A(n18514), .B(n3394), .Z(n3396) );
  XOR U3657 ( .A(b[17]), .B(a[22]), .Z(n3537) );
  NANDN U3658 ( .A(n18585), .B(n3537), .Z(n3395) );
  NAND U3659 ( .A(n3396), .B(n3395), .Z(n3540) );
  XNOR U3660 ( .A(n3541), .B(n3540), .Z(n3542) );
  XOR U3661 ( .A(n3543), .B(n3542), .Z(n3575) );
  XOR U3662 ( .A(n3574), .B(n3575), .Z(n3577) );
  XOR U3663 ( .A(n3576), .B(n3577), .Z(n3511) );
  NANDN U3664 ( .A(n3398), .B(n3397), .Z(n3402) );
  NANDN U3665 ( .A(n3400), .B(n3399), .Z(n3401) );
  AND U3666 ( .A(n3402), .B(n3401), .Z(n3564) );
  NANDN U3667 ( .A(n3404), .B(n3403), .Z(n3408) );
  NANDN U3668 ( .A(n3406), .B(n3405), .Z(n3407) );
  NAND U3669 ( .A(n3408), .B(n3407), .Z(n3565) );
  XNOR U3670 ( .A(n3564), .B(n3565), .Z(n3566) );
  NANDN U3671 ( .A(n3410), .B(n3409), .Z(n3414) );
  NANDN U3672 ( .A(n3412), .B(n3411), .Z(n3413) );
  NAND U3673 ( .A(n3414), .B(n3413), .Z(n3567) );
  XNOR U3674 ( .A(n3566), .B(n3567), .Z(n3510) );
  XNOR U3675 ( .A(n3511), .B(n3510), .Z(n3513) );
  NANDN U3676 ( .A(n3416), .B(n3415), .Z(n3420) );
  NANDN U3677 ( .A(n3418), .B(n3417), .Z(n3419) );
  AND U3678 ( .A(n3420), .B(n3419), .Z(n3512) );
  XOR U3679 ( .A(n3513), .B(n3512), .Z(n3625) );
  NANDN U3680 ( .A(n3422), .B(n3421), .Z(n3426) );
  NANDN U3681 ( .A(n3424), .B(n3423), .Z(n3425) );
  AND U3682 ( .A(n3426), .B(n3425), .Z(n3622) );
  NANDN U3683 ( .A(n3428), .B(n3427), .Z(n3432) );
  NANDN U3684 ( .A(n3430), .B(n3429), .Z(n3431) );
  AND U3685 ( .A(n3432), .B(n3431), .Z(n3507) );
  NANDN U3686 ( .A(n3434), .B(n3433), .Z(n3438) );
  OR U3687 ( .A(n3436), .B(n3435), .Z(n3437) );
  AND U3688 ( .A(n3438), .B(n3437), .Z(n3505) );
  NANDN U3689 ( .A(n3440), .B(n3439), .Z(n3444) );
  NANDN U3690 ( .A(n3442), .B(n3441), .Z(n3443) );
  AND U3691 ( .A(n3444), .B(n3443), .Z(n3571) );
  NANDN U3692 ( .A(n3446), .B(n3445), .Z(n3450) );
  NANDN U3693 ( .A(n3448), .B(n3447), .Z(n3449) );
  NAND U3694 ( .A(n3450), .B(n3449), .Z(n3570) );
  XNOR U3695 ( .A(n3571), .B(n3570), .Z(n3573) );
  NAND U3696 ( .A(b[0]), .B(a[38]), .Z(n3451) );
  XNOR U3697 ( .A(b[1]), .B(n3451), .Z(n3453) );
  NANDN U3698 ( .A(b[0]), .B(a[37]), .Z(n3452) );
  NAND U3699 ( .A(n3453), .B(n3452), .Z(n3519) );
  NANDN U3700 ( .A(n19394), .B(n3454), .Z(n3456) );
  XOR U3701 ( .A(b[29]), .B(a[10]), .Z(n3595) );
  NANDN U3702 ( .A(n19395), .B(n3595), .Z(n3455) );
  AND U3703 ( .A(n3456), .B(n3455), .Z(n3517) );
  AND U3704 ( .A(b[31]), .B(a[6]), .Z(n3516) );
  XNOR U3705 ( .A(n3517), .B(n3516), .Z(n3518) );
  XNOR U3706 ( .A(n3519), .B(n3518), .Z(n3559) );
  NANDN U3707 ( .A(n19005), .B(n3457), .Z(n3459) );
  XOR U3708 ( .A(b[23]), .B(a[16]), .Z(n3598) );
  NANDN U3709 ( .A(n19055), .B(n3598), .Z(n3458) );
  AND U3710 ( .A(n3459), .B(n3458), .Z(n3588) );
  NANDN U3711 ( .A(n17362), .B(n3460), .Z(n3462) );
  XOR U3712 ( .A(b[7]), .B(a[32]), .Z(n3601) );
  NANDN U3713 ( .A(n17522), .B(n3601), .Z(n3461) );
  AND U3714 ( .A(n3462), .B(n3461), .Z(n3587) );
  NANDN U3715 ( .A(n19116), .B(n3463), .Z(n3465) );
  XOR U3716 ( .A(b[25]), .B(a[14]), .Z(n3604) );
  NANDN U3717 ( .A(n19179), .B(n3604), .Z(n3464) );
  NAND U3718 ( .A(n3465), .B(n3464), .Z(n3586) );
  XOR U3719 ( .A(n3587), .B(n3586), .Z(n3589) );
  XOR U3720 ( .A(n3588), .B(n3589), .Z(n3558) );
  XOR U3721 ( .A(n3559), .B(n3558), .Z(n3561) );
  NANDN U3722 ( .A(n18113), .B(n3466), .Z(n3468) );
  XOR U3723 ( .A(b[13]), .B(a[26]), .Z(n3607) );
  NANDN U3724 ( .A(n18229), .B(n3607), .Z(n3467) );
  AND U3725 ( .A(n3468), .B(n3467), .Z(n3553) );
  NANDN U3726 ( .A(n17888), .B(n3469), .Z(n3471) );
  XOR U3727 ( .A(b[11]), .B(a[28]), .Z(n3610) );
  NANDN U3728 ( .A(n18025), .B(n3610), .Z(n3470) );
  NAND U3729 ( .A(n3471), .B(n3470), .Z(n3552) );
  XNOR U3730 ( .A(n3553), .B(n3552), .Z(n3555) );
  NANDN U3731 ( .A(n18487), .B(n3472), .Z(n3474) );
  XOR U3732 ( .A(b[15]), .B(a[24]), .Z(n3613) );
  NANDN U3733 ( .A(n18311), .B(n3613), .Z(n3473) );
  AND U3734 ( .A(n3474), .B(n3473), .Z(n3549) );
  NANDN U3735 ( .A(n18853), .B(n3475), .Z(n3477) );
  XOR U3736 ( .A(b[21]), .B(a[18]), .Z(n3616) );
  NANDN U3737 ( .A(n18926), .B(n3616), .Z(n3476) );
  AND U3738 ( .A(n3477), .B(n3476), .Z(n3547) );
  NANDN U3739 ( .A(n17613), .B(n3478), .Z(n3480) );
  XOR U3740 ( .A(b[9]), .B(a[30]), .Z(n3619) );
  NANDN U3741 ( .A(n17739), .B(n3619), .Z(n3479) );
  NAND U3742 ( .A(n3480), .B(n3479), .Z(n3546) );
  XNOR U3743 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U3744 ( .A(n3549), .B(n3548), .Z(n3554) );
  XOR U3745 ( .A(n3555), .B(n3554), .Z(n3560) );
  XOR U3746 ( .A(n3561), .B(n3560), .Z(n3572) );
  XOR U3747 ( .A(n3573), .B(n3572), .Z(n3504) );
  XNOR U3748 ( .A(n3505), .B(n3504), .Z(n3506) );
  XOR U3749 ( .A(n3507), .B(n3506), .Z(n3623) );
  XNOR U3750 ( .A(n3622), .B(n3623), .Z(n3624) );
  XNOR U3751 ( .A(n3625), .B(n3624), .Z(n3630) );
  XOR U3752 ( .A(n3631), .B(n3630), .Z(n3499) );
  NANDN U3753 ( .A(n3482), .B(n3481), .Z(n3486) );
  NANDN U3754 ( .A(n3484), .B(n3483), .Z(n3485) );
  AND U3755 ( .A(n3486), .B(n3485), .Z(n3498) );
  XOR U3756 ( .A(n3499), .B(n3498), .Z(n3501) );
  XNOR U3757 ( .A(n3500), .B(n3501), .Z(n3492) );
  XNOR U3758 ( .A(n3493), .B(n3492), .Z(n3494) );
  XNOR U3759 ( .A(n3495), .B(n3494), .Z(n3634) );
  XNOR U3760 ( .A(sreg[134]), .B(n3634), .Z(n3636) );
  NANDN U3761 ( .A(sreg[133]), .B(n3487), .Z(n3491) );
  NAND U3762 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND U3763 ( .A(n3491), .B(n3490), .Z(n3635) );
  XNOR U3764 ( .A(n3636), .B(n3635), .Z(c[134]) );
  NANDN U3765 ( .A(n3493), .B(n3492), .Z(n3497) );
  NANDN U3766 ( .A(n3495), .B(n3494), .Z(n3496) );
  AND U3767 ( .A(n3497), .B(n3496), .Z(n3642) );
  NANDN U3768 ( .A(n3499), .B(n3498), .Z(n3503) );
  NANDN U3769 ( .A(n3501), .B(n3500), .Z(n3502) );
  AND U3770 ( .A(n3503), .B(n3502), .Z(n3640) );
  NANDN U3771 ( .A(n3505), .B(n3504), .Z(n3509) );
  NANDN U3772 ( .A(n3507), .B(n3506), .Z(n3508) );
  AND U3773 ( .A(n3509), .B(n3508), .Z(n3778) );
  NANDN U3774 ( .A(n3511), .B(n3510), .Z(n3515) );
  NAND U3775 ( .A(n3513), .B(n3512), .Z(n3514) );
  AND U3776 ( .A(n3515), .B(n3514), .Z(n3777) );
  XNOR U3777 ( .A(n3778), .B(n3777), .Z(n3780) );
  NANDN U3778 ( .A(n3517), .B(n3516), .Z(n3521) );
  NANDN U3779 ( .A(n3519), .B(n3518), .Z(n3520) );
  AND U3780 ( .A(n3521), .B(n3520), .Z(n3713) );
  NANDN U3781 ( .A(n19237), .B(n3522), .Z(n3524) );
  XOR U3782 ( .A(b[27]), .B(a[13]), .Z(n3657) );
  NANDN U3783 ( .A(n19277), .B(n3657), .Z(n3523) );
  AND U3784 ( .A(n3524), .B(n3523), .Z(n3720) );
  NANDN U3785 ( .A(n17072), .B(n3525), .Z(n3527) );
  XOR U3786 ( .A(b[5]), .B(a[35]), .Z(n3660) );
  NANDN U3787 ( .A(n17223), .B(n3660), .Z(n3526) );
  AND U3788 ( .A(n3527), .B(n3526), .Z(n3718) );
  NANDN U3789 ( .A(n18673), .B(n3528), .Z(n3530) );
  XOR U3790 ( .A(b[19]), .B(a[21]), .Z(n3663) );
  NANDN U3791 ( .A(n18758), .B(n3663), .Z(n3529) );
  NAND U3792 ( .A(n3530), .B(n3529), .Z(n3717) );
  XNOR U3793 ( .A(n3718), .B(n3717), .Z(n3719) );
  XNOR U3794 ( .A(n3720), .B(n3719), .Z(n3711) );
  NANDN U3795 ( .A(n19425), .B(n3531), .Z(n3533) );
  XOR U3796 ( .A(b[31]), .B(a[9]), .Z(n3666) );
  NANDN U3797 ( .A(n19426), .B(n3666), .Z(n3532) );
  AND U3798 ( .A(n3533), .B(n3532), .Z(n3678) );
  NANDN U3799 ( .A(n17067), .B(n3534), .Z(n3536) );
  XOR U3800 ( .A(b[3]), .B(a[37]), .Z(n3669) );
  NANDN U3801 ( .A(n17068), .B(n3669), .Z(n3535) );
  AND U3802 ( .A(n3536), .B(n3535), .Z(n3676) );
  NANDN U3803 ( .A(n18514), .B(n3537), .Z(n3539) );
  XOR U3804 ( .A(b[17]), .B(a[23]), .Z(n3672) );
  NANDN U3805 ( .A(n18585), .B(n3672), .Z(n3538) );
  NAND U3806 ( .A(n3539), .B(n3538), .Z(n3675) );
  XNOR U3807 ( .A(n3676), .B(n3675), .Z(n3677) );
  XOR U3808 ( .A(n3678), .B(n3677), .Z(n3712) );
  XOR U3809 ( .A(n3711), .B(n3712), .Z(n3714) );
  XOR U3810 ( .A(n3713), .B(n3714), .Z(n3760) );
  NANDN U3811 ( .A(n3541), .B(n3540), .Z(n3545) );
  NANDN U3812 ( .A(n3543), .B(n3542), .Z(n3544) );
  AND U3813 ( .A(n3545), .B(n3544), .Z(n3699) );
  NANDN U3814 ( .A(n3547), .B(n3546), .Z(n3551) );
  NANDN U3815 ( .A(n3549), .B(n3548), .Z(n3550) );
  NAND U3816 ( .A(n3551), .B(n3550), .Z(n3700) );
  XNOR U3817 ( .A(n3699), .B(n3700), .Z(n3701) );
  NANDN U3818 ( .A(n3553), .B(n3552), .Z(n3557) );
  NAND U3819 ( .A(n3555), .B(n3554), .Z(n3556) );
  NAND U3820 ( .A(n3557), .B(n3556), .Z(n3702) );
  XNOR U3821 ( .A(n3701), .B(n3702), .Z(n3759) );
  XNOR U3822 ( .A(n3760), .B(n3759), .Z(n3762) );
  NAND U3823 ( .A(n3559), .B(n3558), .Z(n3563) );
  NAND U3824 ( .A(n3561), .B(n3560), .Z(n3562) );
  AND U3825 ( .A(n3563), .B(n3562), .Z(n3761) );
  XOR U3826 ( .A(n3762), .B(n3761), .Z(n3774) );
  NANDN U3827 ( .A(n3565), .B(n3564), .Z(n3569) );
  NANDN U3828 ( .A(n3567), .B(n3566), .Z(n3568) );
  AND U3829 ( .A(n3569), .B(n3568), .Z(n3771) );
  NANDN U3830 ( .A(n3575), .B(n3574), .Z(n3579) );
  OR U3831 ( .A(n3577), .B(n3576), .Z(n3578) );
  AND U3832 ( .A(n3579), .B(n3578), .Z(n3766) );
  NANDN U3833 ( .A(n3581), .B(n3580), .Z(n3585) );
  NANDN U3834 ( .A(n3583), .B(n3582), .Z(n3584) );
  AND U3835 ( .A(n3585), .B(n3584), .Z(n3706) );
  NANDN U3836 ( .A(n3587), .B(n3586), .Z(n3591) );
  OR U3837 ( .A(n3589), .B(n3588), .Z(n3590) );
  NAND U3838 ( .A(n3591), .B(n3590), .Z(n3705) );
  XNOR U3839 ( .A(n3706), .B(n3705), .Z(n3707) );
  NAND U3840 ( .A(b[0]), .B(a[39]), .Z(n3592) );
  XNOR U3841 ( .A(b[1]), .B(n3592), .Z(n3594) );
  NANDN U3842 ( .A(b[0]), .B(a[38]), .Z(n3593) );
  NAND U3843 ( .A(n3594), .B(n3593), .Z(n3654) );
  NANDN U3844 ( .A(n19394), .B(n3595), .Z(n3597) );
  XOR U3845 ( .A(b[29]), .B(a[11]), .Z(n3732) );
  NANDN U3846 ( .A(n19395), .B(n3732), .Z(n3596) );
  AND U3847 ( .A(n3597), .B(n3596), .Z(n3652) );
  AND U3848 ( .A(b[31]), .B(a[7]), .Z(n3651) );
  XNOR U3849 ( .A(n3652), .B(n3651), .Z(n3653) );
  XNOR U3850 ( .A(n3654), .B(n3653), .Z(n3693) );
  NANDN U3851 ( .A(n19005), .B(n3598), .Z(n3600) );
  XOR U3852 ( .A(b[23]), .B(a[17]), .Z(n3735) );
  NANDN U3853 ( .A(n19055), .B(n3735), .Z(n3599) );
  AND U3854 ( .A(n3600), .B(n3599), .Z(n3726) );
  NANDN U3855 ( .A(n17362), .B(n3601), .Z(n3603) );
  XOR U3856 ( .A(b[7]), .B(a[33]), .Z(n3738) );
  NANDN U3857 ( .A(n17522), .B(n3738), .Z(n3602) );
  AND U3858 ( .A(n3603), .B(n3602), .Z(n3724) );
  NANDN U3859 ( .A(n19116), .B(n3604), .Z(n3606) );
  XOR U3860 ( .A(b[25]), .B(a[15]), .Z(n3741) );
  NANDN U3861 ( .A(n19179), .B(n3741), .Z(n3605) );
  NAND U3862 ( .A(n3606), .B(n3605), .Z(n3723) );
  XNOR U3863 ( .A(n3724), .B(n3723), .Z(n3725) );
  XOR U3864 ( .A(n3726), .B(n3725), .Z(n3694) );
  XNOR U3865 ( .A(n3693), .B(n3694), .Z(n3695) );
  NANDN U3866 ( .A(n18113), .B(n3607), .Z(n3609) );
  XOR U3867 ( .A(b[13]), .B(a[27]), .Z(n3744) );
  NANDN U3868 ( .A(n18229), .B(n3744), .Z(n3608) );
  AND U3869 ( .A(n3609), .B(n3608), .Z(n3688) );
  NANDN U3870 ( .A(n17888), .B(n3610), .Z(n3612) );
  XOR U3871 ( .A(b[11]), .B(a[29]), .Z(n3747) );
  NANDN U3872 ( .A(n18025), .B(n3747), .Z(n3611) );
  NAND U3873 ( .A(n3612), .B(n3611), .Z(n3687) );
  XNOR U3874 ( .A(n3688), .B(n3687), .Z(n3689) );
  NANDN U3875 ( .A(n18487), .B(n3613), .Z(n3615) );
  XOR U3876 ( .A(b[15]), .B(a[25]), .Z(n3750) );
  NANDN U3877 ( .A(n18311), .B(n3750), .Z(n3614) );
  AND U3878 ( .A(n3615), .B(n3614), .Z(n3684) );
  NANDN U3879 ( .A(n18853), .B(n3616), .Z(n3618) );
  XOR U3880 ( .A(b[21]), .B(a[19]), .Z(n3753) );
  NANDN U3881 ( .A(n18926), .B(n3753), .Z(n3617) );
  AND U3882 ( .A(n3618), .B(n3617), .Z(n3682) );
  NANDN U3883 ( .A(n17613), .B(n3619), .Z(n3621) );
  XOR U3884 ( .A(b[9]), .B(a[31]), .Z(n3756) );
  NANDN U3885 ( .A(n17739), .B(n3756), .Z(n3620) );
  NAND U3886 ( .A(n3621), .B(n3620), .Z(n3681) );
  XNOR U3887 ( .A(n3682), .B(n3681), .Z(n3683) );
  XOR U3888 ( .A(n3684), .B(n3683), .Z(n3690) );
  XOR U3889 ( .A(n3689), .B(n3690), .Z(n3696) );
  XOR U3890 ( .A(n3695), .B(n3696), .Z(n3708) );
  XNOR U3891 ( .A(n3707), .B(n3708), .Z(n3765) );
  XNOR U3892 ( .A(n3766), .B(n3765), .Z(n3767) );
  XOR U3893 ( .A(n3768), .B(n3767), .Z(n3772) );
  XNOR U3894 ( .A(n3771), .B(n3772), .Z(n3773) );
  XNOR U3895 ( .A(n3774), .B(n3773), .Z(n3779) );
  XOR U3896 ( .A(n3780), .B(n3779), .Z(n3646) );
  NANDN U3897 ( .A(n3623), .B(n3622), .Z(n3627) );
  NANDN U3898 ( .A(n3625), .B(n3624), .Z(n3626) );
  AND U3899 ( .A(n3627), .B(n3626), .Z(n3645) );
  XNOR U3900 ( .A(n3646), .B(n3645), .Z(n3647) );
  NANDN U3901 ( .A(n3629), .B(n3628), .Z(n3633) );
  NAND U3902 ( .A(n3631), .B(n3630), .Z(n3632) );
  NAND U3903 ( .A(n3633), .B(n3632), .Z(n3648) );
  XNOR U3904 ( .A(n3647), .B(n3648), .Z(n3639) );
  XNOR U3905 ( .A(n3640), .B(n3639), .Z(n3641) );
  XNOR U3906 ( .A(n3642), .B(n3641), .Z(n3783) );
  XNOR U3907 ( .A(sreg[135]), .B(n3783), .Z(n3785) );
  NANDN U3908 ( .A(sreg[134]), .B(n3634), .Z(n3638) );
  NAND U3909 ( .A(n3636), .B(n3635), .Z(n3637) );
  NAND U3910 ( .A(n3638), .B(n3637), .Z(n3784) );
  XNOR U3911 ( .A(n3785), .B(n3784), .Z(c[135]) );
  NANDN U3912 ( .A(n3640), .B(n3639), .Z(n3644) );
  NANDN U3913 ( .A(n3642), .B(n3641), .Z(n3643) );
  AND U3914 ( .A(n3644), .B(n3643), .Z(n3791) );
  NANDN U3915 ( .A(n3646), .B(n3645), .Z(n3650) );
  NANDN U3916 ( .A(n3648), .B(n3647), .Z(n3649) );
  AND U3917 ( .A(n3650), .B(n3649), .Z(n3789) );
  NANDN U3918 ( .A(n3652), .B(n3651), .Z(n3656) );
  NANDN U3919 ( .A(n3654), .B(n3653), .Z(n3655) );
  AND U3920 ( .A(n3656), .B(n3655), .Z(n3880) );
  NANDN U3921 ( .A(n19237), .B(n3657), .Z(n3659) );
  XOR U3922 ( .A(b[27]), .B(a[14]), .Z(n3824) );
  NANDN U3923 ( .A(n19277), .B(n3824), .Z(n3658) );
  AND U3924 ( .A(n3659), .B(n3658), .Z(n3887) );
  NANDN U3925 ( .A(n17072), .B(n3660), .Z(n3662) );
  XOR U3926 ( .A(b[5]), .B(a[36]), .Z(n3827) );
  NANDN U3927 ( .A(n17223), .B(n3827), .Z(n3661) );
  AND U3928 ( .A(n3662), .B(n3661), .Z(n3885) );
  NANDN U3929 ( .A(n18673), .B(n3663), .Z(n3665) );
  XOR U3930 ( .A(b[19]), .B(a[22]), .Z(n3830) );
  NANDN U3931 ( .A(n18758), .B(n3830), .Z(n3664) );
  NAND U3932 ( .A(n3665), .B(n3664), .Z(n3884) );
  XNOR U3933 ( .A(n3885), .B(n3884), .Z(n3886) );
  XNOR U3934 ( .A(n3887), .B(n3886), .Z(n3878) );
  NANDN U3935 ( .A(n19425), .B(n3666), .Z(n3668) );
  XOR U3936 ( .A(b[31]), .B(a[10]), .Z(n3833) );
  NANDN U3937 ( .A(n19426), .B(n3833), .Z(n3667) );
  AND U3938 ( .A(n3668), .B(n3667), .Z(n3845) );
  NANDN U3939 ( .A(n17067), .B(n3669), .Z(n3671) );
  XOR U3940 ( .A(b[3]), .B(a[38]), .Z(n3836) );
  NANDN U3941 ( .A(n17068), .B(n3836), .Z(n3670) );
  AND U3942 ( .A(n3671), .B(n3670), .Z(n3843) );
  NANDN U3943 ( .A(n18514), .B(n3672), .Z(n3674) );
  XOR U3944 ( .A(b[17]), .B(a[24]), .Z(n3839) );
  NANDN U3945 ( .A(n18585), .B(n3839), .Z(n3673) );
  NAND U3946 ( .A(n3674), .B(n3673), .Z(n3842) );
  XNOR U3947 ( .A(n3843), .B(n3842), .Z(n3844) );
  XOR U3948 ( .A(n3845), .B(n3844), .Z(n3879) );
  XOR U3949 ( .A(n3878), .B(n3879), .Z(n3881) );
  XOR U3950 ( .A(n3880), .B(n3881), .Z(n3813) );
  NANDN U3951 ( .A(n3676), .B(n3675), .Z(n3680) );
  NANDN U3952 ( .A(n3678), .B(n3677), .Z(n3679) );
  AND U3953 ( .A(n3680), .B(n3679), .Z(n3866) );
  NANDN U3954 ( .A(n3682), .B(n3681), .Z(n3686) );
  NANDN U3955 ( .A(n3684), .B(n3683), .Z(n3685) );
  NAND U3956 ( .A(n3686), .B(n3685), .Z(n3867) );
  XNOR U3957 ( .A(n3866), .B(n3867), .Z(n3868) );
  NANDN U3958 ( .A(n3688), .B(n3687), .Z(n3692) );
  NANDN U3959 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U3960 ( .A(n3692), .B(n3691), .Z(n3869) );
  XNOR U3961 ( .A(n3868), .B(n3869), .Z(n3812) );
  XNOR U3962 ( .A(n3813), .B(n3812), .Z(n3815) );
  NANDN U3963 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U3964 ( .A(n3696), .B(n3695), .Z(n3697) );
  AND U3965 ( .A(n3698), .B(n3697), .Z(n3814) );
  XOR U3966 ( .A(n3815), .B(n3814), .Z(n3928) );
  NANDN U3967 ( .A(n3700), .B(n3699), .Z(n3704) );
  NANDN U3968 ( .A(n3702), .B(n3701), .Z(n3703) );
  AND U3969 ( .A(n3704), .B(n3703), .Z(n3926) );
  NANDN U3970 ( .A(n3706), .B(n3705), .Z(n3710) );
  NANDN U3971 ( .A(n3708), .B(n3707), .Z(n3709) );
  AND U3972 ( .A(n3710), .B(n3709), .Z(n3809) );
  NANDN U3973 ( .A(n3712), .B(n3711), .Z(n3716) );
  OR U3974 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U3975 ( .A(n3716), .B(n3715), .Z(n3807) );
  NANDN U3976 ( .A(n3718), .B(n3717), .Z(n3722) );
  NANDN U3977 ( .A(n3720), .B(n3719), .Z(n3721) );
  AND U3978 ( .A(n3722), .B(n3721), .Z(n3873) );
  NANDN U3979 ( .A(n3724), .B(n3723), .Z(n3728) );
  NANDN U3980 ( .A(n3726), .B(n3725), .Z(n3727) );
  NAND U3981 ( .A(n3728), .B(n3727), .Z(n3872) );
  XNOR U3982 ( .A(n3873), .B(n3872), .Z(n3874) );
  NAND U3983 ( .A(b[0]), .B(a[40]), .Z(n3729) );
  XNOR U3984 ( .A(b[1]), .B(n3729), .Z(n3731) );
  NANDN U3985 ( .A(b[0]), .B(a[39]), .Z(n3730) );
  NAND U3986 ( .A(n3731), .B(n3730), .Z(n3821) );
  NANDN U3987 ( .A(n19394), .B(n3732), .Z(n3734) );
  XOR U3988 ( .A(b[29]), .B(a[12]), .Z(n3896) );
  NANDN U3989 ( .A(n19395), .B(n3896), .Z(n3733) );
  AND U3990 ( .A(n3734), .B(n3733), .Z(n3819) );
  AND U3991 ( .A(b[31]), .B(a[8]), .Z(n3818) );
  XNOR U3992 ( .A(n3819), .B(n3818), .Z(n3820) );
  XNOR U3993 ( .A(n3821), .B(n3820), .Z(n3860) );
  NANDN U3994 ( .A(n19005), .B(n3735), .Z(n3737) );
  XOR U3995 ( .A(b[23]), .B(a[18]), .Z(n3902) );
  NANDN U3996 ( .A(n19055), .B(n3902), .Z(n3736) );
  AND U3997 ( .A(n3737), .B(n3736), .Z(n3893) );
  NANDN U3998 ( .A(n17362), .B(n3738), .Z(n3740) );
  XOR U3999 ( .A(b[7]), .B(a[34]), .Z(n3905) );
  NANDN U4000 ( .A(n17522), .B(n3905), .Z(n3739) );
  AND U4001 ( .A(n3740), .B(n3739), .Z(n3891) );
  NANDN U4002 ( .A(n19116), .B(n3741), .Z(n3743) );
  XOR U4003 ( .A(b[25]), .B(a[16]), .Z(n3908) );
  NANDN U4004 ( .A(n19179), .B(n3908), .Z(n3742) );
  NAND U4005 ( .A(n3743), .B(n3742), .Z(n3890) );
  XNOR U4006 ( .A(n3891), .B(n3890), .Z(n3892) );
  XOR U4007 ( .A(n3893), .B(n3892), .Z(n3861) );
  XNOR U4008 ( .A(n3860), .B(n3861), .Z(n3862) );
  NANDN U4009 ( .A(n18113), .B(n3744), .Z(n3746) );
  XOR U4010 ( .A(b[13]), .B(a[28]), .Z(n3911) );
  NANDN U4011 ( .A(n18229), .B(n3911), .Z(n3745) );
  AND U4012 ( .A(n3746), .B(n3745), .Z(n3855) );
  NANDN U4013 ( .A(n17888), .B(n3747), .Z(n3749) );
  XOR U4014 ( .A(b[11]), .B(a[30]), .Z(n3914) );
  NANDN U4015 ( .A(n18025), .B(n3914), .Z(n3748) );
  NAND U4016 ( .A(n3749), .B(n3748), .Z(n3854) );
  XNOR U4017 ( .A(n3855), .B(n3854), .Z(n3856) );
  NANDN U4018 ( .A(n18487), .B(n3750), .Z(n3752) );
  XOR U4019 ( .A(b[15]), .B(a[26]), .Z(n3917) );
  NANDN U4020 ( .A(n18311), .B(n3917), .Z(n3751) );
  AND U4021 ( .A(n3752), .B(n3751), .Z(n3851) );
  NANDN U4022 ( .A(n18853), .B(n3753), .Z(n3755) );
  XOR U4023 ( .A(b[21]), .B(a[20]), .Z(n3920) );
  NANDN U4024 ( .A(n18926), .B(n3920), .Z(n3754) );
  AND U4025 ( .A(n3755), .B(n3754), .Z(n3849) );
  NANDN U4026 ( .A(n17613), .B(n3756), .Z(n3758) );
  XOR U4027 ( .A(b[9]), .B(a[32]), .Z(n3923) );
  NANDN U4028 ( .A(n17739), .B(n3923), .Z(n3757) );
  NAND U4029 ( .A(n3758), .B(n3757), .Z(n3848) );
  XNOR U4030 ( .A(n3849), .B(n3848), .Z(n3850) );
  XOR U4031 ( .A(n3851), .B(n3850), .Z(n3857) );
  XOR U4032 ( .A(n3856), .B(n3857), .Z(n3863) );
  XOR U4033 ( .A(n3862), .B(n3863), .Z(n3875) );
  XNOR U4034 ( .A(n3874), .B(n3875), .Z(n3806) );
  XNOR U4035 ( .A(n3807), .B(n3806), .Z(n3808) );
  XOR U4036 ( .A(n3809), .B(n3808), .Z(n3927) );
  XOR U4037 ( .A(n3926), .B(n3927), .Z(n3929) );
  XOR U4038 ( .A(n3928), .B(n3929), .Z(n3803) );
  NANDN U4039 ( .A(n3760), .B(n3759), .Z(n3764) );
  NAND U4040 ( .A(n3762), .B(n3761), .Z(n3763) );
  AND U4041 ( .A(n3764), .B(n3763), .Z(n3801) );
  NANDN U4042 ( .A(n3766), .B(n3765), .Z(n3770) );
  NANDN U4043 ( .A(n3768), .B(n3767), .Z(n3769) );
  AND U4044 ( .A(n3770), .B(n3769), .Z(n3800) );
  XNOR U4045 ( .A(n3801), .B(n3800), .Z(n3802) );
  XNOR U4046 ( .A(n3803), .B(n3802), .Z(n3794) );
  NANDN U4047 ( .A(n3772), .B(n3771), .Z(n3776) );
  NANDN U4048 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U4049 ( .A(n3776), .B(n3775), .Z(n3795) );
  XNOR U4050 ( .A(n3794), .B(n3795), .Z(n3796) );
  NANDN U4051 ( .A(n3778), .B(n3777), .Z(n3782) );
  NAND U4052 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4053 ( .A(n3782), .B(n3781), .Z(n3797) );
  XNOR U4054 ( .A(n3796), .B(n3797), .Z(n3788) );
  XNOR U4055 ( .A(n3789), .B(n3788), .Z(n3790) );
  XNOR U4056 ( .A(n3791), .B(n3790), .Z(n3932) );
  XNOR U4057 ( .A(sreg[136]), .B(n3932), .Z(n3934) );
  NANDN U4058 ( .A(sreg[135]), .B(n3783), .Z(n3787) );
  NAND U4059 ( .A(n3785), .B(n3784), .Z(n3786) );
  NAND U4060 ( .A(n3787), .B(n3786), .Z(n3933) );
  XNOR U4061 ( .A(n3934), .B(n3933), .Z(c[136]) );
  NANDN U4062 ( .A(n3789), .B(n3788), .Z(n3793) );
  NANDN U4063 ( .A(n3791), .B(n3790), .Z(n3792) );
  AND U4064 ( .A(n3793), .B(n3792), .Z(n3940) );
  NANDN U4065 ( .A(n3795), .B(n3794), .Z(n3799) );
  NANDN U4066 ( .A(n3797), .B(n3796), .Z(n3798) );
  AND U4067 ( .A(n3799), .B(n3798), .Z(n3938) );
  NANDN U4068 ( .A(n3801), .B(n3800), .Z(n3805) );
  NANDN U4069 ( .A(n3803), .B(n3802), .Z(n3804) );
  AND U4070 ( .A(n3805), .B(n3804), .Z(n3946) );
  NANDN U4071 ( .A(n3807), .B(n3806), .Z(n3811) );
  NANDN U4072 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U4073 ( .A(n3811), .B(n3810), .Z(n3950) );
  NANDN U4074 ( .A(n3813), .B(n3812), .Z(n3817) );
  NAND U4075 ( .A(n3815), .B(n3814), .Z(n3816) );
  AND U4076 ( .A(n3817), .B(n3816), .Z(n3949) );
  XNOR U4077 ( .A(n3950), .B(n3949), .Z(n3952) );
  NANDN U4078 ( .A(n3819), .B(n3818), .Z(n3823) );
  NANDN U4079 ( .A(n3821), .B(n3820), .Z(n3822) );
  AND U4080 ( .A(n3823), .B(n3822), .Z(n4029) );
  NANDN U4081 ( .A(n19237), .B(n3824), .Z(n3826) );
  XOR U4082 ( .A(b[27]), .B(a[15]), .Z(n3973) );
  NANDN U4083 ( .A(n19277), .B(n3973), .Z(n3825) );
  AND U4084 ( .A(n3826), .B(n3825), .Z(n4036) );
  NANDN U4085 ( .A(n17072), .B(n3827), .Z(n3829) );
  XOR U4086 ( .A(b[5]), .B(a[37]), .Z(n3976) );
  NANDN U4087 ( .A(n17223), .B(n3976), .Z(n3828) );
  AND U4088 ( .A(n3829), .B(n3828), .Z(n4034) );
  NANDN U4089 ( .A(n18673), .B(n3830), .Z(n3832) );
  XOR U4090 ( .A(b[19]), .B(a[23]), .Z(n3979) );
  NANDN U4091 ( .A(n18758), .B(n3979), .Z(n3831) );
  NAND U4092 ( .A(n3832), .B(n3831), .Z(n4033) );
  XNOR U4093 ( .A(n4034), .B(n4033), .Z(n4035) );
  XNOR U4094 ( .A(n4036), .B(n4035), .Z(n4027) );
  NANDN U4095 ( .A(n19425), .B(n3833), .Z(n3835) );
  XOR U4096 ( .A(b[31]), .B(a[11]), .Z(n3982) );
  NANDN U4097 ( .A(n19426), .B(n3982), .Z(n3834) );
  AND U4098 ( .A(n3835), .B(n3834), .Z(n3994) );
  NANDN U4099 ( .A(n17067), .B(n3836), .Z(n3838) );
  XOR U4100 ( .A(b[3]), .B(a[39]), .Z(n3985) );
  NANDN U4101 ( .A(n17068), .B(n3985), .Z(n3837) );
  AND U4102 ( .A(n3838), .B(n3837), .Z(n3992) );
  NANDN U4103 ( .A(n18514), .B(n3839), .Z(n3841) );
  XOR U4104 ( .A(b[17]), .B(a[25]), .Z(n3988) );
  NANDN U4105 ( .A(n18585), .B(n3988), .Z(n3840) );
  NAND U4106 ( .A(n3841), .B(n3840), .Z(n3991) );
  XNOR U4107 ( .A(n3992), .B(n3991), .Z(n3993) );
  XOR U4108 ( .A(n3994), .B(n3993), .Z(n4028) );
  XOR U4109 ( .A(n4027), .B(n4028), .Z(n4030) );
  XOR U4110 ( .A(n4029), .B(n4030), .Z(n3962) );
  NANDN U4111 ( .A(n3843), .B(n3842), .Z(n3847) );
  NANDN U4112 ( .A(n3845), .B(n3844), .Z(n3846) );
  AND U4113 ( .A(n3847), .B(n3846), .Z(n4015) );
  NANDN U4114 ( .A(n3849), .B(n3848), .Z(n3853) );
  NANDN U4115 ( .A(n3851), .B(n3850), .Z(n3852) );
  NAND U4116 ( .A(n3853), .B(n3852), .Z(n4016) );
  XNOR U4117 ( .A(n4015), .B(n4016), .Z(n4017) );
  NANDN U4118 ( .A(n3855), .B(n3854), .Z(n3859) );
  NANDN U4119 ( .A(n3857), .B(n3856), .Z(n3858) );
  NAND U4120 ( .A(n3859), .B(n3858), .Z(n4018) );
  XNOR U4121 ( .A(n4017), .B(n4018), .Z(n3961) );
  XNOR U4122 ( .A(n3962), .B(n3961), .Z(n3964) );
  NANDN U4123 ( .A(n3861), .B(n3860), .Z(n3865) );
  NANDN U4124 ( .A(n3863), .B(n3862), .Z(n3864) );
  AND U4125 ( .A(n3865), .B(n3864), .Z(n3963) );
  XOR U4126 ( .A(n3964), .B(n3963), .Z(n4078) );
  NANDN U4127 ( .A(n3867), .B(n3866), .Z(n3871) );
  NANDN U4128 ( .A(n3869), .B(n3868), .Z(n3870) );
  AND U4129 ( .A(n3871), .B(n3870), .Z(n4075) );
  NANDN U4130 ( .A(n3873), .B(n3872), .Z(n3877) );
  NANDN U4131 ( .A(n3875), .B(n3874), .Z(n3876) );
  AND U4132 ( .A(n3877), .B(n3876), .Z(n3958) );
  NANDN U4133 ( .A(n3879), .B(n3878), .Z(n3883) );
  OR U4134 ( .A(n3881), .B(n3880), .Z(n3882) );
  AND U4135 ( .A(n3883), .B(n3882), .Z(n3956) );
  NANDN U4136 ( .A(n3885), .B(n3884), .Z(n3889) );
  NANDN U4137 ( .A(n3887), .B(n3886), .Z(n3888) );
  AND U4138 ( .A(n3889), .B(n3888), .Z(n4022) );
  NANDN U4139 ( .A(n3891), .B(n3890), .Z(n3895) );
  NANDN U4140 ( .A(n3893), .B(n3892), .Z(n3894) );
  NAND U4141 ( .A(n3895), .B(n3894), .Z(n4021) );
  XNOR U4142 ( .A(n4022), .B(n4021), .Z(n4023) );
  NANDN U4143 ( .A(n19394), .B(n3896), .Z(n3898) );
  XOR U4144 ( .A(b[29]), .B(a[13]), .Z(n4048) );
  NANDN U4145 ( .A(n19395), .B(n4048), .Z(n3897) );
  AND U4146 ( .A(n3898), .B(n3897), .Z(n3968) );
  AND U4147 ( .A(b[31]), .B(a[9]), .Z(n3967) );
  XNOR U4148 ( .A(n3968), .B(n3967), .Z(n3969) );
  NAND U4149 ( .A(b[0]), .B(a[41]), .Z(n3899) );
  XNOR U4150 ( .A(b[1]), .B(n3899), .Z(n3901) );
  NANDN U4151 ( .A(b[0]), .B(a[40]), .Z(n3900) );
  NAND U4152 ( .A(n3901), .B(n3900), .Z(n3970) );
  XNOR U4153 ( .A(n3969), .B(n3970), .Z(n4009) );
  NANDN U4154 ( .A(n19005), .B(n3902), .Z(n3904) );
  XOR U4155 ( .A(b[23]), .B(a[19]), .Z(n4051) );
  NANDN U4156 ( .A(n19055), .B(n4051), .Z(n3903) );
  AND U4157 ( .A(n3904), .B(n3903), .Z(n4042) );
  NANDN U4158 ( .A(n17362), .B(n3905), .Z(n3907) );
  XOR U4159 ( .A(b[7]), .B(a[35]), .Z(n4054) );
  NANDN U4160 ( .A(n17522), .B(n4054), .Z(n3906) );
  AND U4161 ( .A(n3907), .B(n3906), .Z(n4040) );
  NANDN U4162 ( .A(n19116), .B(n3908), .Z(n3910) );
  XOR U4163 ( .A(b[25]), .B(a[17]), .Z(n4057) );
  NANDN U4164 ( .A(n19179), .B(n4057), .Z(n3909) );
  NAND U4165 ( .A(n3910), .B(n3909), .Z(n4039) );
  XNOR U4166 ( .A(n4040), .B(n4039), .Z(n4041) );
  XOR U4167 ( .A(n4042), .B(n4041), .Z(n4010) );
  XNOR U4168 ( .A(n4009), .B(n4010), .Z(n4011) );
  NANDN U4169 ( .A(n18113), .B(n3911), .Z(n3913) );
  XOR U4170 ( .A(b[13]), .B(a[29]), .Z(n4060) );
  NANDN U4171 ( .A(n18229), .B(n4060), .Z(n3912) );
  AND U4172 ( .A(n3913), .B(n3912), .Z(n4004) );
  NANDN U4173 ( .A(n17888), .B(n3914), .Z(n3916) );
  XOR U4174 ( .A(b[11]), .B(a[31]), .Z(n4063) );
  NANDN U4175 ( .A(n18025), .B(n4063), .Z(n3915) );
  NAND U4176 ( .A(n3916), .B(n3915), .Z(n4003) );
  XNOR U4177 ( .A(n4004), .B(n4003), .Z(n4005) );
  NANDN U4178 ( .A(n18487), .B(n3917), .Z(n3919) );
  XOR U4179 ( .A(b[15]), .B(a[27]), .Z(n4066) );
  NANDN U4180 ( .A(n18311), .B(n4066), .Z(n3918) );
  AND U4181 ( .A(n3919), .B(n3918), .Z(n4000) );
  NANDN U4182 ( .A(n18853), .B(n3920), .Z(n3922) );
  XOR U4183 ( .A(b[21]), .B(a[21]), .Z(n4069) );
  NANDN U4184 ( .A(n18926), .B(n4069), .Z(n3921) );
  AND U4185 ( .A(n3922), .B(n3921), .Z(n3998) );
  NANDN U4186 ( .A(n17613), .B(n3923), .Z(n3925) );
  XOR U4187 ( .A(b[9]), .B(a[33]), .Z(n4072) );
  NANDN U4188 ( .A(n17739), .B(n4072), .Z(n3924) );
  NAND U4189 ( .A(n3925), .B(n3924), .Z(n3997) );
  XNOR U4190 ( .A(n3998), .B(n3997), .Z(n3999) );
  XOR U4191 ( .A(n4000), .B(n3999), .Z(n4006) );
  XOR U4192 ( .A(n4005), .B(n4006), .Z(n4012) );
  XOR U4193 ( .A(n4011), .B(n4012), .Z(n4024) );
  XNOR U4194 ( .A(n4023), .B(n4024), .Z(n3955) );
  XNOR U4195 ( .A(n3956), .B(n3955), .Z(n3957) );
  XOR U4196 ( .A(n3958), .B(n3957), .Z(n4076) );
  XNOR U4197 ( .A(n4075), .B(n4076), .Z(n4077) );
  XNOR U4198 ( .A(n4078), .B(n4077), .Z(n3951) );
  XOR U4199 ( .A(n3952), .B(n3951), .Z(n3944) );
  NANDN U4200 ( .A(n3927), .B(n3926), .Z(n3931) );
  OR U4201 ( .A(n3929), .B(n3928), .Z(n3930) );
  AND U4202 ( .A(n3931), .B(n3930), .Z(n3943) );
  XNOR U4203 ( .A(n3944), .B(n3943), .Z(n3945) );
  XNOR U4204 ( .A(n3946), .B(n3945), .Z(n3937) );
  XNOR U4205 ( .A(n3938), .B(n3937), .Z(n3939) );
  XNOR U4206 ( .A(n3940), .B(n3939), .Z(n4081) );
  XNOR U4207 ( .A(sreg[137]), .B(n4081), .Z(n4083) );
  NANDN U4208 ( .A(sreg[136]), .B(n3932), .Z(n3936) );
  NAND U4209 ( .A(n3934), .B(n3933), .Z(n3935) );
  NAND U4210 ( .A(n3936), .B(n3935), .Z(n4082) );
  XNOR U4211 ( .A(n4083), .B(n4082), .Z(c[137]) );
  NANDN U4212 ( .A(n3938), .B(n3937), .Z(n3942) );
  NANDN U4213 ( .A(n3940), .B(n3939), .Z(n3941) );
  AND U4214 ( .A(n3942), .B(n3941), .Z(n4089) );
  NANDN U4215 ( .A(n3944), .B(n3943), .Z(n3948) );
  NANDN U4216 ( .A(n3946), .B(n3945), .Z(n3947) );
  AND U4217 ( .A(n3948), .B(n3947), .Z(n4087) );
  NANDN U4218 ( .A(n3950), .B(n3949), .Z(n3954) );
  NAND U4219 ( .A(n3952), .B(n3951), .Z(n3953) );
  AND U4220 ( .A(n3954), .B(n3953), .Z(n4094) );
  NANDN U4221 ( .A(n3956), .B(n3955), .Z(n3960) );
  NANDN U4222 ( .A(n3958), .B(n3957), .Z(n3959) );
  AND U4223 ( .A(n3960), .B(n3959), .Z(n4099) );
  NANDN U4224 ( .A(n3962), .B(n3961), .Z(n3966) );
  NAND U4225 ( .A(n3964), .B(n3963), .Z(n3965) );
  AND U4226 ( .A(n3966), .B(n3965), .Z(n4098) );
  XNOR U4227 ( .A(n4099), .B(n4098), .Z(n4101) );
  NANDN U4228 ( .A(n3968), .B(n3967), .Z(n3972) );
  NANDN U4229 ( .A(n3970), .B(n3969), .Z(n3971) );
  AND U4230 ( .A(n3972), .B(n3971), .Z(n4178) );
  NANDN U4231 ( .A(n19237), .B(n3973), .Z(n3975) );
  XOR U4232 ( .A(b[27]), .B(a[16]), .Z(n4122) );
  NANDN U4233 ( .A(n19277), .B(n4122), .Z(n3974) );
  AND U4234 ( .A(n3975), .B(n3974), .Z(n4185) );
  NANDN U4235 ( .A(n17072), .B(n3976), .Z(n3978) );
  XOR U4236 ( .A(b[5]), .B(a[38]), .Z(n4125) );
  NANDN U4237 ( .A(n17223), .B(n4125), .Z(n3977) );
  AND U4238 ( .A(n3978), .B(n3977), .Z(n4183) );
  NANDN U4239 ( .A(n18673), .B(n3979), .Z(n3981) );
  XOR U4240 ( .A(b[19]), .B(a[24]), .Z(n4128) );
  NANDN U4241 ( .A(n18758), .B(n4128), .Z(n3980) );
  NAND U4242 ( .A(n3981), .B(n3980), .Z(n4182) );
  XNOR U4243 ( .A(n4183), .B(n4182), .Z(n4184) );
  XNOR U4244 ( .A(n4185), .B(n4184), .Z(n4176) );
  NANDN U4245 ( .A(n19425), .B(n3982), .Z(n3984) );
  XOR U4246 ( .A(b[31]), .B(a[12]), .Z(n4131) );
  NANDN U4247 ( .A(n19426), .B(n4131), .Z(n3983) );
  AND U4248 ( .A(n3984), .B(n3983), .Z(n4143) );
  NANDN U4249 ( .A(n17067), .B(n3985), .Z(n3987) );
  XOR U4250 ( .A(b[3]), .B(a[40]), .Z(n4134) );
  NANDN U4251 ( .A(n17068), .B(n4134), .Z(n3986) );
  AND U4252 ( .A(n3987), .B(n3986), .Z(n4141) );
  NANDN U4253 ( .A(n18514), .B(n3988), .Z(n3990) );
  XOR U4254 ( .A(b[17]), .B(a[26]), .Z(n4137) );
  NANDN U4255 ( .A(n18585), .B(n4137), .Z(n3989) );
  NAND U4256 ( .A(n3990), .B(n3989), .Z(n4140) );
  XNOR U4257 ( .A(n4141), .B(n4140), .Z(n4142) );
  XOR U4258 ( .A(n4143), .B(n4142), .Z(n4177) );
  XOR U4259 ( .A(n4176), .B(n4177), .Z(n4179) );
  XOR U4260 ( .A(n4178), .B(n4179), .Z(n4111) );
  NANDN U4261 ( .A(n3992), .B(n3991), .Z(n3996) );
  NANDN U4262 ( .A(n3994), .B(n3993), .Z(n3995) );
  AND U4263 ( .A(n3996), .B(n3995), .Z(n4164) );
  NANDN U4264 ( .A(n3998), .B(n3997), .Z(n4002) );
  NANDN U4265 ( .A(n4000), .B(n3999), .Z(n4001) );
  NAND U4266 ( .A(n4002), .B(n4001), .Z(n4165) );
  XNOR U4267 ( .A(n4164), .B(n4165), .Z(n4166) );
  NANDN U4268 ( .A(n4004), .B(n4003), .Z(n4008) );
  NANDN U4269 ( .A(n4006), .B(n4005), .Z(n4007) );
  NAND U4270 ( .A(n4008), .B(n4007), .Z(n4167) );
  XNOR U4271 ( .A(n4166), .B(n4167), .Z(n4110) );
  XNOR U4272 ( .A(n4111), .B(n4110), .Z(n4113) );
  NANDN U4273 ( .A(n4010), .B(n4009), .Z(n4014) );
  NANDN U4274 ( .A(n4012), .B(n4011), .Z(n4013) );
  AND U4275 ( .A(n4014), .B(n4013), .Z(n4112) );
  XOR U4276 ( .A(n4113), .B(n4112), .Z(n4227) );
  NANDN U4277 ( .A(n4016), .B(n4015), .Z(n4020) );
  NANDN U4278 ( .A(n4018), .B(n4017), .Z(n4019) );
  AND U4279 ( .A(n4020), .B(n4019), .Z(n4224) );
  NANDN U4280 ( .A(n4022), .B(n4021), .Z(n4026) );
  NANDN U4281 ( .A(n4024), .B(n4023), .Z(n4025) );
  AND U4282 ( .A(n4026), .B(n4025), .Z(n4107) );
  NANDN U4283 ( .A(n4028), .B(n4027), .Z(n4032) );
  OR U4284 ( .A(n4030), .B(n4029), .Z(n4031) );
  AND U4285 ( .A(n4032), .B(n4031), .Z(n4105) );
  NANDN U4286 ( .A(n4034), .B(n4033), .Z(n4038) );
  NANDN U4287 ( .A(n4036), .B(n4035), .Z(n4037) );
  AND U4288 ( .A(n4038), .B(n4037), .Z(n4171) );
  NANDN U4289 ( .A(n4040), .B(n4039), .Z(n4044) );
  NANDN U4290 ( .A(n4042), .B(n4041), .Z(n4043) );
  NAND U4291 ( .A(n4044), .B(n4043), .Z(n4170) );
  XNOR U4292 ( .A(n4171), .B(n4170), .Z(n4172) );
  NAND U4293 ( .A(b[0]), .B(a[42]), .Z(n4045) );
  XNOR U4294 ( .A(b[1]), .B(n4045), .Z(n4047) );
  NANDN U4295 ( .A(b[0]), .B(a[41]), .Z(n4046) );
  NAND U4296 ( .A(n4047), .B(n4046), .Z(n4119) );
  NANDN U4297 ( .A(n19394), .B(n4048), .Z(n4050) );
  XOR U4298 ( .A(b[29]), .B(a[14]), .Z(n4197) );
  NANDN U4299 ( .A(n19395), .B(n4197), .Z(n4049) );
  AND U4300 ( .A(n4050), .B(n4049), .Z(n4117) );
  AND U4301 ( .A(b[31]), .B(a[10]), .Z(n4116) );
  XNOR U4302 ( .A(n4117), .B(n4116), .Z(n4118) );
  XNOR U4303 ( .A(n4119), .B(n4118), .Z(n4158) );
  NANDN U4304 ( .A(n19005), .B(n4051), .Z(n4053) );
  XOR U4305 ( .A(b[23]), .B(a[20]), .Z(n4200) );
  NANDN U4306 ( .A(n19055), .B(n4200), .Z(n4052) );
  AND U4307 ( .A(n4053), .B(n4052), .Z(n4191) );
  NANDN U4308 ( .A(n17362), .B(n4054), .Z(n4056) );
  XOR U4309 ( .A(b[7]), .B(a[36]), .Z(n4203) );
  NANDN U4310 ( .A(n17522), .B(n4203), .Z(n4055) );
  AND U4311 ( .A(n4056), .B(n4055), .Z(n4189) );
  NANDN U4312 ( .A(n19116), .B(n4057), .Z(n4059) );
  XOR U4313 ( .A(b[25]), .B(a[18]), .Z(n4206) );
  NANDN U4314 ( .A(n19179), .B(n4206), .Z(n4058) );
  NAND U4315 ( .A(n4059), .B(n4058), .Z(n4188) );
  XNOR U4316 ( .A(n4189), .B(n4188), .Z(n4190) );
  XOR U4317 ( .A(n4191), .B(n4190), .Z(n4159) );
  XNOR U4318 ( .A(n4158), .B(n4159), .Z(n4160) );
  NANDN U4319 ( .A(n18113), .B(n4060), .Z(n4062) );
  XOR U4320 ( .A(b[13]), .B(a[30]), .Z(n4209) );
  NANDN U4321 ( .A(n18229), .B(n4209), .Z(n4061) );
  AND U4322 ( .A(n4062), .B(n4061), .Z(n4153) );
  NANDN U4323 ( .A(n17888), .B(n4063), .Z(n4065) );
  XOR U4324 ( .A(b[11]), .B(a[32]), .Z(n4212) );
  NANDN U4325 ( .A(n18025), .B(n4212), .Z(n4064) );
  NAND U4326 ( .A(n4065), .B(n4064), .Z(n4152) );
  XNOR U4327 ( .A(n4153), .B(n4152), .Z(n4154) );
  NANDN U4328 ( .A(n18487), .B(n4066), .Z(n4068) );
  XOR U4329 ( .A(b[15]), .B(a[28]), .Z(n4215) );
  NANDN U4330 ( .A(n18311), .B(n4215), .Z(n4067) );
  AND U4331 ( .A(n4068), .B(n4067), .Z(n4149) );
  NANDN U4332 ( .A(n18853), .B(n4069), .Z(n4071) );
  XOR U4333 ( .A(b[21]), .B(a[22]), .Z(n4218) );
  NANDN U4334 ( .A(n18926), .B(n4218), .Z(n4070) );
  AND U4335 ( .A(n4071), .B(n4070), .Z(n4147) );
  NANDN U4336 ( .A(n17613), .B(n4072), .Z(n4074) );
  XOR U4337 ( .A(b[9]), .B(a[34]), .Z(n4221) );
  NANDN U4338 ( .A(n17739), .B(n4221), .Z(n4073) );
  NAND U4339 ( .A(n4074), .B(n4073), .Z(n4146) );
  XNOR U4340 ( .A(n4147), .B(n4146), .Z(n4148) );
  XOR U4341 ( .A(n4149), .B(n4148), .Z(n4155) );
  XOR U4342 ( .A(n4154), .B(n4155), .Z(n4161) );
  XOR U4343 ( .A(n4160), .B(n4161), .Z(n4173) );
  XNOR U4344 ( .A(n4172), .B(n4173), .Z(n4104) );
  XNOR U4345 ( .A(n4105), .B(n4104), .Z(n4106) );
  XOR U4346 ( .A(n4107), .B(n4106), .Z(n4225) );
  XNOR U4347 ( .A(n4224), .B(n4225), .Z(n4226) );
  XNOR U4348 ( .A(n4227), .B(n4226), .Z(n4100) );
  XOR U4349 ( .A(n4101), .B(n4100), .Z(n4093) );
  NANDN U4350 ( .A(n4076), .B(n4075), .Z(n4080) );
  NANDN U4351 ( .A(n4078), .B(n4077), .Z(n4079) );
  AND U4352 ( .A(n4080), .B(n4079), .Z(n4092) );
  XOR U4353 ( .A(n4093), .B(n4092), .Z(n4095) );
  XNOR U4354 ( .A(n4094), .B(n4095), .Z(n4086) );
  XNOR U4355 ( .A(n4087), .B(n4086), .Z(n4088) );
  XNOR U4356 ( .A(n4089), .B(n4088), .Z(n4230) );
  XNOR U4357 ( .A(sreg[138]), .B(n4230), .Z(n4232) );
  NANDN U4358 ( .A(sreg[137]), .B(n4081), .Z(n4085) );
  NAND U4359 ( .A(n4083), .B(n4082), .Z(n4084) );
  NAND U4360 ( .A(n4085), .B(n4084), .Z(n4231) );
  XNOR U4361 ( .A(n4232), .B(n4231), .Z(c[138]) );
  NANDN U4362 ( .A(n4087), .B(n4086), .Z(n4091) );
  NANDN U4363 ( .A(n4089), .B(n4088), .Z(n4090) );
  AND U4364 ( .A(n4091), .B(n4090), .Z(n4238) );
  NANDN U4365 ( .A(n4093), .B(n4092), .Z(n4097) );
  NANDN U4366 ( .A(n4095), .B(n4094), .Z(n4096) );
  AND U4367 ( .A(n4097), .B(n4096), .Z(n4236) );
  NANDN U4368 ( .A(n4099), .B(n4098), .Z(n4103) );
  NAND U4369 ( .A(n4101), .B(n4100), .Z(n4102) );
  AND U4370 ( .A(n4103), .B(n4102), .Z(n4243) );
  NANDN U4371 ( .A(n4105), .B(n4104), .Z(n4109) );
  NANDN U4372 ( .A(n4107), .B(n4106), .Z(n4108) );
  AND U4373 ( .A(n4109), .B(n4108), .Z(n4372) );
  NANDN U4374 ( .A(n4111), .B(n4110), .Z(n4115) );
  NAND U4375 ( .A(n4113), .B(n4112), .Z(n4114) );
  AND U4376 ( .A(n4115), .B(n4114), .Z(n4371) );
  XNOR U4377 ( .A(n4372), .B(n4371), .Z(n4374) );
  NANDN U4378 ( .A(n4117), .B(n4116), .Z(n4121) );
  NANDN U4379 ( .A(n4119), .B(n4118), .Z(n4120) );
  AND U4380 ( .A(n4121), .B(n4120), .Z(n4319) );
  NANDN U4381 ( .A(n19237), .B(n4122), .Z(n4124) );
  XOR U4382 ( .A(b[27]), .B(a[17]), .Z(n4265) );
  NANDN U4383 ( .A(n19277), .B(n4265), .Z(n4123) );
  AND U4384 ( .A(n4124), .B(n4123), .Z(n4326) );
  NANDN U4385 ( .A(n17072), .B(n4125), .Z(n4127) );
  XOR U4386 ( .A(b[5]), .B(a[39]), .Z(n4268) );
  NANDN U4387 ( .A(n17223), .B(n4268), .Z(n4126) );
  AND U4388 ( .A(n4127), .B(n4126), .Z(n4324) );
  NANDN U4389 ( .A(n18673), .B(n4128), .Z(n4130) );
  XOR U4390 ( .A(b[19]), .B(a[25]), .Z(n4271) );
  NANDN U4391 ( .A(n18758), .B(n4271), .Z(n4129) );
  NAND U4392 ( .A(n4130), .B(n4129), .Z(n4323) );
  XNOR U4393 ( .A(n4324), .B(n4323), .Z(n4325) );
  XNOR U4394 ( .A(n4326), .B(n4325), .Z(n4317) );
  NANDN U4395 ( .A(n19425), .B(n4131), .Z(n4133) );
  XOR U4396 ( .A(b[31]), .B(a[13]), .Z(n4274) );
  NANDN U4397 ( .A(n19426), .B(n4274), .Z(n4132) );
  AND U4398 ( .A(n4133), .B(n4132), .Z(n4286) );
  NANDN U4399 ( .A(n17067), .B(n4134), .Z(n4136) );
  XOR U4400 ( .A(b[3]), .B(a[41]), .Z(n4277) );
  NANDN U4401 ( .A(n17068), .B(n4277), .Z(n4135) );
  AND U4402 ( .A(n4136), .B(n4135), .Z(n4284) );
  NANDN U4403 ( .A(n18514), .B(n4137), .Z(n4139) );
  XOR U4404 ( .A(b[17]), .B(a[27]), .Z(n4280) );
  NANDN U4405 ( .A(n18585), .B(n4280), .Z(n4138) );
  NAND U4406 ( .A(n4139), .B(n4138), .Z(n4283) );
  XNOR U4407 ( .A(n4284), .B(n4283), .Z(n4285) );
  XOR U4408 ( .A(n4286), .B(n4285), .Z(n4318) );
  XOR U4409 ( .A(n4317), .B(n4318), .Z(n4320) );
  XOR U4410 ( .A(n4319), .B(n4320), .Z(n4254) );
  NANDN U4411 ( .A(n4141), .B(n4140), .Z(n4145) );
  NANDN U4412 ( .A(n4143), .B(n4142), .Z(n4144) );
  AND U4413 ( .A(n4145), .B(n4144), .Z(n4307) );
  NANDN U4414 ( .A(n4147), .B(n4146), .Z(n4151) );
  NANDN U4415 ( .A(n4149), .B(n4148), .Z(n4150) );
  NAND U4416 ( .A(n4151), .B(n4150), .Z(n4308) );
  XNOR U4417 ( .A(n4307), .B(n4308), .Z(n4309) );
  NANDN U4418 ( .A(n4153), .B(n4152), .Z(n4157) );
  NANDN U4419 ( .A(n4155), .B(n4154), .Z(n4156) );
  NAND U4420 ( .A(n4157), .B(n4156), .Z(n4310) );
  XNOR U4421 ( .A(n4309), .B(n4310), .Z(n4253) );
  XNOR U4422 ( .A(n4254), .B(n4253), .Z(n4256) );
  NANDN U4423 ( .A(n4159), .B(n4158), .Z(n4163) );
  NANDN U4424 ( .A(n4161), .B(n4160), .Z(n4162) );
  AND U4425 ( .A(n4163), .B(n4162), .Z(n4255) );
  XOR U4426 ( .A(n4256), .B(n4255), .Z(n4368) );
  NANDN U4427 ( .A(n4165), .B(n4164), .Z(n4169) );
  NANDN U4428 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U4429 ( .A(n4169), .B(n4168), .Z(n4365) );
  NANDN U4430 ( .A(n4171), .B(n4170), .Z(n4175) );
  NANDN U4431 ( .A(n4173), .B(n4172), .Z(n4174) );
  AND U4432 ( .A(n4175), .B(n4174), .Z(n4250) );
  NANDN U4433 ( .A(n4177), .B(n4176), .Z(n4181) );
  OR U4434 ( .A(n4179), .B(n4178), .Z(n4180) );
  AND U4435 ( .A(n4181), .B(n4180), .Z(n4248) );
  NANDN U4436 ( .A(n4183), .B(n4182), .Z(n4187) );
  NANDN U4437 ( .A(n4185), .B(n4184), .Z(n4186) );
  AND U4438 ( .A(n4187), .B(n4186), .Z(n4314) );
  NANDN U4439 ( .A(n4189), .B(n4188), .Z(n4193) );
  NANDN U4440 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND U4441 ( .A(n4193), .B(n4192), .Z(n4313) );
  XNOR U4442 ( .A(n4314), .B(n4313), .Z(n4316) );
  NAND U4443 ( .A(b[0]), .B(a[43]), .Z(n4194) );
  XNOR U4444 ( .A(b[1]), .B(n4194), .Z(n4196) );
  NANDN U4445 ( .A(b[0]), .B(a[42]), .Z(n4195) );
  NAND U4446 ( .A(n4196), .B(n4195), .Z(n4262) );
  NANDN U4447 ( .A(n19394), .B(n4197), .Z(n4199) );
  XOR U4448 ( .A(b[29]), .B(a[15]), .Z(n4338) );
  NANDN U4449 ( .A(n19395), .B(n4338), .Z(n4198) );
  AND U4450 ( .A(n4199), .B(n4198), .Z(n4260) );
  AND U4451 ( .A(b[31]), .B(a[11]), .Z(n4259) );
  XNOR U4452 ( .A(n4260), .B(n4259), .Z(n4261) );
  XNOR U4453 ( .A(n4262), .B(n4261), .Z(n4302) );
  NANDN U4454 ( .A(n19005), .B(n4200), .Z(n4202) );
  XOR U4455 ( .A(b[23]), .B(a[21]), .Z(n4341) );
  NANDN U4456 ( .A(n19055), .B(n4341), .Z(n4201) );
  AND U4457 ( .A(n4202), .B(n4201), .Z(n4331) );
  NANDN U4458 ( .A(n17362), .B(n4203), .Z(n4205) );
  XOR U4459 ( .A(b[7]), .B(a[37]), .Z(n4344) );
  NANDN U4460 ( .A(n17522), .B(n4344), .Z(n4204) );
  AND U4461 ( .A(n4205), .B(n4204), .Z(n4330) );
  NANDN U4462 ( .A(n19116), .B(n4206), .Z(n4208) );
  XOR U4463 ( .A(b[25]), .B(a[19]), .Z(n4347) );
  NANDN U4464 ( .A(n19179), .B(n4347), .Z(n4207) );
  NAND U4465 ( .A(n4208), .B(n4207), .Z(n4329) );
  XOR U4466 ( .A(n4330), .B(n4329), .Z(n4332) );
  XOR U4467 ( .A(n4331), .B(n4332), .Z(n4301) );
  XOR U4468 ( .A(n4302), .B(n4301), .Z(n4304) );
  NANDN U4469 ( .A(n18113), .B(n4209), .Z(n4211) );
  XOR U4470 ( .A(b[13]), .B(a[31]), .Z(n4350) );
  NANDN U4471 ( .A(n18229), .B(n4350), .Z(n4210) );
  AND U4472 ( .A(n4211), .B(n4210), .Z(n4296) );
  NANDN U4473 ( .A(n17888), .B(n4212), .Z(n4214) );
  XOR U4474 ( .A(b[11]), .B(a[33]), .Z(n4353) );
  NANDN U4475 ( .A(n18025), .B(n4353), .Z(n4213) );
  NAND U4476 ( .A(n4214), .B(n4213), .Z(n4295) );
  XNOR U4477 ( .A(n4296), .B(n4295), .Z(n4298) );
  NANDN U4478 ( .A(n18487), .B(n4215), .Z(n4217) );
  XOR U4479 ( .A(b[15]), .B(a[29]), .Z(n4356) );
  NANDN U4480 ( .A(n18311), .B(n4356), .Z(n4216) );
  AND U4481 ( .A(n4217), .B(n4216), .Z(n4292) );
  NANDN U4482 ( .A(n18853), .B(n4218), .Z(n4220) );
  XOR U4483 ( .A(b[21]), .B(a[23]), .Z(n4359) );
  NANDN U4484 ( .A(n18926), .B(n4359), .Z(n4219) );
  AND U4485 ( .A(n4220), .B(n4219), .Z(n4290) );
  NANDN U4486 ( .A(n17613), .B(n4221), .Z(n4223) );
  XOR U4487 ( .A(b[9]), .B(a[35]), .Z(n4362) );
  NANDN U4488 ( .A(n17739), .B(n4362), .Z(n4222) );
  NAND U4489 ( .A(n4223), .B(n4222), .Z(n4289) );
  XNOR U4490 ( .A(n4290), .B(n4289), .Z(n4291) );
  XNOR U4491 ( .A(n4292), .B(n4291), .Z(n4297) );
  XOR U4492 ( .A(n4298), .B(n4297), .Z(n4303) );
  XOR U4493 ( .A(n4304), .B(n4303), .Z(n4315) );
  XOR U4494 ( .A(n4316), .B(n4315), .Z(n4247) );
  XNOR U4495 ( .A(n4248), .B(n4247), .Z(n4249) );
  XOR U4496 ( .A(n4250), .B(n4249), .Z(n4366) );
  XNOR U4497 ( .A(n4365), .B(n4366), .Z(n4367) );
  XNOR U4498 ( .A(n4368), .B(n4367), .Z(n4373) );
  XOR U4499 ( .A(n4374), .B(n4373), .Z(n4242) );
  NANDN U4500 ( .A(n4225), .B(n4224), .Z(n4229) );
  NANDN U4501 ( .A(n4227), .B(n4226), .Z(n4228) );
  AND U4502 ( .A(n4229), .B(n4228), .Z(n4241) );
  XOR U4503 ( .A(n4242), .B(n4241), .Z(n4244) );
  XNOR U4504 ( .A(n4243), .B(n4244), .Z(n4235) );
  XNOR U4505 ( .A(n4236), .B(n4235), .Z(n4237) );
  XNOR U4506 ( .A(n4238), .B(n4237), .Z(n4377) );
  XNOR U4507 ( .A(sreg[139]), .B(n4377), .Z(n4379) );
  NANDN U4508 ( .A(sreg[138]), .B(n4230), .Z(n4234) );
  NAND U4509 ( .A(n4232), .B(n4231), .Z(n4233) );
  NAND U4510 ( .A(n4234), .B(n4233), .Z(n4378) );
  XNOR U4511 ( .A(n4379), .B(n4378), .Z(c[139]) );
  NANDN U4512 ( .A(n4236), .B(n4235), .Z(n4240) );
  NANDN U4513 ( .A(n4238), .B(n4237), .Z(n4239) );
  AND U4514 ( .A(n4240), .B(n4239), .Z(n4385) );
  NANDN U4515 ( .A(n4242), .B(n4241), .Z(n4246) );
  NANDN U4516 ( .A(n4244), .B(n4243), .Z(n4245) );
  AND U4517 ( .A(n4246), .B(n4245), .Z(n4383) );
  NANDN U4518 ( .A(n4248), .B(n4247), .Z(n4252) );
  NANDN U4519 ( .A(n4250), .B(n4249), .Z(n4251) );
  AND U4520 ( .A(n4252), .B(n4251), .Z(n4395) );
  NANDN U4521 ( .A(n4254), .B(n4253), .Z(n4258) );
  NAND U4522 ( .A(n4256), .B(n4255), .Z(n4257) );
  AND U4523 ( .A(n4258), .B(n4257), .Z(n4394) );
  XNOR U4524 ( .A(n4395), .B(n4394), .Z(n4397) );
  NANDN U4525 ( .A(n4260), .B(n4259), .Z(n4264) );
  NANDN U4526 ( .A(n4262), .B(n4261), .Z(n4263) );
  AND U4527 ( .A(n4264), .B(n4263), .Z(n4462) );
  NANDN U4528 ( .A(n19237), .B(n4265), .Z(n4267) );
  XOR U4529 ( .A(b[27]), .B(a[18]), .Z(n4406) );
  NANDN U4530 ( .A(n19277), .B(n4406), .Z(n4266) );
  AND U4531 ( .A(n4267), .B(n4266), .Z(n4469) );
  NANDN U4532 ( .A(n17072), .B(n4268), .Z(n4270) );
  XOR U4533 ( .A(b[5]), .B(a[40]), .Z(n4409) );
  NANDN U4534 ( .A(n17223), .B(n4409), .Z(n4269) );
  AND U4535 ( .A(n4270), .B(n4269), .Z(n4467) );
  NANDN U4536 ( .A(n18673), .B(n4271), .Z(n4273) );
  XOR U4537 ( .A(b[19]), .B(a[26]), .Z(n4412) );
  NANDN U4538 ( .A(n18758), .B(n4412), .Z(n4272) );
  NAND U4539 ( .A(n4273), .B(n4272), .Z(n4466) );
  XNOR U4540 ( .A(n4467), .B(n4466), .Z(n4468) );
  XNOR U4541 ( .A(n4469), .B(n4468), .Z(n4460) );
  NANDN U4542 ( .A(n19425), .B(n4274), .Z(n4276) );
  XOR U4543 ( .A(b[31]), .B(a[14]), .Z(n4415) );
  NANDN U4544 ( .A(n19426), .B(n4415), .Z(n4275) );
  AND U4545 ( .A(n4276), .B(n4275), .Z(n4427) );
  NANDN U4546 ( .A(n17067), .B(n4277), .Z(n4279) );
  XOR U4547 ( .A(b[3]), .B(a[42]), .Z(n4418) );
  NANDN U4548 ( .A(n17068), .B(n4418), .Z(n4278) );
  AND U4549 ( .A(n4279), .B(n4278), .Z(n4425) );
  NANDN U4550 ( .A(n18514), .B(n4280), .Z(n4282) );
  XOR U4551 ( .A(b[17]), .B(a[28]), .Z(n4421) );
  NANDN U4552 ( .A(n18585), .B(n4421), .Z(n4281) );
  NAND U4553 ( .A(n4282), .B(n4281), .Z(n4424) );
  XNOR U4554 ( .A(n4425), .B(n4424), .Z(n4426) );
  XOR U4555 ( .A(n4427), .B(n4426), .Z(n4461) );
  XOR U4556 ( .A(n4460), .B(n4461), .Z(n4463) );
  XOR U4557 ( .A(n4462), .B(n4463), .Z(n4509) );
  NANDN U4558 ( .A(n4284), .B(n4283), .Z(n4288) );
  NANDN U4559 ( .A(n4286), .B(n4285), .Z(n4287) );
  AND U4560 ( .A(n4288), .B(n4287), .Z(n4448) );
  NANDN U4561 ( .A(n4290), .B(n4289), .Z(n4294) );
  NANDN U4562 ( .A(n4292), .B(n4291), .Z(n4293) );
  NAND U4563 ( .A(n4294), .B(n4293), .Z(n4449) );
  XNOR U4564 ( .A(n4448), .B(n4449), .Z(n4450) );
  NANDN U4565 ( .A(n4296), .B(n4295), .Z(n4300) );
  NAND U4566 ( .A(n4298), .B(n4297), .Z(n4299) );
  NAND U4567 ( .A(n4300), .B(n4299), .Z(n4451) );
  XNOR U4568 ( .A(n4450), .B(n4451), .Z(n4508) );
  XNOR U4569 ( .A(n4509), .B(n4508), .Z(n4511) );
  NAND U4570 ( .A(n4302), .B(n4301), .Z(n4306) );
  NAND U4571 ( .A(n4304), .B(n4303), .Z(n4305) );
  AND U4572 ( .A(n4306), .B(n4305), .Z(n4510) );
  XOR U4573 ( .A(n4511), .B(n4510), .Z(n4523) );
  NANDN U4574 ( .A(n4308), .B(n4307), .Z(n4312) );
  NANDN U4575 ( .A(n4310), .B(n4309), .Z(n4311) );
  AND U4576 ( .A(n4312), .B(n4311), .Z(n4520) );
  NANDN U4577 ( .A(n4318), .B(n4317), .Z(n4322) );
  OR U4578 ( .A(n4320), .B(n4319), .Z(n4321) );
  AND U4579 ( .A(n4322), .B(n4321), .Z(n4515) );
  NANDN U4580 ( .A(n4324), .B(n4323), .Z(n4328) );
  NANDN U4581 ( .A(n4326), .B(n4325), .Z(n4327) );
  AND U4582 ( .A(n4328), .B(n4327), .Z(n4455) );
  NANDN U4583 ( .A(n4330), .B(n4329), .Z(n4334) );
  OR U4584 ( .A(n4332), .B(n4331), .Z(n4333) );
  NAND U4585 ( .A(n4334), .B(n4333), .Z(n4454) );
  XNOR U4586 ( .A(n4455), .B(n4454), .Z(n4456) );
  NAND U4587 ( .A(b[0]), .B(a[44]), .Z(n4335) );
  XNOR U4588 ( .A(b[1]), .B(n4335), .Z(n4337) );
  NANDN U4589 ( .A(b[0]), .B(a[43]), .Z(n4336) );
  NAND U4590 ( .A(n4337), .B(n4336), .Z(n4403) );
  NANDN U4591 ( .A(n19394), .B(n4338), .Z(n4340) );
  XOR U4592 ( .A(b[29]), .B(a[16]), .Z(n4478) );
  NANDN U4593 ( .A(n19395), .B(n4478), .Z(n4339) );
  AND U4594 ( .A(n4340), .B(n4339), .Z(n4401) );
  AND U4595 ( .A(b[31]), .B(a[12]), .Z(n4400) );
  XNOR U4596 ( .A(n4401), .B(n4400), .Z(n4402) );
  XNOR U4597 ( .A(n4403), .B(n4402), .Z(n4442) );
  NANDN U4598 ( .A(n19005), .B(n4341), .Z(n4343) );
  XOR U4599 ( .A(b[23]), .B(a[22]), .Z(n4484) );
  NANDN U4600 ( .A(n19055), .B(n4484), .Z(n4342) );
  AND U4601 ( .A(n4343), .B(n4342), .Z(n4475) );
  NANDN U4602 ( .A(n17362), .B(n4344), .Z(n4346) );
  XOR U4603 ( .A(b[7]), .B(a[38]), .Z(n4487) );
  NANDN U4604 ( .A(n17522), .B(n4487), .Z(n4345) );
  AND U4605 ( .A(n4346), .B(n4345), .Z(n4473) );
  NANDN U4606 ( .A(n19116), .B(n4347), .Z(n4349) );
  XOR U4607 ( .A(b[25]), .B(a[20]), .Z(n4490) );
  NANDN U4608 ( .A(n19179), .B(n4490), .Z(n4348) );
  NAND U4609 ( .A(n4349), .B(n4348), .Z(n4472) );
  XNOR U4610 ( .A(n4473), .B(n4472), .Z(n4474) );
  XOR U4611 ( .A(n4475), .B(n4474), .Z(n4443) );
  XNOR U4612 ( .A(n4442), .B(n4443), .Z(n4444) );
  NANDN U4613 ( .A(n18113), .B(n4350), .Z(n4352) );
  XOR U4614 ( .A(b[13]), .B(a[32]), .Z(n4493) );
  NANDN U4615 ( .A(n18229), .B(n4493), .Z(n4351) );
  AND U4616 ( .A(n4352), .B(n4351), .Z(n4437) );
  NANDN U4617 ( .A(n17888), .B(n4353), .Z(n4355) );
  XOR U4618 ( .A(b[11]), .B(a[34]), .Z(n4496) );
  NANDN U4619 ( .A(n18025), .B(n4496), .Z(n4354) );
  NAND U4620 ( .A(n4355), .B(n4354), .Z(n4436) );
  XNOR U4621 ( .A(n4437), .B(n4436), .Z(n4438) );
  NANDN U4622 ( .A(n18487), .B(n4356), .Z(n4358) );
  XOR U4623 ( .A(b[15]), .B(a[30]), .Z(n4499) );
  NANDN U4624 ( .A(n18311), .B(n4499), .Z(n4357) );
  AND U4625 ( .A(n4358), .B(n4357), .Z(n4433) );
  NANDN U4626 ( .A(n18853), .B(n4359), .Z(n4361) );
  XOR U4627 ( .A(b[21]), .B(a[24]), .Z(n4502) );
  NANDN U4628 ( .A(n18926), .B(n4502), .Z(n4360) );
  AND U4629 ( .A(n4361), .B(n4360), .Z(n4431) );
  NANDN U4630 ( .A(n17613), .B(n4362), .Z(n4364) );
  XOR U4631 ( .A(b[9]), .B(a[36]), .Z(n4505) );
  NANDN U4632 ( .A(n17739), .B(n4505), .Z(n4363) );
  NAND U4633 ( .A(n4364), .B(n4363), .Z(n4430) );
  XNOR U4634 ( .A(n4431), .B(n4430), .Z(n4432) );
  XOR U4635 ( .A(n4433), .B(n4432), .Z(n4439) );
  XOR U4636 ( .A(n4438), .B(n4439), .Z(n4445) );
  XOR U4637 ( .A(n4444), .B(n4445), .Z(n4457) );
  XNOR U4638 ( .A(n4456), .B(n4457), .Z(n4514) );
  XNOR U4639 ( .A(n4515), .B(n4514), .Z(n4516) );
  XOR U4640 ( .A(n4517), .B(n4516), .Z(n4521) );
  XNOR U4641 ( .A(n4520), .B(n4521), .Z(n4522) );
  XNOR U4642 ( .A(n4523), .B(n4522), .Z(n4396) );
  XOR U4643 ( .A(n4397), .B(n4396), .Z(n4389) );
  NANDN U4644 ( .A(n4366), .B(n4365), .Z(n4370) );
  NANDN U4645 ( .A(n4368), .B(n4367), .Z(n4369) );
  AND U4646 ( .A(n4370), .B(n4369), .Z(n4388) );
  XNOR U4647 ( .A(n4389), .B(n4388), .Z(n4390) );
  NANDN U4648 ( .A(n4372), .B(n4371), .Z(n4376) );
  NAND U4649 ( .A(n4374), .B(n4373), .Z(n4375) );
  NAND U4650 ( .A(n4376), .B(n4375), .Z(n4391) );
  XNOR U4651 ( .A(n4390), .B(n4391), .Z(n4382) );
  XNOR U4652 ( .A(n4383), .B(n4382), .Z(n4384) );
  XNOR U4653 ( .A(n4385), .B(n4384), .Z(n4526) );
  XNOR U4654 ( .A(sreg[140]), .B(n4526), .Z(n4528) );
  NANDN U4655 ( .A(sreg[139]), .B(n4377), .Z(n4381) );
  NAND U4656 ( .A(n4379), .B(n4378), .Z(n4380) );
  NAND U4657 ( .A(n4381), .B(n4380), .Z(n4527) );
  XNOR U4658 ( .A(n4528), .B(n4527), .Z(c[140]) );
  NANDN U4659 ( .A(n4383), .B(n4382), .Z(n4387) );
  NANDN U4660 ( .A(n4385), .B(n4384), .Z(n4386) );
  AND U4661 ( .A(n4387), .B(n4386), .Z(n4534) );
  NANDN U4662 ( .A(n4389), .B(n4388), .Z(n4393) );
  NANDN U4663 ( .A(n4391), .B(n4390), .Z(n4392) );
  AND U4664 ( .A(n4393), .B(n4392), .Z(n4532) );
  NANDN U4665 ( .A(n4395), .B(n4394), .Z(n4399) );
  NAND U4666 ( .A(n4397), .B(n4396), .Z(n4398) );
  AND U4667 ( .A(n4399), .B(n4398), .Z(n4539) );
  NANDN U4668 ( .A(n4401), .B(n4400), .Z(n4405) );
  NANDN U4669 ( .A(n4403), .B(n4402), .Z(n4404) );
  AND U4670 ( .A(n4405), .B(n4404), .Z(n4623) );
  NANDN U4671 ( .A(n19237), .B(n4406), .Z(n4408) );
  XOR U4672 ( .A(b[27]), .B(a[19]), .Z(n4567) );
  NANDN U4673 ( .A(n19277), .B(n4567), .Z(n4407) );
  AND U4674 ( .A(n4408), .B(n4407), .Z(n4630) );
  NANDN U4675 ( .A(n17072), .B(n4409), .Z(n4411) );
  XOR U4676 ( .A(b[5]), .B(a[41]), .Z(n4570) );
  NANDN U4677 ( .A(n17223), .B(n4570), .Z(n4410) );
  AND U4678 ( .A(n4411), .B(n4410), .Z(n4628) );
  NANDN U4679 ( .A(n18673), .B(n4412), .Z(n4414) );
  XOR U4680 ( .A(b[19]), .B(a[27]), .Z(n4573) );
  NANDN U4681 ( .A(n18758), .B(n4573), .Z(n4413) );
  NAND U4682 ( .A(n4414), .B(n4413), .Z(n4627) );
  XNOR U4683 ( .A(n4628), .B(n4627), .Z(n4629) );
  XNOR U4684 ( .A(n4630), .B(n4629), .Z(n4621) );
  NANDN U4685 ( .A(n19425), .B(n4415), .Z(n4417) );
  XOR U4686 ( .A(b[31]), .B(a[15]), .Z(n4576) );
  NANDN U4687 ( .A(n19426), .B(n4576), .Z(n4416) );
  AND U4688 ( .A(n4417), .B(n4416), .Z(n4588) );
  NANDN U4689 ( .A(n17067), .B(n4418), .Z(n4420) );
  XOR U4690 ( .A(b[3]), .B(a[43]), .Z(n4579) );
  NANDN U4691 ( .A(n17068), .B(n4579), .Z(n4419) );
  AND U4692 ( .A(n4420), .B(n4419), .Z(n4586) );
  NANDN U4693 ( .A(n18514), .B(n4421), .Z(n4423) );
  XOR U4694 ( .A(b[17]), .B(a[29]), .Z(n4582) );
  NANDN U4695 ( .A(n18585), .B(n4582), .Z(n4422) );
  NAND U4696 ( .A(n4423), .B(n4422), .Z(n4585) );
  XNOR U4697 ( .A(n4586), .B(n4585), .Z(n4587) );
  XOR U4698 ( .A(n4588), .B(n4587), .Z(n4622) );
  XOR U4699 ( .A(n4621), .B(n4622), .Z(n4624) );
  XOR U4700 ( .A(n4623), .B(n4624), .Z(n4556) );
  NANDN U4701 ( .A(n4425), .B(n4424), .Z(n4429) );
  NANDN U4702 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U4703 ( .A(n4429), .B(n4428), .Z(n4609) );
  NANDN U4704 ( .A(n4431), .B(n4430), .Z(n4435) );
  NANDN U4705 ( .A(n4433), .B(n4432), .Z(n4434) );
  NAND U4706 ( .A(n4435), .B(n4434), .Z(n4610) );
  XNOR U4707 ( .A(n4609), .B(n4610), .Z(n4611) );
  NANDN U4708 ( .A(n4437), .B(n4436), .Z(n4441) );
  NANDN U4709 ( .A(n4439), .B(n4438), .Z(n4440) );
  NAND U4710 ( .A(n4441), .B(n4440), .Z(n4612) );
  XNOR U4711 ( .A(n4611), .B(n4612), .Z(n4555) );
  XNOR U4712 ( .A(n4556), .B(n4555), .Z(n4558) );
  NANDN U4713 ( .A(n4443), .B(n4442), .Z(n4447) );
  NANDN U4714 ( .A(n4445), .B(n4444), .Z(n4446) );
  AND U4715 ( .A(n4447), .B(n4446), .Z(n4557) );
  XOR U4716 ( .A(n4558), .B(n4557), .Z(n4671) );
  NANDN U4717 ( .A(n4449), .B(n4448), .Z(n4453) );
  NANDN U4718 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U4719 ( .A(n4453), .B(n4452), .Z(n4669) );
  NANDN U4720 ( .A(n4455), .B(n4454), .Z(n4459) );
  NANDN U4721 ( .A(n4457), .B(n4456), .Z(n4458) );
  AND U4722 ( .A(n4459), .B(n4458), .Z(n4552) );
  NANDN U4723 ( .A(n4461), .B(n4460), .Z(n4465) );
  OR U4724 ( .A(n4463), .B(n4462), .Z(n4464) );
  AND U4725 ( .A(n4465), .B(n4464), .Z(n4550) );
  NANDN U4726 ( .A(n4467), .B(n4466), .Z(n4471) );
  NANDN U4727 ( .A(n4469), .B(n4468), .Z(n4470) );
  AND U4728 ( .A(n4471), .B(n4470), .Z(n4616) );
  NANDN U4729 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U4730 ( .A(n4475), .B(n4474), .Z(n4476) );
  NAND U4731 ( .A(n4477), .B(n4476), .Z(n4615) );
  XNOR U4732 ( .A(n4616), .B(n4615), .Z(n4617) );
  NANDN U4733 ( .A(n19394), .B(n4478), .Z(n4480) );
  XOR U4734 ( .A(b[29]), .B(a[17]), .Z(n4642) );
  NANDN U4735 ( .A(n19395), .B(n4642), .Z(n4479) );
  AND U4736 ( .A(n4480), .B(n4479), .Z(n4562) );
  AND U4737 ( .A(b[31]), .B(a[13]), .Z(n4561) );
  XNOR U4738 ( .A(n4562), .B(n4561), .Z(n4563) );
  NAND U4739 ( .A(b[0]), .B(a[45]), .Z(n4481) );
  XNOR U4740 ( .A(b[1]), .B(n4481), .Z(n4483) );
  NANDN U4741 ( .A(b[0]), .B(a[44]), .Z(n4482) );
  NAND U4742 ( .A(n4483), .B(n4482), .Z(n4564) );
  XNOR U4743 ( .A(n4563), .B(n4564), .Z(n4603) );
  NANDN U4744 ( .A(n19005), .B(n4484), .Z(n4486) );
  XOR U4745 ( .A(b[23]), .B(a[23]), .Z(n4645) );
  NANDN U4746 ( .A(n19055), .B(n4645), .Z(n4485) );
  AND U4747 ( .A(n4486), .B(n4485), .Z(n4636) );
  NANDN U4748 ( .A(n17362), .B(n4487), .Z(n4489) );
  XOR U4749 ( .A(b[7]), .B(a[39]), .Z(n4648) );
  NANDN U4750 ( .A(n17522), .B(n4648), .Z(n4488) );
  AND U4751 ( .A(n4489), .B(n4488), .Z(n4634) );
  NANDN U4752 ( .A(n19116), .B(n4490), .Z(n4492) );
  XOR U4753 ( .A(b[25]), .B(a[21]), .Z(n4651) );
  NANDN U4754 ( .A(n19179), .B(n4651), .Z(n4491) );
  NAND U4755 ( .A(n4492), .B(n4491), .Z(n4633) );
  XNOR U4756 ( .A(n4634), .B(n4633), .Z(n4635) );
  XOR U4757 ( .A(n4636), .B(n4635), .Z(n4604) );
  XNOR U4758 ( .A(n4603), .B(n4604), .Z(n4605) );
  NANDN U4759 ( .A(n18113), .B(n4493), .Z(n4495) );
  XOR U4760 ( .A(b[13]), .B(a[33]), .Z(n4654) );
  NANDN U4761 ( .A(n18229), .B(n4654), .Z(n4494) );
  AND U4762 ( .A(n4495), .B(n4494), .Z(n4598) );
  NANDN U4763 ( .A(n17888), .B(n4496), .Z(n4498) );
  XOR U4764 ( .A(b[11]), .B(a[35]), .Z(n4657) );
  NANDN U4765 ( .A(n18025), .B(n4657), .Z(n4497) );
  NAND U4766 ( .A(n4498), .B(n4497), .Z(n4597) );
  XNOR U4767 ( .A(n4598), .B(n4597), .Z(n4599) );
  NANDN U4768 ( .A(n18487), .B(n4499), .Z(n4501) );
  XOR U4769 ( .A(b[15]), .B(a[31]), .Z(n4660) );
  NANDN U4770 ( .A(n18311), .B(n4660), .Z(n4500) );
  AND U4771 ( .A(n4501), .B(n4500), .Z(n4594) );
  NANDN U4772 ( .A(n18853), .B(n4502), .Z(n4504) );
  XOR U4773 ( .A(b[21]), .B(a[25]), .Z(n4663) );
  NANDN U4774 ( .A(n18926), .B(n4663), .Z(n4503) );
  AND U4775 ( .A(n4504), .B(n4503), .Z(n4592) );
  NANDN U4776 ( .A(n17613), .B(n4505), .Z(n4507) );
  XOR U4777 ( .A(b[9]), .B(a[37]), .Z(n4666) );
  NANDN U4778 ( .A(n17739), .B(n4666), .Z(n4506) );
  NAND U4779 ( .A(n4507), .B(n4506), .Z(n4591) );
  XNOR U4780 ( .A(n4592), .B(n4591), .Z(n4593) );
  XOR U4781 ( .A(n4594), .B(n4593), .Z(n4600) );
  XOR U4782 ( .A(n4599), .B(n4600), .Z(n4606) );
  XOR U4783 ( .A(n4605), .B(n4606), .Z(n4618) );
  XNOR U4784 ( .A(n4617), .B(n4618), .Z(n4549) );
  XNOR U4785 ( .A(n4550), .B(n4549), .Z(n4551) );
  XOR U4786 ( .A(n4552), .B(n4551), .Z(n4670) );
  XOR U4787 ( .A(n4669), .B(n4670), .Z(n4672) );
  XOR U4788 ( .A(n4671), .B(n4672), .Z(n4546) );
  NANDN U4789 ( .A(n4509), .B(n4508), .Z(n4513) );
  NAND U4790 ( .A(n4511), .B(n4510), .Z(n4512) );
  AND U4791 ( .A(n4513), .B(n4512), .Z(n4544) );
  NANDN U4792 ( .A(n4515), .B(n4514), .Z(n4519) );
  NANDN U4793 ( .A(n4517), .B(n4516), .Z(n4518) );
  AND U4794 ( .A(n4519), .B(n4518), .Z(n4543) );
  XNOR U4795 ( .A(n4544), .B(n4543), .Z(n4545) );
  XNOR U4796 ( .A(n4546), .B(n4545), .Z(n4537) );
  NANDN U4797 ( .A(n4521), .B(n4520), .Z(n4525) );
  NANDN U4798 ( .A(n4523), .B(n4522), .Z(n4524) );
  NAND U4799 ( .A(n4525), .B(n4524), .Z(n4538) );
  XOR U4800 ( .A(n4537), .B(n4538), .Z(n4540) );
  XNOR U4801 ( .A(n4539), .B(n4540), .Z(n4531) );
  XNOR U4802 ( .A(n4532), .B(n4531), .Z(n4533) );
  XNOR U4803 ( .A(n4534), .B(n4533), .Z(n4675) );
  XNOR U4804 ( .A(sreg[141]), .B(n4675), .Z(n4677) );
  NANDN U4805 ( .A(sreg[140]), .B(n4526), .Z(n4530) );
  NAND U4806 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U4807 ( .A(n4530), .B(n4529), .Z(n4676) );
  XNOR U4808 ( .A(n4677), .B(n4676), .Z(c[141]) );
  NANDN U4809 ( .A(n4532), .B(n4531), .Z(n4536) );
  NANDN U4810 ( .A(n4534), .B(n4533), .Z(n4535) );
  AND U4811 ( .A(n4536), .B(n4535), .Z(n4683) );
  NANDN U4812 ( .A(n4538), .B(n4537), .Z(n4542) );
  NANDN U4813 ( .A(n4540), .B(n4539), .Z(n4541) );
  AND U4814 ( .A(n4542), .B(n4541), .Z(n4681) );
  NANDN U4815 ( .A(n4544), .B(n4543), .Z(n4548) );
  NANDN U4816 ( .A(n4546), .B(n4545), .Z(n4547) );
  AND U4817 ( .A(n4548), .B(n4547), .Z(n4689) );
  NANDN U4818 ( .A(n4550), .B(n4549), .Z(n4554) );
  NANDN U4819 ( .A(n4552), .B(n4551), .Z(n4553) );
  AND U4820 ( .A(n4554), .B(n4553), .Z(n4819) );
  NANDN U4821 ( .A(n4556), .B(n4555), .Z(n4560) );
  NAND U4822 ( .A(n4558), .B(n4557), .Z(n4559) );
  AND U4823 ( .A(n4560), .B(n4559), .Z(n4818) );
  XNOR U4824 ( .A(n4819), .B(n4818), .Z(n4821) );
  NANDN U4825 ( .A(n4562), .B(n4561), .Z(n4566) );
  NANDN U4826 ( .A(n4564), .B(n4563), .Z(n4565) );
  AND U4827 ( .A(n4566), .B(n4565), .Z(n4766) );
  NANDN U4828 ( .A(n19237), .B(n4567), .Z(n4569) );
  XOR U4829 ( .A(b[27]), .B(a[20]), .Z(n4710) );
  NANDN U4830 ( .A(n19277), .B(n4710), .Z(n4568) );
  AND U4831 ( .A(n4569), .B(n4568), .Z(n4773) );
  NANDN U4832 ( .A(n17072), .B(n4570), .Z(n4572) );
  XOR U4833 ( .A(b[5]), .B(a[42]), .Z(n4713) );
  NANDN U4834 ( .A(n17223), .B(n4713), .Z(n4571) );
  AND U4835 ( .A(n4572), .B(n4571), .Z(n4771) );
  NANDN U4836 ( .A(n18673), .B(n4573), .Z(n4575) );
  XOR U4837 ( .A(b[19]), .B(a[28]), .Z(n4716) );
  NANDN U4838 ( .A(n18758), .B(n4716), .Z(n4574) );
  NAND U4839 ( .A(n4575), .B(n4574), .Z(n4770) );
  XNOR U4840 ( .A(n4771), .B(n4770), .Z(n4772) );
  XNOR U4841 ( .A(n4773), .B(n4772), .Z(n4764) );
  NANDN U4842 ( .A(n19425), .B(n4576), .Z(n4578) );
  XOR U4843 ( .A(b[31]), .B(a[16]), .Z(n4719) );
  NANDN U4844 ( .A(n19426), .B(n4719), .Z(n4577) );
  AND U4845 ( .A(n4578), .B(n4577), .Z(n4731) );
  NANDN U4846 ( .A(n17067), .B(n4579), .Z(n4581) );
  XOR U4847 ( .A(b[3]), .B(a[44]), .Z(n4722) );
  NANDN U4848 ( .A(n17068), .B(n4722), .Z(n4580) );
  AND U4849 ( .A(n4581), .B(n4580), .Z(n4729) );
  NANDN U4850 ( .A(n18514), .B(n4582), .Z(n4584) );
  XOR U4851 ( .A(b[17]), .B(a[30]), .Z(n4725) );
  NANDN U4852 ( .A(n18585), .B(n4725), .Z(n4583) );
  NAND U4853 ( .A(n4584), .B(n4583), .Z(n4728) );
  XNOR U4854 ( .A(n4729), .B(n4728), .Z(n4730) );
  XOR U4855 ( .A(n4731), .B(n4730), .Z(n4765) );
  XOR U4856 ( .A(n4764), .B(n4765), .Z(n4767) );
  XOR U4857 ( .A(n4766), .B(n4767), .Z(n4699) );
  NANDN U4858 ( .A(n4586), .B(n4585), .Z(n4590) );
  NANDN U4859 ( .A(n4588), .B(n4587), .Z(n4589) );
  AND U4860 ( .A(n4590), .B(n4589), .Z(n4752) );
  NANDN U4861 ( .A(n4592), .B(n4591), .Z(n4596) );
  NANDN U4862 ( .A(n4594), .B(n4593), .Z(n4595) );
  NAND U4863 ( .A(n4596), .B(n4595), .Z(n4753) );
  XNOR U4864 ( .A(n4752), .B(n4753), .Z(n4754) );
  NANDN U4865 ( .A(n4598), .B(n4597), .Z(n4602) );
  NANDN U4866 ( .A(n4600), .B(n4599), .Z(n4601) );
  NAND U4867 ( .A(n4602), .B(n4601), .Z(n4755) );
  XNOR U4868 ( .A(n4754), .B(n4755), .Z(n4698) );
  XNOR U4869 ( .A(n4699), .B(n4698), .Z(n4701) );
  NANDN U4870 ( .A(n4604), .B(n4603), .Z(n4608) );
  NANDN U4871 ( .A(n4606), .B(n4605), .Z(n4607) );
  AND U4872 ( .A(n4608), .B(n4607), .Z(n4700) );
  XOR U4873 ( .A(n4701), .B(n4700), .Z(n4815) );
  NANDN U4874 ( .A(n4610), .B(n4609), .Z(n4614) );
  NANDN U4875 ( .A(n4612), .B(n4611), .Z(n4613) );
  AND U4876 ( .A(n4614), .B(n4613), .Z(n4812) );
  NANDN U4877 ( .A(n4616), .B(n4615), .Z(n4620) );
  NANDN U4878 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U4879 ( .A(n4620), .B(n4619), .Z(n4695) );
  NANDN U4880 ( .A(n4622), .B(n4621), .Z(n4626) );
  OR U4881 ( .A(n4624), .B(n4623), .Z(n4625) );
  AND U4882 ( .A(n4626), .B(n4625), .Z(n4693) );
  NANDN U4883 ( .A(n4628), .B(n4627), .Z(n4632) );
  NANDN U4884 ( .A(n4630), .B(n4629), .Z(n4631) );
  AND U4885 ( .A(n4632), .B(n4631), .Z(n4759) );
  NANDN U4886 ( .A(n4634), .B(n4633), .Z(n4638) );
  NANDN U4887 ( .A(n4636), .B(n4635), .Z(n4637) );
  NAND U4888 ( .A(n4638), .B(n4637), .Z(n4758) );
  XNOR U4889 ( .A(n4759), .B(n4758), .Z(n4760) );
  NAND U4890 ( .A(b[0]), .B(a[46]), .Z(n4639) );
  XNOR U4891 ( .A(b[1]), .B(n4639), .Z(n4641) );
  NANDN U4892 ( .A(b[0]), .B(a[45]), .Z(n4640) );
  NAND U4893 ( .A(n4641), .B(n4640), .Z(n4707) );
  NANDN U4894 ( .A(n19394), .B(n4642), .Z(n4644) );
  XOR U4895 ( .A(b[29]), .B(a[18]), .Z(n4785) );
  NANDN U4896 ( .A(n19395), .B(n4785), .Z(n4643) );
  AND U4897 ( .A(n4644), .B(n4643), .Z(n4705) );
  AND U4898 ( .A(b[31]), .B(a[14]), .Z(n4704) );
  XNOR U4899 ( .A(n4705), .B(n4704), .Z(n4706) );
  XNOR U4900 ( .A(n4707), .B(n4706), .Z(n4746) );
  NANDN U4901 ( .A(n19005), .B(n4645), .Z(n4647) );
  XOR U4902 ( .A(b[23]), .B(a[24]), .Z(n4788) );
  NANDN U4903 ( .A(n19055), .B(n4788), .Z(n4646) );
  AND U4904 ( .A(n4647), .B(n4646), .Z(n4779) );
  NANDN U4905 ( .A(n17362), .B(n4648), .Z(n4650) );
  XOR U4906 ( .A(b[7]), .B(a[40]), .Z(n4791) );
  NANDN U4907 ( .A(n17522), .B(n4791), .Z(n4649) );
  AND U4908 ( .A(n4650), .B(n4649), .Z(n4777) );
  NANDN U4909 ( .A(n19116), .B(n4651), .Z(n4653) );
  XOR U4910 ( .A(b[25]), .B(a[22]), .Z(n4794) );
  NANDN U4911 ( .A(n19179), .B(n4794), .Z(n4652) );
  NAND U4912 ( .A(n4653), .B(n4652), .Z(n4776) );
  XNOR U4913 ( .A(n4777), .B(n4776), .Z(n4778) );
  XOR U4914 ( .A(n4779), .B(n4778), .Z(n4747) );
  XNOR U4915 ( .A(n4746), .B(n4747), .Z(n4748) );
  NANDN U4916 ( .A(n18113), .B(n4654), .Z(n4656) );
  XOR U4917 ( .A(b[13]), .B(a[34]), .Z(n4797) );
  NANDN U4918 ( .A(n18229), .B(n4797), .Z(n4655) );
  AND U4919 ( .A(n4656), .B(n4655), .Z(n4741) );
  NANDN U4920 ( .A(n17888), .B(n4657), .Z(n4659) );
  XOR U4921 ( .A(b[11]), .B(a[36]), .Z(n4800) );
  NANDN U4922 ( .A(n18025), .B(n4800), .Z(n4658) );
  NAND U4923 ( .A(n4659), .B(n4658), .Z(n4740) );
  XNOR U4924 ( .A(n4741), .B(n4740), .Z(n4742) );
  NANDN U4925 ( .A(n18487), .B(n4660), .Z(n4662) );
  XOR U4926 ( .A(b[15]), .B(a[32]), .Z(n4803) );
  NANDN U4927 ( .A(n18311), .B(n4803), .Z(n4661) );
  AND U4928 ( .A(n4662), .B(n4661), .Z(n4737) );
  NANDN U4929 ( .A(n18853), .B(n4663), .Z(n4665) );
  XOR U4930 ( .A(b[21]), .B(a[26]), .Z(n4806) );
  NANDN U4931 ( .A(n18926), .B(n4806), .Z(n4664) );
  AND U4932 ( .A(n4665), .B(n4664), .Z(n4735) );
  NANDN U4933 ( .A(n17613), .B(n4666), .Z(n4668) );
  XOR U4934 ( .A(b[9]), .B(a[38]), .Z(n4809) );
  NANDN U4935 ( .A(n17739), .B(n4809), .Z(n4667) );
  NAND U4936 ( .A(n4668), .B(n4667), .Z(n4734) );
  XNOR U4937 ( .A(n4735), .B(n4734), .Z(n4736) );
  XOR U4938 ( .A(n4737), .B(n4736), .Z(n4743) );
  XOR U4939 ( .A(n4742), .B(n4743), .Z(n4749) );
  XOR U4940 ( .A(n4748), .B(n4749), .Z(n4761) );
  XNOR U4941 ( .A(n4760), .B(n4761), .Z(n4692) );
  XNOR U4942 ( .A(n4693), .B(n4692), .Z(n4694) );
  XOR U4943 ( .A(n4695), .B(n4694), .Z(n4813) );
  XNOR U4944 ( .A(n4812), .B(n4813), .Z(n4814) );
  XNOR U4945 ( .A(n4815), .B(n4814), .Z(n4820) );
  XOR U4946 ( .A(n4821), .B(n4820), .Z(n4687) );
  NANDN U4947 ( .A(n4670), .B(n4669), .Z(n4674) );
  OR U4948 ( .A(n4672), .B(n4671), .Z(n4673) );
  AND U4949 ( .A(n4674), .B(n4673), .Z(n4686) );
  XNOR U4950 ( .A(n4687), .B(n4686), .Z(n4688) );
  XNOR U4951 ( .A(n4689), .B(n4688), .Z(n4680) );
  XNOR U4952 ( .A(n4681), .B(n4680), .Z(n4682) );
  XNOR U4953 ( .A(n4683), .B(n4682), .Z(n4824) );
  XNOR U4954 ( .A(sreg[142]), .B(n4824), .Z(n4826) );
  NANDN U4955 ( .A(sreg[141]), .B(n4675), .Z(n4679) );
  NAND U4956 ( .A(n4677), .B(n4676), .Z(n4678) );
  NAND U4957 ( .A(n4679), .B(n4678), .Z(n4825) );
  XNOR U4958 ( .A(n4826), .B(n4825), .Z(c[142]) );
  NANDN U4959 ( .A(n4681), .B(n4680), .Z(n4685) );
  NANDN U4960 ( .A(n4683), .B(n4682), .Z(n4684) );
  AND U4961 ( .A(n4685), .B(n4684), .Z(n4832) );
  NANDN U4962 ( .A(n4687), .B(n4686), .Z(n4691) );
  NANDN U4963 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U4964 ( .A(n4691), .B(n4690), .Z(n4830) );
  NANDN U4965 ( .A(n4693), .B(n4692), .Z(n4697) );
  NANDN U4966 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U4967 ( .A(n4697), .B(n4696), .Z(n4842) );
  NANDN U4968 ( .A(n4699), .B(n4698), .Z(n4703) );
  NAND U4969 ( .A(n4701), .B(n4700), .Z(n4702) );
  AND U4970 ( .A(n4703), .B(n4702), .Z(n4841) );
  XNOR U4971 ( .A(n4842), .B(n4841), .Z(n4844) );
  NANDN U4972 ( .A(n4705), .B(n4704), .Z(n4709) );
  NANDN U4973 ( .A(n4707), .B(n4706), .Z(n4708) );
  AND U4974 ( .A(n4709), .B(n4708), .Z(n4919) );
  NANDN U4975 ( .A(n19237), .B(n4710), .Z(n4712) );
  XOR U4976 ( .A(b[27]), .B(a[21]), .Z(n4865) );
  NANDN U4977 ( .A(n19277), .B(n4865), .Z(n4711) );
  AND U4978 ( .A(n4712), .B(n4711), .Z(n4926) );
  NANDN U4979 ( .A(n17072), .B(n4713), .Z(n4715) );
  XOR U4980 ( .A(b[5]), .B(a[43]), .Z(n4868) );
  NANDN U4981 ( .A(n17223), .B(n4868), .Z(n4714) );
  AND U4982 ( .A(n4715), .B(n4714), .Z(n4924) );
  NANDN U4983 ( .A(n18673), .B(n4716), .Z(n4718) );
  XOR U4984 ( .A(b[19]), .B(a[29]), .Z(n4871) );
  NANDN U4985 ( .A(n18758), .B(n4871), .Z(n4717) );
  NAND U4986 ( .A(n4718), .B(n4717), .Z(n4923) );
  XNOR U4987 ( .A(n4924), .B(n4923), .Z(n4925) );
  XNOR U4988 ( .A(n4926), .B(n4925), .Z(n4917) );
  NANDN U4989 ( .A(n19425), .B(n4719), .Z(n4721) );
  XOR U4990 ( .A(b[31]), .B(a[17]), .Z(n4874) );
  NANDN U4991 ( .A(n19426), .B(n4874), .Z(n4720) );
  AND U4992 ( .A(n4721), .B(n4720), .Z(n4886) );
  NANDN U4993 ( .A(n17067), .B(n4722), .Z(n4724) );
  XOR U4994 ( .A(b[3]), .B(a[45]), .Z(n4877) );
  NANDN U4995 ( .A(n17068), .B(n4877), .Z(n4723) );
  AND U4996 ( .A(n4724), .B(n4723), .Z(n4884) );
  NANDN U4997 ( .A(n18514), .B(n4725), .Z(n4727) );
  XOR U4998 ( .A(b[17]), .B(a[31]), .Z(n4880) );
  NANDN U4999 ( .A(n18585), .B(n4880), .Z(n4726) );
  NAND U5000 ( .A(n4727), .B(n4726), .Z(n4883) );
  XNOR U5001 ( .A(n4884), .B(n4883), .Z(n4885) );
  XOR U5002 ( .A(n4886), .B(n4885), .Z(n4918) );
  XOR U5003 ( .A(n4917), .B(n4918), .Z(n4920) );
  XOR U5004 ( .A(n4919), .B(n4920), .Z(n4854) );
  NANDN U5005 ( .A(n4729), .B(n4728), .Z(n4733) );
  NANDN U5006 ( .A(n4731), .B(n4730), .Z(n4732) );
  AND U5007 ( .A(n4733), .B(n4732), .Z(n4907) );
  NANDN U5008 ( .A(n4735), .B(n4734), .Z(n4739) );
  NANDN U5009 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U5010 ( .A(n4739), .B(n4738), .Z(n4908) );
  XNOR U5011 ( .A(n4907), .B(n4908), .Z(n4909) );
  NANDN U5012 ( .A(n4741), .B(n4740), .Z(n4745) );
  NANDN U5013 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U5014 ( .A(n4745), .B(n4744), .Z(n4910) );
  XNOR U5015 ( .A(n4909), .B(n4910), .Z(n4853) );
  XNOR U5016 ( .A(n4854), .B(n4853), .Z(n4856) );
  NANDN U5017 ( .A(n4747), .B(n4746), .Z(n4751) );
  NANDN U5018 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U5019 ( .A(n4751), .B(n4750), .Z(n4855) );
  XOR U5020 ( .A(n4856), .B(n4855), .Z(n4968) );
  NANDN U5021 ( .A(n4753), .B(n4752), .Z(n4757) );
  NANDN U5022 ( .A(n4755), .B(n4754), .Z(n4756) );
  AND U5023 ( .A(n4757), .B(n4756), .Z(n4965) );
  NANDN U5024 ( .A(n4759), .B(n4758), .Z(n4763) );
  NANDN U5025 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U5026 ( .A(n4763), .B(n4762), .Z(n4850) );
  NANDN U5027 ( .A(n4765), .B(n4764), .Z(n4769) );
  OR U5028 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U5029 ( .A(n4769), .B(n4768), .Z(n4848) );
  NANDN U5030 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U5031 ( .A(n4773), .B(n4772), .Z(n4774) );
  AND U5032 ( .A(n4775), .B(n4774), .Z(n4914) );
  NANDN U5033 ( .A(n4777), .B(n4776), .Z(n4781) );
  NANDN U5034 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U5035 ( .A(n4781), .B(n4780), .Z(n4913) );
  XNOR U5036 ( .A(n4914), .B(n4913), .Z(n4916) );
  NAND U5037 ( .A(b[0]), .B(a[47]), .Z(n4782) );
  XNOR U5038 ( .A(b[1]), .B(n4782), .Z(n4784) );
  NANDN U5039 ( .A(b[0]), .B(a[46]), .Z(n4783) );
  NAND U5040 ( .A(n4784), .B(n4783), .Z(n4862) );
  NANDN U5041 ( .A(n19394), .B(n4785), .Z(n4787) );
  XOR U5042 ( .A(b[29]), .B(a[19]), .Z(n4938) );
  NANDN U5043 ( .A(n19395), .B(n4938), .Z(n4786) );
  AND U5044 ( .A(n4787), .B(n4786), .Z(n4860) );
  AND U5045 ( .A(b[31]), .B(a[15]), .Z(n4859) );
  XNOR U5046 ( .A(n4860), .B(n4859), .Z(n4861) );
  XNOR U5047 ( .A(n4862), .B(n4861), .Z(n4902) );
  NANDN U5048 ( .A(n19005), .B(n4788), .Z(n4790) );
  XOR U5049 ( .A(b[23]), .B(a[25]), .Z(n4941) );
  NANDN U5050 ( .A(n19055), .B(n4941), .Z(n4789) );
  AND U5051 ( .A(n4790), .B(n4789), .Z(n4931) );
  NANDN U5052 ( .A(n17362), .B(n4791), .Z(n4793) );
  XOR U5053 ( .A(b[7]), .B(a[41]), .Z(n4944) );
  NANDN U5054 ( .A(n17522), .B(n4944), .Z(n4792) );
  AND U5055 ( .A(n4793), .B(n4792), .Z(n4930) );
  NANDN U5056 ( .A(n19116), .B(n4794), .Z(n4796) );
  XOR U5057 ( .A(b[25]), .B(a[23]), .Z(n4947) );
  NANDN U5058 ( .A(n19179), .B(n4947), .Z(n4795) );
  NAND U5059 ( .A(n4796), .B(n4795), .Z(n4929) );
  XOR U5060 ( .A(n4930), .B(n4929), .Z(n4932) );
  XOR U5061 ( .A(n4931), .B(n4932), .Z(n4901) );
  XOR U5062 ( .A(n4902), .B(n4901), .Z(n4904) );
  NANDN U5063 ( .A(n18113), .B(n4797), .Z(n4799) );
  XOR U5064 ( .A(b[13]), .B(a[35]), .Z(n4950) );
  NANDN U5065 ( .A(n18229), .B(n4950), .Z(n4798) );
  AND U5066 ( .A(n4799), .B(n4798), .Z(n4896) );
  NANDN U5067 ( .A(n17888), .B(n4800), .Z(n4802) );
  XOR U5068 ( .A(b[11]), .B(a[37]), .Z(n4953) );
  NANDN U5069 ( .A(n18025), .B(n4953), .Z(n4801) );
  NAND U5070 ( .A(n4802), .B(n4801), .Z(n4895) );
  XNOR U5071 ( .A(n4896), .B(n4895), .Z(n4898) );
  NANDN U5072 ( .A(n18487), .B(n4803), .Z(n4805) );
  XOR U5073 ( .A(b[15]), .B(a[33]), .Z(n4956) );
  NANDN U5074 ( .A(n18311), .B(n4956), .Z(n4804) );
  AND U5075 ( .A(n4805), .B(n4804), .Z(n4892) );
  NANDN U5076 ( .A(n18853), .B(n4806), .Z(n4808) );
  XOR U5077 ( .A(b[21]), .B(a[27]), .Z(n4959) );
  NANDN U5078 ( .A(n18926), .B(n4959), .Z(n4807) );
  AND U5079 ( .A(n4808), .B(n4807), .Z(n4890) );
  NANDN U5080 ( .A(n17613), .B(n4809), .Z(n4811) );
  XOR U5081 ( .A(b[9]), .B(a[39]), .Z(n4962) );
  NANDN U5082 ( .A(n17739), .B(n4962), .Z(n4810) );
  NAND U5083 ( .A(n4811), .B(n4810), .Z(n4889) );
  XNOR U5084 ( .A(n4890), .B(n4889), .Z(n4891) );
  XNOR U5085 ( .A(n4892), .B(n4891), .Z(n4897) );
  XOR U5086 ( .A(n4898), .B(n4897), .Z(n4903) );
  XOR U5087 ( .A(n4904), .B(n4903), .Z(n4915) );
  XOR U5088 ( .A(n4916), .B(n4915), .Z(n4847) );
  XNOR U5089 ( .A(n4848), .B(n4847), .Z(n4849) );
  XOR U5090 ( .A(n4850), .B(n4849), .Z(n4966) );
  XNOR U5091 ( .A(n4965), .B(n4966), .Z(n4967) );
  XNOR U5092 ( .A(n4968), .B(n4967), .Z(n4843) );
  XOR U5093 ( .A(n4844), .B(n4843), .Z(n4836) );
  NANDN U5094 ( .A(n4813), .B(n4812), .Z(n4817) );
  NANDN U5095 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U5096 ( .A(n4817), .B(n4816), .Z(n4835) );
  XNOR U5097 ( .A(n4836), .B(n4835), .Z(n4837) );
  NANDN U5098 ( .A(n4819), .B(n4818), .Z(n4823) );
  NAND U5099 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U5100 ( .A(n4823), .B(n4822), .Z(n4838) );
  XNOR U5101 ( .A(n4837), .B(n4838), .Z(n4829) );
  XNOR U5102 ( .A(n4830), .B(n4829), .Z(n4831) );
  XNOR U5103 ( .A(n4832), .B(n4831), .Z(n4971) );
  XNOR U5104 ( .A(sreg[143]), .B(n4971), .Z(n4973) );
  NANDN U5105 ( .A(sreg[142]), .B(n4824), .Z(n4828) );
  NAND U5106 ( .A(n4826), .B(n4825), .Z(n4827) );
  NAND U5107 ( .A(n4828), .B(n4827), .Z(n4972) );
  XNOR U5108 ( .A(n4973), .B(n4972), .Z(c[143]) );
  NANDN U5109 ( .A(n4830), .B(n4829), .Z(n4834) );
  NANDN U5110 ( .A(n4832), .B(n4831), .Z(n4833) );
  AND U5111 ( .A(n4834), .B(n4833), .Z(n4979) );
  NANDN U5112 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U5113 ( .A(n4838), .B(n4837), .Z(n4839) );
  AND U5114 ( .A(n4840), .B(n4839), .Z(n4977) );
  NANDN U5115 ( .A(n4842), .B(n4841), .Z(n4846) );
  NAND U5116 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U5117 ( .A(n4846), .B(n4845), .Z(n4984) );
  NANDN U5118 ( .A(n4848), .B(n4847), .Z(n4852) );
  NANDN U5119 ( .A(n4850), .B(n4849), .Z(n4851) );
  AND U5120 ( .A(n4852), .B(n4851), .Z(n4989) );
  NANDN U5121 ( .A(n4854), .B(n4853), .Z(n4858) );
  NAND U5122 ( .A(n4856), .B(n4855), .Z(n4857) );
  AND U5123 ( .A(n4858), .B(n4857), .Z(n4988) );
  XNOR U5124 ( .A(n4989), .B(n4988), .Z(n4991) );
  NANDN U5125 ( .A(n4860), .B(n4859), .Z(n4864) );
  NANDN U5126 ( .A(n4862), .B(n4861), .Z(n4863) );
  AND U5127 ( .A(n4864), .B(n4863), .Z(n5056) );
  NANDN U5128 ( .A(n19237), .B(n4865), .Z(n4867) );
  XOR U5129 ( .A(b[27]), .B(a[22]), .Z(n5000) );
  NANDN U5130 ( .A(n19277), .B(n5000), .Z(n4866) );
  AND U5131 ( .A(n4867), .B(n4866), .Z(n5063) );
  NANDN U5132 ( .A(n17072), .B(n4868), .Z(n4870) );
  XOR U5133 ( .A(b[5]), .B(a[44]), .Z(n5003) );
  NANDN U5134 ( .A(n17223), .B(n5003), .Z(n4869) );
  AND U5135 ( .A(n4870), .B(n4869), .Z(n5061) );
  NANDN U5136 ( .A(n18673), .B(n4871), .Z(n4873) );
  XOR U5137 ( .A(b[19]), .B(a[30]), .Z(n5006) );
  NANDN U5138 ( .A(n18758), .B(n5006), .Z(n4872) );
  NAND U5139 ( .A(n4873), .B(n4872), .Z(n5060) );
  XNOR U5140 ( .A(n5061), .B(n5060), .Z(n5062) );
  XNOR U5141 ( .A(n5063), .B(n5062), .Z(n5054) );
  NANDN U5142 ( .A(n19425), .B(n4874), .Z(n4876) );
  XOR U5143 ( .A(b[31]), .B(a[18]), .Z(n5009) );
  NANDN U5144 ( .A(n19426), .B(n5009), .Z(n4875) );
  AND U5145 ( .A(n4876), .B(n4875), .Z(n5021) );
  NANDN U5146 ( .A(n17067), .B(n4877), .Z(n4879) );
  XOR U5147 ( .A(b[3]), .B(a[46]), .Z(n5012) );
  NANDN U5148 ( .A(n17068), .B(n5012), .Z(n4878) );
  AND U5149 ( .A(n4879), .B(n4878), .Z(n5019) );
  NANDN U5150 ( .A(n18514), .B(n4880), .Z(n4882) );
  XOR U5151 ( .A(b[17]), .B(a[32]), .Z(n5015) );
  NANDN U5152 ( .A(n18585), .B(n5015), .Z(n4881) );
  NAND U5153 ( .A(n4882), .B(n4881), .Z(n5018) );
  XNOR U5154 ( .A(n5019), .B(n5018), .Z(n5020) );
  XOR U5155 ( .A(n5021), .B(n5020), .Z(n5055) );
  XOR U5156 ( .A(n5054), .B(n5055), .Z(n5057) );
  XOR U5157 ( .A(n5056), .B(n5057), .Z(n5103) );
  NANDN U5158 ( .A(n4884), .B(n4883), .Z(n4888) );
  NANDN U5159 ( .A(n4886), .B(n4885), .Z(n4887) );
  AND U5160 ( .A(n4888), .B(n4887), .Z(n5042) );
  NANDN U5161 ( .A(n4890), .B(n4889), .Z(n4894) );
  NANDN U5162 ( .A(n4892), .B(n4891), .Z(n4893) );
  NAND U5163 ( .A(n4894), .B(n4893), .Z(n5043) );
  XNOR U5164 ( .A(n5042), .B(n5043), .Z(n5044) );
  NANDN U5165 ( .A(n4896), .B(n4895), .Z(n4900) );
  NAND U5166 ( .A(n4898), .B(n4897), .Z(n4899) );
  NAND U5167 ( .A(n4900), .B(n4899), .Z(n5045) );
  XNOR U5168 ( .A(n5044), .B(n5045), .Z(n5102) );
  XNOR U5169 ( .A(n5103), .B(n5102), .Z(n5105) );
  NAND U5170 ( .A(n4902), .B(n4901), .Z(n4906) );
  NAND U5171 ( .A(n4904), .B(n4903), .Z(n4905) );
  AND U5172 ( .A(n4906), .B(n4905), .Z(n5104) );
  XOR U5173 ( .A(n5105), .B(n5104), .Z(n5117) );
  NANDN U5174 ( .A(n4908), .B(n4907), .Z(n4912) );
  NANDN U5175 ( .A(n4910), .B(n4909), .Z(n4911) );
  AND U5176 ( .A(n4912), .B(n4911), .Z(n5114) );
  NANDN U5177 ( .A(n4918), .B(n4917), .Z(n4922) );
  OR U5178 ( .A(n4920), .B(n4919), .Z(n4921) );
  AND U5179 ( .A(n4922), .B(n4921), .Z(n5109) );
  NANDN U5180 ( .A(n4924), .B(n4923), .Z(n4928) );
  NANDN U5181 ( .A(n4926), .B(n4925), .Z(n4927) );
  AND U5182 ( .A(n4928), .B(n4927), .Z(n5049) );
  NANDN U5183 ( .A(n4930), .B(n4929), .Z(n4934) );
  OR U5184 ( .A(n4932), .B(n4931), .Z(n4933) );
  NAND U5185 ( .A(n4934), .B(n4933), .Z(n5048) );
  XNOR U5186 ( .A(n5049), .B(n5048), .Z(n5050) );
  NAND U5187 ( .A(b[0]), .B(a[48]), .Z(n4935) );
  XNOR U5188 ( .A(b[1]), .B(n4935), .Z(n4937) );
  NANDN U5189 ( .A(b[0]), .B(a[47]), .Z(n4936) );
  NAND U5190 ( .A(n4937), .B(n4936), .Z(n4997) );
  NANDN U5191 ( .A(n19394), .B(n4938), .Z(n4940) );
  XOR U5192 ( .A(b[29]), .B(a[20]), .Z(n5072) );
  NANDN U5193 ( .A(n19395), .B(n5072), .Z(n4939) );
  AND U5194 ( .A(n4940), .B(n4939), .Z(n4995) );
  AND U5195 ( .A(b[31]), .B(a[16]), .Z(n4994) );
  XNOR U5196 ( .A(n4995), .B(n4994), .Z(n4996) );
  XNOR U5197 ( .A(n4997), .B(n4996), .Z(n5036) );
  NANDN U5198 ( .A(n19005), .B(n4941), .Z(n4943) );
  XOR U5199 ( .A(b[23]), .B(a[26]), .Z(n5078) );
  NANDN U5200 ( .A(n19055), .B(n5078), .Z(n4942) );
  AND U5201 ( .A(n4943), .B(n4942), .Z(n5069) );
  NANDN U5202 ( .A(n17362), .B(n4944), .Z(n4946) );
  XOR U5203 ( .A(b[7]), .B(a[42]), .Z(n5081) );
  NANDN U5204 ( .A(n17522), .B(n5081), .Z(n4945) );
  AND U5205 ( .A(n4946), .B(n4945), .Z(n5067) );
  NANDN U5206 ( .A(n19116), .B(n4947), .Z(n4949) );
  XOR U5207 ( .A(b[25]), .B(a[24]), .Z(n5084) );
  NANDN U5208 ( .A(n19179), .B(n5084), .Z(n4948) );
  NAND U5209 ( .A(n4949), .B(n4948), .Z(n5066) );
  XNOR U5210 ( .A(n5067), .B(n5066), .Z(n5068) );
  XOR U5211 ( .A(n5069), .B(n5068), .Z(n5037) );
  XNOR U5212 ( .A(n5036), .B(n5037), .Z(n5038) );
  NANDN U5213 ( .A(n18113), .B(n4950), .Z(n4952) );
  XOR U5214 ( .A(b[13]), .B(a[36]), .Z(n5087) );
  NANDN U5215 ( .A(n18229), .B(n5087), .Z(n4951) );
  AND U5216 ( .A(n4952), .B(n4951), .Z(n5031) );
  NANDN U5217 ( .A(n17888), .B(n4953), .Z(n4955) );
  XOR U5218 ( .A(b[11]), .B(a[38]), .Z(n5090) );
  NANDN U5219 ( .A(n18025), .B(n5090), .Z(n4954) );
  NAND U5220 ( .A(n4955), .B(n4954), .Z(n5030) );
  XNOR U5221 ( .A(n5031), .B(n5030), .Z(n5032) );
  NANDN U5222 ( .A(n18487), .B(n4956), .Z(n4958) );
  XOR U5223 ( .A(b[15]), .B(a[34]), .Z(n5093) );
  NANDN U5224 ( .A(n18311), .B(n5093), .Z(n4957) );
  AND U5225 ( .A(n4958), .B(n4957), .Z(n5027) );
  NANDN U5226 ( .A(n18853), .B(n4959), .Z(n4961) );
  XOR U5227 ( .A(b[21]), .B(a[28]), .Z(n5096) );
  NANDN U5228 ( .A(n18926), .B(n5096), .Z(n4960) );
  AND U5229 ( .A(n4961), .B(n4960), .Z(n5025) );
  NANDN U5230 ( .A(n17613), .B(n4962), .Z(n4964) );
  XOR U5231 ( .A(b[9]), .B(a[40]), .Z(n5099) );
  NANDN U5232 ( .A(n17739), .B(n5099), .Z(n4963) );
  NAND U5233 ( .A(n4964), .B(n4963), .Z(n5024) );
  XNOR U5234 ( .A(n5025), .B(n5024), .Z(n5026) );
  XOR U5235 ( .A(n5027), .B(n5026), .Z(n5033) );
  XOR U5236 ( .A(n5032), .B(n5033), .Z(n5039) );
  XOR U5237 ( .A(n5038), .B(n5039), .Z(n5051) );
  XNOR U5238 ( .A(n5050), .B(n5051), .Z(n5108) );
  XNOR U5239 ( .A(n5109), .B(n5108), .Z(n5110) );
  XOR U5240 ( .A(n5111), .B(n5110), .Z(n5115) );
  XNOR U5241 ( .A(n5114), .B(n5115), .Z(n5116) );
  XNOR U5242 ( .A(n5117), .B(n5116), .Z(n4990) );
  XOR U5243 ( .A(n4991), .B(n4990), .Z(n4983) );
  NANDN U5244 ( .A(n4966), .B(n4965), .Z(n4970) );
  NANDN U5245 ( .A(n4968), .B(n4967), .Z(n4969) );
  AND U5246 ( .A(n4970), .B(n4969), .Z(n4982) );
  XOR U5247 ( .A(n4983), .B(n4982), .Z(n4985) );
  XNOR U5248 ( .A(n4984), .B(n4985), .Z(n4976) );
  XNOR U5249 ( .A(n4977), .B(n4976), .Z(n4978) );
  XNOR U5250 ( .A(n4979), .B(n4978), .Z(n5120) );
  XNOR U5251 ( .A(sreg[144]), .B(n5120), .Z(n5122) );
  NANDN U5252 ( .A(sreg[143]), .B(n4971), .Z(n4975) );
  NAND U5253 ( .A(n4973), .B(n4972), .Z(n4974) );
  NAND U5254 ( .A(n4975), .B(n4974), .Z(n5121) );
  XNOR U5255 ( .A(n5122), .B(n5121), .Z(c[144]) );
  NANDN U5256 ( .A(n4977), .B(n4976), .Z(n4981) );
  NANDN U5257 ( .A(n4979), .B(n4978), .Z(n4980) );
  AND U5258 ( .A(n4981), .B(n4980), .Z(n5128) );
  NANDN U5259 ( .A(n4983), .B(n4982), .Z(n4987) );
  NANDN U5260 ( .A(n4985), .B(n4984), .Z(n4986) );
  AND U5261 ( .A(n4987), .B(n4986), .Z(n5126) );
  NANDN U5262 ( .A(n4989), .B(n4988), .Z(n4993) );
  NAND U5263 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U5264 ( .A(n4993), .B(n4992), .Z(n5133) );
  NANDN U5265 ( .A(n4995), .B(n4994), .Z(n4999) );
  NANDN U5266 ( .A(n4997), .B(n4996), .Z(n4998) );
  AND U5267 ( .A(n4999), .B(n4998), .Z(n5215) );
  NANDN U5268 ( .A(n19237), .B(n5000), .Z(n5002) );
  XOR U5269 ( .A(b[27]), .B(a[23]), .Z(n5161) );
  NANDN U5270 ( .A(n19277), .B(n5161), .Z(n5001) );
  AND U5271 ( .A(n5002), .B(n5001), .Z(n5222) );
  NANDN U5272 ( .A(n17072), .B(n5003), .Z(n5005) );
  XOR U5273 ( .A(b[5]), .B(a[45]), .Z(n5164) );
  NANDN U5274 ( .A(n17223), .B(n5164), .Z(n5004) );
  AND U5275 ( .A(n5005), .B(n5004), .Z(n5220) );
  NANDN U5276 ( .A(n18673), .B(n5006), .Z(n5008) );
  XOR U5277 ( .A(b[19]), .B(a[31]), .Z(n5167) );
  NANDN U5278 ( .A(n18758), .B(n5167), .Z(n5007) );
  NAND U5279 ( .A(n5008), .B(n5007), .Z(n5219) );
  XNOR U5280 ( .A(n5220), .B(n5219), .Z(n5221) );
  XNOR U5281 ( .A(n5222), .B(n5221), .Z(n5213) );
  NANDN U5282 ( .A(n19425), .B(n5009), .Z(n5011) );
  XOR U5283 ( .A(b[31]), .B(a[19]), .Z(n5170) );
  NANDN U5284 ( .A(n19426), .B(n5170), .Z(n5010) );
  AND U5285 ( .A(n5011), .B(n5010), .Z(n5182) );
  NANDN U5286 ( .A(n17067), .B(n5012), .Z(n5014) );
  XOR U5287 ( .A(b[3]), .B(a[47]), .Z(n5173) );
  NANDN U5288 ( .A(n17068), .B(n5173), .Z(n5013) );
  AND U5289 ( .A(n5014), .B(n5013), .Z(n5180) );
  NANDN U5290 ( .A(n18514), .B(n5015), .Z(n5017) );
  XOR U5291 ( .A(b[17]), .B(a[33]), .Z(n5176) );
  NANDN U5292 ( .A(n18585), .B(n5176), .Z(n5016) );
  NAND U5293 ( .A(n5017), .B(n5016), .Z(n5179) );
  XNOR U5294 ( .A(n5180), .B(n5179), .Z(n5181) );
  XOR U5295 ( .A(n5182), .B(n5181), .Z(n5214) );
  XOR U5296 ( .A(n5213), .B(n5214), .Z(n5216) );
  XOR U5297 ( .A(n5215), .B(n5216), .Z(n5150) );
  NANDN U5298 ( .A(n5019), .B(n5018), .Z(n5023) );
  NANDN U5299 ( .A(n5021), .B(n5020), .Z(n5022) );
  AND U5300 ( .A(n5023), .B(n5022), .Z(n5203) );
  NANDN U5301 ( .A(n5025), .B(n5024), .Z(n5029) );
  NANDN U5302 ( .A(n5027), .B(n5026), .Z(n5028) );
  NAND U5303 ( .A(n5029), .B(n5028), .Z(n5204) );
  XNOR U5304 ( .A(n5203), .B(n5204), .Z(n5205) );
  NANDN U5305 ( .A(n5031), .B(n5030), .Z(n5035) );
  NANDN U5306 ( .A(n5033), .B(n5032), .Z(n5034) );
  NAND U5307 ( .A(n5035), .B(n5034), .Z(n5206) );
  XNOR U5308 ( .A(n5205), .B(n5206), .Z(n5149) );
  XNOR U5309 ( .A(n5150), .B(n5149), .Z(n5152) );
  NANDN U5310 ( .A(n5037), .B(n5036), .Z(n5041) );
  NANDN U5311 ( .A(n5039), .B(n5038), .Z(n5040) );
  AND U5312 ( .A(n5041), .B(n5040), .Z(n5151) );
  XOR U5313 ( .A(n5152), .B(n5151), .Z(n5263) );
  NANDN U5314 ( .A(n5043), .B(n5042), .Z(n5047) );
  NANDN U5315 ( .A(n5045), .B(n5044), .Z(n5046) );
  AND U5316 ( .A(n5047), .B(n5046), .Z(n5261) );
  NANDN U5317 ( .A(n5049), .B(n5048), .Z(n5053) );
  NANDN U5318 ( .A(n5051), .B(n5050), .Z(n5052) );
  AND U5319 ( .A(n5053), .B(n5052), .Z(n5146) );
  NANDN U5320 ( .A(n5055), .B(n5054), .Z(n5059) );
  OR U5321 ( .A(n5057), .B(n5056), .Z(n5058) );
  AND U5322 ( .A(n5059), .B(n5058), .Z(n5144) );
  NANDN U5323 ( .A(n5061), .B(n5060), .Z(n5065) );
  NANDN U5324 ( .A(n5063), .B(n5062), .Z(n5064) );
  AND U5325 ( .A(n5065), .B(n5064), .Z(n5210) );
  NANDN U5326 ( .A(n5067), .B(n5066), .Z(n5071) );
  NANDN U5327 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND U5328 ( .A(n5071), .B(n5070), .Z(n5209) );
  XNOR U5329 ( .A(n5210), .B(n5209), .Z(n5212) );
  NANDN U5330 ( .A(n19394), .B(n5072), .Z(n5074) );
  XOR U5331 ( .A(b[29]), .B(a[21]), .Z(n5234) );
  NANDN U5332 ( .A(n19395), .B(n5234), .Z(n5073) );
  AND U5333 ( .A(n5074), .B(n5073), .Z(n5156) );
  AND U5334 ( .A(b[31]), .B(a[17]), .Z(n5155) );
  XNOR U5335 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U5336 ( .A(b[0]), .B(a[49]), .Z(n5075) );
  XNOR U5337 ( .A(b[1]), .B(n5075), .Z(n5077) );
  NANDN U5338 ( .A(b[0]), .B(a[48]), .Z(n5076) );
  NAND U5339 ( .A(n5077), .B(n5076), .Z(n5158) );
  XNOR U5340 ( .A(n5157), .B(n5158), .Z(n5198) );
  NANDN U5341 ( .A(n19005), .B(n5078), .Z(n5080) );
  XOR U5342 ( .A(b[23]), .B(a[27]), .Z(n5237) );
  NANDN U5343 ( .A(n19055), .B(n5237), .Z(n5079) );
  AND U5344 ( .A(n5080), .B(n5079), .Z(n5227) );
  NANDN U5345 ( .A(n17362), .B(n5081), .Z(n5083) );
  XOR U5346 ( .A(b[7]), .B(a[43]), .Z(n5240) );
  NANDN U5347 ( .A(n17522), .B(n5240), .Z(n5082) );
  AND U5348 ( .A(n5083), .B(n5082), .Z(n5226) );
  NANDN U5349 ( .A(n19116), .B(n5084), .Z(n5086) );
  XOR U5350 ( .A(b[25]), .B(a[25]), .Z(n5243) );
  NANDN U5351 ( .A(n19179), .B(n5243), .Z(n5085) );
  NAND U5352 ( .A(n5086), .B(n5085), .Z(n5225) );
  XOR U5353 ( .A(n5226), .B(n5225), .Z(n5228) );
  XOR U5354 ( .A(n5227), .B(n5228), .Z(n5197) );
  XOR U5355 ( .A(n5198), .B(n5197), .Z(n5200) );
  NANDN U5356 ( .A(n18113), .B(n5087), .Z(n5089) );
  XOR U5357 ( .A(b[13]), .B(a[37]), .Z(n5246) );
  NANDN U5358 ( .A(n18229), .B(n5246), .Z(n5088) );
  AND U5359 ( .A(n5089), .B(n5088), .Z(n5192) );
  NANDN U5360 ( .A(n17888), .B(n5090), .Z(n5092) );
  XOR U5361 ( .A(b[11]), .B(a[39]), .Z(n5249) );
  NANDN U5362 ( .A(n18025), .B(n5249), .Z(n5091) );
  NAND U5363 ( .A(n5092), .B(n5091), .Z(n5191) );
  XNOR U5364 ( .A(n5192), .B(n5191), .Z(n5194) );
  NANDN U5365 ( .A(n18487), .B(n5093), .Z(n5095) );
  XOR U5366 ( .A(b[15]), .B(a[35]), .Z(n5252) );
  NANDN U5367 ( .A(n18311), .B(n5252), .Z(n5094) );
  AND U5368 ( .A(n5095), .B(n5094), .Z(n5188) );
  NANDN U5369 ( .A(n18853), .B(n5096), .Z(n5098) );
  XOR U5370 ( .A(b[21]), .B(a[29]), .Z(n5255) );
  NANDN U5371 ( .A(n18926), .B(n5255), .Z(n5097) );
  AND U5372 ( .A(n5098), .B(n5097), .Z(n5186) );
  NANDN U5373 ( .A(n17613), .B(n5099), .Z(n5101) );
  XOR U5374 ( .A(b[9]), .B(a[41]), .Z(n5258) );
  NANDN U5375 ( .A(n17739), .B(n5258), .Z(n5100) );
  NAND U5376 ( .A(n5101), .B(n5100), .Z(n5185) );
  XNOR U5377 ( .A(n5186), .B(n5185), .Z(n5187) );
  XNOR U5378 ( .A(n5188), .B(n5187), .Z(n5193) );
  XOR U5379 ( .A(n5194), .B(n5193), .Z(n5199) );
  XOR U5380 ( .A(n5200), .B(n5199), .Z(n5211) );
  XOR U5381 ( .A(n5212), .B(n5211), .Z(n5143) );
  XNOR U5382 ( .A(n5144), .B(n5143), .Z(n5145) );
  XOR U5383 ( .A(n5146), .B(n5145), .Z(n5262) );
  XOR U5384 ( .A(n5261), .B(n5262), .Z(n5264) );
  XOR U5385 ( .A(n5263), .B(n5264), .Z(n5140) );
  NANDN U5386 ( .A(n5103), .B(n5102), .Z(n5107) );
  NAND U5387 ( .A(n5105), .B(n5104), .Z(n5106) );
  AND U5388 ( .A(n5107), .B(n5106), .Z(n5138) );
  NANDN U5389 ( .A(n5109), .B(n5108), .Z(n5113) );
  NANDN U5390 ( .A(n5111), .B(n5110), .Z(n5112) );
  AND U5391 ( .A(n5113), .B(n5112), .Z(n5137) );
  XNOR U5392 ( .A(n5138), .B(n5137), .Z(n5139) );
  XNOR U5393 ( .A(n5140), .B(n5139), .Z(n5131) );
  NANDN U5394 ( .A(n5115), .B(n5114), .Z(n5119) );
  NANDN U5395 ( .A(n5117), .B(n5116), .Z(n5118) );
  NAND U5396 ( .A(n5119), .B(n5118), .Z(n5132) );
  XOR U5397 ( .A(n5131), .B(n5132), .Z(n5134) );
  XNOR U5398 ( .A(n5133), .B(n5134), .Z(n5125) );
  XNOR U5399 ( .A(n5126), .B(n5125), .Z(n5127) );
  XNOR U5400 ( .A(n5128), .B(n5127), .Z(n5267) );
  XNOR U5401 ( .A(sreg[145]), .B(n5267), .Z(n5269) );
  NANDN U5402 ( .A(sreg[144]), .B(n5120), .Z(n5124) );
  NAND U5403 ( .A(n5122), .B(n5121), .Z(n5123) );
  NAND U5404 ( .A(n5124), .B(n5123), .Z(n5268) );
  XNOR U5405 ( .A(n5269), .B(n5268), .Z(c[145]) );
  NANDN U5406 ( .A(n5126), .B(n5125), .Z(n5130) );
  NANDN U5407 ( .A(n5128), .B(n5127), .Z(n5129) );
  AND U5408 ( .A(n5130), .B(n5129), .Z(n5275) );
  NANDN U5409 ( .A(n5132), .B(n5131), .Z(n5136) );
  NANDN U5410 ( .A(n5134), .B(n5133), .Z(n5135) );
  AND U5411 ( .A(n5136), .B(n5135), .Z(n5273) );
  NANDN U5412 ( .A(n5138), .B(n5137), .Z(n5142) );
  NANDN U5413 ( .A(n5140), .B(n5139), .Z(n5141) );
  AND U5414 ( .A(n5142), .B(n5141), .Z(n5281) );
  NANDN U5415 ( .A(n5144), .B(n5143), .Z(n5148) );
  NANDN U5416 ( .A(n5146), .B(n5145), .Z(n5147) );
  AND U5417 ( .A(n5148), .B(n5147), .Z(n5285) );
  NANDN U5418 ( .A(n5150), .B(n5149), .Z(n5154) );
  NAND U5419 ( .A(n5152), .B(n5151), .Z(n5153) );
  AND U5420 ( .A(n5154), .B(n5153), .Z(n5284) );
  XNOR U5421 ( .A(n5285), .B(n5284), .Z(n5287) );
  NANDN U5422 ( .A(n5156), .B(n5155), .Z(n5160) );
  NANDN U5423 ( .A(n5158), .B(n5157), .Z(n5159) );
  AND U5424 ( .A(n5160), .B(n5159), .Z(n5350) );
  NANDN U5425 ( .A(n19237), .B(n5161), .Z(n5163) );
  XOR U5426 ( .A(b[27]), .B(a[24]), .Z(n5296) );
  NANDN U5427 ( .A(n19277), .B(n5296), .Z(n5162) );
  AND U5428 ( .A(n5163), .B(n5162), .Z(n5357) );
  NANDN U5429 ( .A(n17072), .B(n5164), .Z(n5166) );
  XOR U5430 ( .A(b[5]), .B(a[46]), .Z(n5299) );
  NANDN U5431 ( .A(n17223), .B(n5299), .Z(n5165) );
  AND U5432 ( .A(n5166), .B(n5165), .Z(n5355) );
  NANDN U5433 ( .A(n18673), .B(n5167), .Z(n5169) );
  XOR U5434 ( .A(b[19]), .B(a[32]), .Z(n5302) );
  NANDN U5435 ( .A(n18758), .B(n5302), .Z(n5168) );
  NAND U5436 ( .A(n5169), .B(n5168), .Z(n5354) );
  XNOR U5437 ( .A(n5355), .B(n5354), .Z(n5356) );
  XNOR U5438 ( .A(n5357), .B(n5356), .Z(n5348) );
  NANDN U5439 ( .A(n19425), .B(n5170), .Z(n5172) );
  XOR U5440 ( .A(b[31]), .B(a[20]), .Z(n5305) );
  NANDN U5441 ( .A(n19426), .B(n5305), .Z(n5171) );
  AND U5442 ( .A(n5172), .B(n5171), .Z(n5317) );
  NANDN U5443 ( .A(n17067), .B(n5173), .Z(n5175) );
  XOR U5444 ( .A(b[3]), .B(a[48]), .Z(n5308) );
  NANDN U5445 ( .A(n17068), .B(n5308), .Z(n5174) );
  AND U5446 ( .A(n5175), .B(n5174), .Z(n5315) );
  NANDN U5447 ( .A(n18514), .B(n5176), .Z(n5178) );
  XOR U5448 ( .A(b[17]), .B(a[34]), .Z(n5311) );
  NANDN U5449 ( .A(n18585), .B(n5311), .Z(n5177) );
  NAND U5450 ( .A(n5178), .B(n5177), .Z(n5314) );
  XNOR U5451 ( .A(n5315), .B(n5314), .Z(n5316) );
  XOR U5452 ( .A(n5317), .B(n5316), .Z(n5349) );
  XOR U5453 ( .A(n5348), .B(n5349), .Z(n5351) );
  XOR U5454 ( .A(n5350), .B(n5351), .Z(n5397) );
  NANDN U5455 ( .A(n5180), .B(n5179), .Z(n5184) );
  NANDN U5456 ( .A(n5182), .B(n5181), .Z(n5183) );
  AND U5457 ( .A(n5184), .B(n5183), .Z(n5338) );
  NANDN U5458 ( .A(n5186), .B(n5185), .Z(n5190) );
  NANDN U5459 ( .A(n5188), .B(n5187), .Z(n5189) );
  NAND U5460 ( .A(n5190), .B(n5189), .Z(n5339) );
  XNOR U5461 ( .A(n5338), .B(n5339), .Z(n5340) );
  NANDN U5462 ( .A(n5192), .B(n5191), .Z(n5196) );
  NAND U5463 ( .A(n5194), .B(n5193), .Z(n5195) );
  NAND U5464 ( .A(n5196), .B(n5195), .Z(n5341) );
  XNOR U5465 ( .A(n5340), .B(n5341), .Z(n5396) );
  XNOR U5466 ( .A(n5397), .B(n5396), .Z(n5399) );
  NAND U5467 ( .A(n5198), .B(n5197), .Z(n5202) );
  NAND U5468 ( .A(n5200), .B(n5199), .Z(n5201) );
  AND U5469 ( .A(n5202), .B(n5201), .Z(n5398) );
  XOR U5470 ( .A(n5399), .B(n5398), .Z(n5411) );
  NANDN U5471 ( .A(n5204), .B(n5203), .Z(n5208) );
  NANDN U5472 ( .A(n5206), .B(n5205), .Z(n5207) );
  AND U5473 ( .A(n5208), .B(n5207), .Z(n5408) );
  NANDN U5474 ( .A(n5214), .B(n5213), .Z(n5218) );
  OR U5475 ( .A(n5216), .B(n5215), .Z(n5217) );
  AND U5476 ( .A(n5218), .B(n5217), .Z(n5403) );
  NANDN U5477 ( .A(n5220), .B(n5219), .Z(n5224) );
  NANDN U5478 ( .A(n5222), .B(n5221), .Z(n5223) );
  AND U5479 ( .A(n5224), .B(n5223), .Z(n5345) );
  NANDN U5480 ( .A(n5226), .B(n5225), .Z(n5230) );
  OR U5481 ( .A(n5228), .B(n5227), .Z(n5229) );
  NAND U5482 ( .A(n5230), .B(n5229), .Z(n5344) );
  XNOR U5483 ( .A(n5345), .B(n5344), .Z(n5347) );
  NAND U5484 ( .A(b[0]), .B(a[50]), .Z(n5231) );
  XNOR U5485 ( .A(b[1]), .B(n5231), .Z(n5233) );
  NANDN U5486 ( .A(b[0]), .B(a[49]), .Z(n5232) );
  NAND U5487 ( .A(n5233), .B(n5232), .Z(n5293) );
  NANDN U5488 ( .A(n19394), .B(n5234), .Z(n5236) );
  XOR U5489 ( .A(b[29]), .B(a[22]), .Z(n5369) );
  NANDN U5490 ( .A(n19395), .B(n5369), .Z(n5235) );
  AND U5491 ( .A(n5236), .B(n5235), .Z(n5291) );
  AND U5492 ( .A(b[31]), .B(a[18]), .Z(n5290) );
  XNOR U5493 ( .A(n5291), .B(n5290), .Z(n5292) );
  XNOR U5494 ( .A(n5293), .B(n5292), .Z(n5333) );
  NANDN U5495 ( .A(n19005), .B(n5237), .Z(n5239) );
  XOR U5496 ( .A(b[23]), .B(a[28]), .Z(n5372) );
  NANDN U5497 ( .A(n19055), .B(n5372), .Z(n5238) );
  AND U5498 ( .A(n5239), .B(n5238), .Z(n5362) );
  NANDN U5499 ( .A(n17362), .B(n5240), .Z(n5242) );
  XOR U5500 ( .A(b[7]), .B(a[44]), .Z(n5375) );
  NANDN U5501 ( .A(n17522), .B(n5375), .Z(n5241) );
  AND U5502 ( .A(n5242), .B(n5241), .Z(n5361) );
  NANDN U5503 ( .A(n19116), .B(n5243), .Z(n5245) );
  XOR U5504 ( .A(b[25]), .B(a[26]), .Z(n5378) );
  NANDN U5505 ( .A(n19179), .B(n5378), .Z(n5244) );
  NAND U5506 ( .A(n5245), .B(n5244), .Z(n5360) );
  XOR U5507 ( .A(n5361), .B(n5360), .Z(n5363) );
  XOR U5508 ( .A(n5362), .B(n5363), .Z(n5332) );
  XOR U5509 ( .A(n5333), .B(n5332), .Z(n5335) );
  NANDN U5510 ( .A(n18113), .B(n5246), .Z(n5248) );
  XOR U5511 ( .A(b[13]), .B(a[38]), .Z(n5381) );
  NANDN U5512 ( .A(n18229), .B(n5381), .Z(n5247) );
  AND U5513 ( .A(n5248), .B(n5247), .Z(n5327) );
  NANDN U5514 ( .A(n17888), .B(n5249), .Z(n5251) );
  XOR U5515 ( .A(b[11]), .B(a[40]), .Z(n5384) );
  NANDN U5516 ( .A(n18025), .B(n5384), .Z(n5250) );
  NAND U5517 ( .A(n5251), .B(n5250), .Z(n5326) );
  XNOR U5518 ( .A(n5327), .B(n5326), .Z(n5329) );
  NANDN U5519 ( .A(n18487), .B(n5252), .Z(n5254) );
  XOR U5520 ( .A(b[15]), .B(a[36]), .Z(n5387) );
  NANDN U5521 ( .A(n18311), .B(n5387), .Z(n5253) );
  AND U5522 ( .A(n5254), .B(n5253), .Z(n5323) );
  NANDN U5523 ( .A(n18853), .B(n5255), .Z(n5257) );
  XOR U5524 ( .A(b[21]), .B(a[30]), .Z(n5390) );
  NANDN U5525 ( .A(n18926), .B(n5390), .Z(n5256) );
  AND U5526 ( .A(n5257), .B(n5256), .Z(n5321) );
  NANDN U5527 ( .A(n17613), .B(n5258), .Z(n5260) );
  XOR U5528 ( .A(b[9]), .B(a[42]), .Z(n5393) );
  NANDN U5529 ( .A(n17739), .B(n5393), .Z(n5259) );
  NAND U5530 ( .A(n5260), .B(n5259), .Z(n5320) );
  XNOR U5531 ( .A(n5321), .B(n5320), .Z(n5322) );
  XNOR U5532 ( .A(n5323), .B(n5322), .Z(n5328) );
  XOR U5533 ( .A(n5329), .B(n5328), .Z(n5334) );
  XOR U5534 ( .A(n5335), .B(n5334), .Z(n5346) );
  XOR U5535 ( .A(n5347), .B(n5346), .Z(n5402) );
  XNOR U5536 ( .A(n5403), .B(n5402), .Z(n5404) );
  XOR U5537 ( .A(n5405), .B(n5404), .Z(n5409) );
  XNOR U5538 ( .A(n5408), .B(n5409), .Z(n5410) );
  XNOR U5539 ( .A(n5411), .B(n5410), .Z(n5286) );
  XOR U5540 ( .A(n5287), .B(n5286), .Z(n5279) );
  NANDN U5541 ( .A(n5262), .B(n5261), .Z(n5266) );
  OR U5542 ( .A(n5264), .B(n5263), .Z(n5265) );
  AND U5543 ( .A(n5266), .B(n5265), .Z(n5278) );
  XNOR U5544 ( .A(n5279), .B(n5278), .Z(n5280) );
  XNOR U5545 ( .A(n5281), .B(n5280), .Z(n5272) );
  XNOR U5546 ( .A(n5273), .B(n5272), .Z(n5274) );
  XNOR U5547 ( .A(n5275), .B(n5274), .Z(n5414) );
  XNOR U5548 ( .A(sreg[146]), .B(n5414), .Z(n5416) );
  NANDN U5549 ( .A(sreg[145]), .B(n5267), .Z(n5271) );
  NAND U5550 ( .A(n5269), .B(n5268), .Z(n5270) );
  NAND U5551 ( .A(n5271), .B(n5270), .Z(n5415) );
  XNOR U5552 ( .A(n5416), .B(n5415), .Z(c[146]) );
  NANDN U5553 ( .A(n5273), .B(n5272), .Z(n5277) );
  NANDN U5554 ( .A(n5275), .B(n5274), .Z(n5276) );
  AND U5555 ( .A(n5277), .B(n5276), .Z(n5422) );
  NANDN U5556 ( .A(n5279), .B(n5278), .Z(n5283) );
  NANDN U5557 ( .A(n5281), .B(n5280), .Z(n5282) );
  AND U5558 ( .A(n5283), .B(n5282), .Z(n5420) );
  NANDN U5559 ( .A(n5285), .B(n5284), .Z(n5289) );
  NAND U5560 ( .A(n5287), .B(n5286), .Z(n5288) );
  AND U5561 ( .A(n5289), .B(n5288), .Z(n5427) );
  NANDN U5562 ( .A(n5291), .B(n5290), .Z(n5295) );
  NANDN U5563 ( .A(n5293), .B(n5292), .Z(n5294) );
  AND U5564 ( .A(n5295), .B(n5294), .Z(n5499) );
  NANDN U5565 ( .A(n19237), .B(n5296), .Z(n5298) );
  XOR U5566 ( .A(b[27]), .B(a[25]), .Z(n5443) );
  NANDN U5567 ( .A(n19277), .B(n5443), .Z(n5297) );
  AND U5568 ( .A(n5298), .B(n5297), .Z(n5506) );
  NANDN U5569 ( .A(n17072), .B(n5299), .Z(n5301) );
  XOR U5570 ( .A(b[5]), .B(a[47]), .Z(n5446) );
  NANDN U5571 ( .A(n17223), .B(n5446), .Z(n5300) );
  AND U5572 ( .A(n5301), .B(n5300), .Z(n5504) );
  NANDN U5573 ( .A(n18673), .B(n5302), .Z(n5304) );
  XOR U5574 ( .A(b[19]), .B(a[33]), .Z(n5449) );
  NANDN U5575 ( .A(n18758), .B(n5449), .Z(n5303) );
  NAND U5576 ( .A(n5304), .B(n5303), .Z(n5503) );
  XNOR U5577 ( .A(n5504), .B(n5503), .Z(n5505) );
  XNOR U5578 ( .A(n5506), .B(n5505), .Z(n5497) );
  NANDN U5579 ( .A(n19425), .B(n5305), .Z(n5307) );
  XOR U5580 ( .A(b[31]), .B(a[21]), .Z(n5452) );
  NANDN U5581 ( .A(n19426), .B(n5452), .Z(n5306) );
  AND U5582 ( .A(n5307), .B(n5306), .Z(n5464) );
  NANDN U5583 ( .A(n17067), .B(n5308), .Z(n5310) );
  XOR U5584 ( .A(b[3]), .B(a[49]), .Z(n5455) );
  NANDN U5585 ( .A(n17068), .B(n5455), .Z(n5309) );
  AND U5586 ( .A(n5310), .B(n5309), .Z(n5462) );
  NANDN U5587 ( .A(n18514), .B(n5311), .Z(n5313) );
  XOR U5588 ( .A(b[17]), .B(a[35]), .Z(n5458) );
  NANDN U5589 ( .A(n18585), .B(n5458), .Z(n5312) );
  NAND U5590 ( .A(n5313), .B(n5312), .Z(n5461) );
  XNOR U5591 ( .A(n5462), .B(n5461), .Z(n5463) );
  XOR U5592 ( .A(n5464), .B(n5463), .Z(n5498) );
  XOR U5593 ( .A(n5497), .B(n5498), .Z(n5500) );
  XOR U5594 ( .A(n5499), .B(n5500), .Z(n5546) );
  NANDN U5595 ( .A(n5315), .B(n5314), .Z(n5319) );
  NANDN U5596 ( .A(n5317), .B(n5316), .Z(n5318) );
  AND U5597 ( .A(n5319), .B(n5318), .Z(n5485) );
  NANDN U5598 ( .A(n5321), .B(n5320), .Z(n5325) );
  NANDN U5599 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U5600 ( .A(n5325), .B(n5324), .Z(n5486) );
  XNOR U5601 ( .A(n5485), .B(n5486), .Z(n5487) );
  NANDN U5602 ( .A(n5327), .B(n5326), .Z(n5331) );
  NAND U5603 ( .A(n5329), .B(n5328), .Z(n5330) );
  NAND U5604 ( .A(n5331), .B(n5330), .Z(n5488) );
  XNOR U5605 ( .A(n5487), .B(n5488), .Z(n5545) );
  XNOR U5606 ( .A(n5546), .B(n5545), .Z(n5548) );
  NAND U5607 ( .A(n5333), .B(n5332), .Z(n5337) );
  NAND U5608 ( .A(n5335), .B(n5334), .Z(n5336) );
  AND U5609 ( .A(n5337), .B(n5336), .Z(n5547) );
  XOR U5610 ( .A(n5548), .B(n5547), .Z(n5559) );
  NANDN U5611 ( .A(n5339), .B(n5338), .Z(n5343) );
  NANDN U5612 ( .A(n5341), .B(n5340), .Z(n5342) );
  AND U5613 ( .A(n5343), .B(n5342), .Z(n5557) );
  NANDN U5614 ( .A(n5349), .B(n5348), .Z(n5353) );
  OR U5615 ( .A(n5351), .B(n5350), .Z(n5352) );
  AND U5616 ( .A(n5353), .B(n5352), .Z(n5552) );
  NANDN U5617 ( .A(n5355), .B(n5354), .Z(n5359) );
  NANDN U5618 ( .A(n5357), .B(n5356), .Z(n5358) );
  AND U5619 ( .A(n5359), .B(n5358), .Z(n5492) );
  NANDN U5620 ( .A(n5361), .B(n5360), .Z(n5365) );
  OR U5621 ( .A(n5363), .B(n5362), .Z(n5364) );
  NAND U5622 ( .A(n5365), .B(n5364), .Z(n5491) );
  XNOR U5623 ( .A(n5492), .B(n5491), .Z(n5493) );
  NAND U5624 ( .A(b[0]), .B(a[51]), .Z(n5366) );
  XNOR U5625 ( .A(b[1]), .B(n5366), .Z(n5368) );
  NANDN U5626 ( .A(b[0]), .B(a[50]), .Z(n5367) );
  NAND U5627 ( .A(n5368), .B(n5367), .Z(n5440) );
  NANDN U5628 ( .A(n19394), .B(n5369), .Z(n5371) );
  XOR U5629 ( .A(b[29]), .B(a[23]), .Z(n5518) );
  NANDN U5630 ( .A(n19395), .B(n5518), .Z(n5370) );
  AND U5631 ( .A(n5371), .B(n5370), .Z(n5438) );
  AND U5632 ( .A(b[31]), .B(a[19]), .Z(n5437) );
  XNOR U5633 ( .A(n5438), .B(n5437), .Z(n5439) );
  XNOR U5634 ( .A(n5440), .B(n5439), .Z(n5479) );
  NANDN U5635 ( .A(n19005), .B(n5372), .Z(n5374) );
  XOR U5636 ( .A(b[23]), .B(a[29]), .Z(n5521) );
  NANDN U5637 ( .A(n19055), .B(n5521), .Z(n5373) );
  AND U5638 ( .A(n5374), .B(n5373), .Z(n5512) );
  NANDN U5639 ( .A(n17362), .B(n5375), .Z(n5377) );
  XOR U5640 ( .A(b[7]), .B(a[45]), .Z(n5524) );
  NANDN U5641 ( .A(n17522), .B(n5524), .Z(n5376) );
  AND U5642 ( .A(n5377), .B(n5376), .Z(n5510) );
  NANDN U5643 ( .A(n19116), .B(n5378), .Z(n5380) );
  XOR U5644 ( .A(b[25]), .B(a[27]), .Z(n5527) );
  NANDN U5645 ( .A(n19179), .B(n5527), .Z(n5379) );
  NAND U5646 ( .A(n5380), .B(n5379), .Z(n5509) );
  XNOR U5647 ( .A(n5510), .B(n5509), .Z(n5511) );
  XOR U5648 ( .A(n5512), .B(n5511), .Z(n5480) );
  XNOR U5649 ( .A(n5479), .B(n5480), .Z(n5481) );
  NANDN U5650 ( .A(n18113), .B(n5381), .Z(n5383) );
  XOR U5651 ( .A(b[13]), .B(a[39]), .Z(n5530) );
  NANDN U5652 ( .A(n18229), .B(n5530), .Z(n5382) );
  AND U5653 ( .A(n5383), .B(n5382), .Z(n5474) );
  NANDN U5654 ( .A(n17888), .B(n5384), .Z(n5386) );
  XOR U5655 ( .A(b[11]), .B(a[41]), .Z(n5533) );
  NANDN U5656 ( .A(n18025), .B(n5533), .Z(n5385) );
  NAND U5657 ( .A(n5386), .B(n5385), .Z(n5473) );
  XNOR U5658 ( .A(n5474), .B(n5473), .Z(n5475) );
  NANDN U5659 ( .A(n18487), .B(n5387), .Z(n5389) );
  XOR U5660 ( .A(b[15]), .B(a[37]), .Z(n5536) );
  NANDN U5661 ( .A(n18311), .B(n5536), .Z(n5388) );
  AND U5662 ( .A(n5389), .B(n5388), .Z(n5470) );
  NANDN U5663 ( .A(n18853), .B(n5390), .Z(n5392) );
  XOR U5664 ( .A(b[21]), .B(a[31]), .Z(n5539) );
  NANDN U5665 ( .A(n18926), .B(n5539), .Z(n5391) );
  AND U5666 ( .A(n5392), .B(n5391), .Z(n5468) );
  NANDN U5667 ( .A(n17613), .B(n5393), .Z(n5395) );
  XOR U5668 ( .A(b[9]), .B(a[43]), .Z(n5542) );
  NANDN U5669 ( .A(n17739), .B(n5542), .Z(n5394) );
  NAND U5670 ( .A(n5395), .B(n5394), .Z(n5467) );
  XNOR U5671 ( .A(n5468), .B(n5467), .Z(n5469) );
  XOR U5672 ( .A(n5470), .B(n5469), .Z(n5476) );
  XOR U5673 ( .A(n5475), .B(n5476), .Z(n5482) );
  XOR U5674 ( .A(n5481), .B(n5482), .Z(n5494) );
  XNOR U5675 ( .A(n5493), .B(n5494), .Z(n5551) );
  XNOR U5676 ( .A(n5552), .B(n5551), .Z(n5553) );
  XOR U5677 ( .A(n5554), .B(n5553), .Z(n5558) );
  XOR U5678 ( .A(n5557), .B(n5558), .Z(n5560) );
  XOR U5679 ( .A(n5559), .B(n5560), .Z(n5434) );
  NANDN U5680 ( .A(n5397), .B(n5396), .Z(n5401) );
  NAND U5681 ( .A(n5399), .B(n5398), .Z(n5400) );
  AND U5682 ( .A(n5401), .B(n5400), .Z(n5432) );
  NANDN U5683 ( .A(n5403), .B(n5402), .Z(n5407) );
  NANDN U5684 ( .A(n5405), .B(n5404), .Z(n5406) );
  AND U5685 ( .A(n5407), .B(n5406), .Z(n5431) );
  XNOR U5686 ( .A(n5432), .B(n5431), .Z(n5433) );
  XNOR U5687 ( .A(n5434), .B(n5433), .Z(n5425) );
  NANDN U5688 ( .A(n5409), .B(n5408), .Z(n5413) );
  NANDN U5689 ( .A(n5411), .B(n5410), .Z(n5412) );
  NAND U5690 ( .A(n5413), .B(n5412), .Z(n5426) );
  XOR U5691 ( .A(n5425), .B(n5426), .Z(n5428) );
  XNOR U5692 ( .A(n5427), .B(n5428), .Z(n5419) );
  XNOR U5693 ( .A(n5420), .B(n5419), .Z(n5421) );
  XNOR U5694 ( .A(n5422), .B(n5421), .Z(n5563) );
  XNOR U5695 ( .A(sreg[147]), .B(n5563), .Z(n5565) );
  NANDN U5696 ( .A(sreg[146]), .B(n5414), .Z(n5418) );
  NAND U5697 ( .A(n5416), .B(n5415), .Z(n5417) );
  NAND U5698 ( .A(n5418), .B(n5417), .Z(n5564) );
  XNOR U5699 ( .A(n5565), .B(n5564), .Z(c[147]) );
  NANDN U5700 ( .A(n5420), .B(n5419), .Z(n5424) );
  NANDN U5701 ( .A(n5422), .B(n5421), .Z(n5423) );
  AND U5702 ( .A(n5424), .B(n5423), .Z(n5571) );
  NANDN U5703 ( .A(n5426), .B(n5425), .Z(n5430) );
  NANDN U5704 ( .A(n5428), .B(n5427), .Z(n5429) );
  AND U5705 ( .A(n5430), .B(n5429), .Z(n5569) );
  NANDN U5706 ( .A(n5432), .B(n5431), .Z(n5436) );
  NANDN U5707 ( .A(n5434), .B(n5433), .Z(n5435) );
  AND U5708 ( .A(n5436), .B(n5435), .Z(n5577) );
  NANDN U5709 ( .A(n5438), .B(n5437), .Z(n5442) );
  NANDN U5710 ( .A(n5440), .B(n5439), .Z(n5441) );
  AND U5711 ( .A(n5442), .B(n5441), .Z(n5660) );
  NANDN U5712 ( .A(n19237), .B(n5443), .Z(n5445) );
  XOR U5713 ( .A(b[27]), .B(a[26]), .Z(n5604) );
  NANDN U5714 ( .A(n19277), .B(n5604), .Z(n5444) );
  AND U5715 ( .A(n5445), .B(n5444), .Z(n5667) );
  NANDN U5716 ( .A(n17072), .B(n5446), .Z(n5448) );
  XOR U5717 ( .A(b[5]), .B(a[48]), .Z(n5607) );
  NANDN U5718 ( .A(n17223), .B(n5607), .Z(n5447) );
  AND U5719 ( .A(n5448), .B(n5447), .Z(n5665) );
  NANDN U5720 ( .A(n18673), .B(n5449), .Z(n5451) );
  XOR U5721 ( .A(b[19]), .B(a[34]), .Z(n5610) );
  NANDN U5722 ( .A(n18758), .B(n5610), .Z(n5450) );
  NAND U5723 ( .A(n5451), .B(n5450), .Z(n5664) );
  XNOR U5724 ( .A(n5665), .B(n5664), .Z(n5666) );
  XNOR U5725 ( .A(n5667), .B(n5666), .Z(n5658) );
  NANDN U5726 ( .A(n19425), .B(n5452), .Z(n5454) );
  XOR U5727 ( .A(b[31]), .B(a[22]), .Z(n5613) );
  NANDN U5728 ( .A(n19426), .B(n5613), .Z(n5453) );
  AND U5729 ( .A(n5454), .B(n5453), .Z(n5625) );
  NANDN U5730 ( .A(n17067), .B(n5455), .Z(n5457) );
  XOR U5731 ( .A(b[3]), .B(a[50]), .Z(n5616) );
  NANDN U5732 ( .A(n17068), .B(n5616), .Z(n5456) );
  AND U5733 ( .A(n5457), .B(n5456), .Z(n5623) );
  NANDN U5734 ( .A(n18514), .B(n5458), .Z(n5460) );
  XOR U5735 ( .A(b[17]), .B(a[36]), .Z(n5619) );
  NANDN U5736 ( .A(n18585), .B(n5619), .Z(n5459) );
  NAND U5737 ( .A(n5460), .B(n5459), .Z(n5622) );
  XNOR U5738 ( .A(n5623), .B(n5622), .Z(n5624) );
  XOR U5739 ( .A(n5625), .B(n5624), .Z(n5659) );
  XOR U5740 ( .A(n5658), .B(n5659), .Z(n5661) );
  XOR U5741 ( .A(n5660), .B(n5661), .Z(n5593) );
  NANDN U5742 ( .A(n5462), .B(n5461), .Z(n5466) );
  NANDN U5743 ( .A(n5464), .B(n5463), .Z(n5465) );
  AND U5744 ( .A(n5466), .B(n5465), .Z(n5646) );
  NANDN U5745 ( .A(n5468), .B(n5467), .Z(n5472) );
  NANDN U5746 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U5747 ( .A(n5472), .B(n5471), .Z(n5647) );
  XNOR U5748 ( .A(n5646), .B(n5647), .Z(n5648) );
  NANDN U5749 ( .A(n5474), .B(n5473), .Z(n5478) );
  NANDN U5750 ( .A(n5476), .B(n5475), .Z(n5477) );
  NAND U5751 ( .A(n5478), .B(n5477), .Z(n5649) );
  XNOR U5752 ( .A(n5648), .B(n5649), .Z(n5592) );
  XNOR U5753 ( .A(n5593), .B(n5592), .Z(n5595) );
  NANDN U5754 ( .A(n5480), .B(n5479), .Z(n5484) );
  NANDN U5755 ( .A(n5482), .B(n5481), .Z(n5483) );
  AND U5756 ( .A(n5484), .B(n5483), .Z(n5594) );
  XOR U5757 ( .A(n5595), .B(n5594), .Z(n5708) );
  NANDN U5758 ( .A(n5486), .B(n5485), .Z(n5490) );
  NANDN U5759 ( .A(n5488), .B(n5487), .Z(n5489) );
  AND U5760 ( .A(n5490), .B(n5489), .Z(n5706) );
  NANDN U5761 ( .A(n5492), .B(n5491), .Z(n5496) );
  NANDN U5762 ( .A(n5494), .B(n5493), .Z(n5495) );
  AND U5763 ( .A(n5496), .B(n5495), .Z(n5589) );
  NANDN U5764 ( .A(n5498), .B(n5497), .Z(n5502) );
  OR U5765 ( .A(n5500), .B(n5499), .Z(n5501) );
  AND U5766 ( .A(n5502), .B(n5501), .Z(n5587) );
  NANDN U5767 ( .A(n5504), .B(n5503), .Z(n5508) );
  NANDN U5768 ( .A(n5506), .B(n5505), .Z(n5507) );
  AND U5769 ( .A(n5508), .B(n5507), .Z(n5653) );
  NANDN U5770 ( .A(n5510), .B(n5509), .Z(n5514) );
  NANDN U5771 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U5772 ( .A(n5514), .B(n5513), .Z(n5652) );
  XNOR U5773 ( .A(n5653), .B(n5652), .Z(n5654) );
  NAND U5774 ( .A(b[0]), .B(a[52]), .Z(n5515) );
  XNOR U5775 ( .A(b[1]), .B(n5515), .Z(n5517) );
  NANDN U5776 ( .A(b[0]), .B(a[51]), .Z(n5516) );
  NAND U5777 ( .A(n5517), .B(n5516), .Z(n5601) );
  NANDN U5778 ( .A(n19394), .B(n5518), .Z(n5520) );
  XOR U5779 ( .A(b[29]), .B(a[24]), .Z(n5679) );
  NANDN U5780 ( .A(n19395), .B(n5679), .Z(n5519) );
  AND U5781 ( .A(n5520), .B(n5519), .Z(n5599) );
  AND U5782 ( .A(b[31]), .B(a[20]), .Z(n5598) );
  XNOR U5783 ( .A(n5599), .B(n5598), .Z(n5600) );
  XNOR U5784 ( .A(n5601), .B(n5600), .Z(n5640) );
  NANDN U5785 ( .A(n19005), .B(n5521), .Z(n5523) );
  XOR U5786 ( .A(b[23]), .B(a[30]), .Z(n5682) );
  NANDN U5787 ( .A(n19055), .B(n5682), .Z(n5522) );
  AND U5788 ( .A(n5523), .B(n5522), .Z(n5673) );
  NANDN U5789 ( .A(n17362), .B(n5524), .Z(n5526) );
  XOR U5790 ( .A(b[7]), .B(a[46]), .Z(n5685) );
  NANDN U5791 ( .A(n17522), .B(n5685), .Z(n5525) );
  AND U5792 ( .A(n5526), .B(n5525), .Z(n5671) );
  NANDN U5793 ( .A(n19116), .B(n5527), .Z(n5529) );
  XOR U5794 ( .A(b[25]), .B(a[28]), .Z(n5688) );
  NANDN U5795 ( .A(n19179), .B(n5688), .Z(n5528) );
  NAND U5796 ( .A(n5529), .B(n5528), .Z(n5670) );
  XNOR U5797 ( .A(n5671), .B(n5670), .Z(n5672) );
  XOR U5798 ( .A(n5673), .B(n5672), .Z(n5641) );
  XNOR U5799 ( .A(n5640), .B(n5641), .Z(n5642) );
  NANDN U5800 ( .A(n18113), .B(n5530), .Z(n5532) );
  XOR U5801 ( .A(b[13]), .B(a[40]), .Z(n5691) );
  NANDN U5802 ( .A(n18229), .B(n5691), .Z(n5531) );
  AND U5803 ( .A(n5532), .B(n5531), .Z(n5635) );
  NANDN U5804 ( .A(n17888), .B(n5533), .Z(n5535) );
  XOR U5805 ( .A(b[11]), .B(a[42]), .Z(n5694) );
  NANDN U5806 ( .A(n18025), .B(n5694), .Z(n5534) );
  NAND U5807 ( .A(n5535), .B(n5534), .Z(n5634) );
  XNOR U5808 ( .A(n5635), .B(n5634), .Z(n5636) );
  NANDN U5809 ( .A(n18487), .B(n5536), .Z(n5538) );
  XOR U5810 ( .A(b[15]), .B(a[38]), .Z(n5697) );
  NANDN U5811 ( .A(n18311), .B(n5697), .Z(n5537) );
  AND U5812 ( .A(n5538), .B(n5537), .Z(n5631) );
  NANDN U5813 ( .A(n18853), .B(n5539), .Z(n5541) );
  XOR U5814 ( .A(b[21]), .B(a[32]), .Z(n5700) );
  NANDN U5815 ( .A(n18926), .B(n5700), .Z(n5540) );
  AND U5816 ( .A(n5541), .B(n5540), .Z(n5629) );
  NANDN U5817 ( .A(n17613), .B(n5542), .Z(n5544) );
  XOR U5818 ( .A(b[9]), .B(a[44]), .Z(n5703) );
  NANDN U5819 ( .A(n17739), .B(n5703), .Z(n5543) );
  NAND U5820 ( .A(n5544), .B(n5543), .Z(n5628) );
  XNOR U5821 ( .A(n5629), .B(n5628), .Z(n5630) );
  XOR U5822 ( .A(n5631), .B(n5630), .Z(n5637) );
  XOR U5823 ( .A(n5636), .B(n5637), .Z(n5643) );
  XOR U5824 ( .A(n5642), .B(n5643), .Z(n5655) );
  XNOR U5825 ( .A(n5654), .B(n5655), .Z(n5586) );
  XNOR U5826 ( .A(n5587), .B(n5586), .Z(n5588) );
  XOR U5827 ( .A(n5589), .B(n5588), .Z(n5707) );
  XOR U5828 ( .A(n5706), .B(n5707), .Z(n5709) );
  XOR U5829 ( .A(n5708), .B(n5709), .Z(n5583) );
  NANDN U5830 ( .A(n5546), .B(n5545), .Z(n5550) );
  NAND U5831 ( .A(n5548), .B(n5547), .Z(n5549) );
  AND U5832 ( .A(n5550), .B(n5549), .Z(n5581) );
  NANDN U5833 ( .A(n5552), .B(n5551), .Z(n5556) );
  NANDN U5834 ( .A(n5554), .B(n5553), .Z(n5555) );
  AND U5835 ( .A(n5556), .B(n5555), .Z(n5580) );
  XNOR U5836 ( .A(n5581), .B(n5580), .Z(n5582) );
  XNOR U5837 ( .A(n5583), .B(n5582), .Z(n5574) );
  NANDN U5838 ( .A(n5558), .B(n5557), .Z(n5562) );
  OR U5839 ( .A(n5560), .B(n5559), .Z(n5561) );
  NAND U5840 ( .A(n5562), .B(n5561), .Z(n5575) );
  XNOR U5841 ( .A(n5574), .B(n5575), .Z(n5576) );
  XNOR U5842 ( .A(n5577), .B(n5576), .Z(n5568) );
  XNOR U5843 ( .A(n5569), .B(n5568), .Z(n5570) );
  XNOR U5844 ( .A(n5571), .B(n5570), .Z(n5712) );
  XNOR U5845 ( .A(sreg[148]), .B(n5712), .Z(n5714) );
  NANDN U5846 ( .A(sreg[147]), .B(n5563), .Z(n5567) );
  NAND U5847 ( .A(n5565), .B(n5564), .Z(n5566) );
  NAND U5848 ( .A(n5567), .B(n5566), .Z(n5713) );
  XNOR U5849 ( .A(n5714), .B(n5713), .Z(c[148]) );
  NANDN U5850 ( .A(n5569), .B(n5568), .Z(n5573) );
  NANDN U5851 ( .A(n5571), .B(n5570), .Z(n5572) );
  AND U5852 ( .A(n5573), .B(n5572), .Z(n5720) );
  NANDN U5853 ( .A(n5575), .B(n5574), .Z(n5579) );
  NANDN U5854 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U5855 ( .A(n5579), .B(n5578), .Z(n5718) );
  NANDN U5856 ( .A(n5581), .B(n5580), .Z(n5585) );
  NANDN U5857 ( .A(n5583), .B(n5582), .Z(n5584) );
  AND U5858 ( .A(n5585), .B(n5584), .Z(n5726) );
  NANDN U5859 ( .A(n5587), .B(n5586), .Z(n5591) );
  NANDN U5860 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U5861 ( .A(n5591), .B(n5590), .Z(n5730) );
  NANDN U5862 ( .A(n5593), .B(n5592), .Z(n5597) );
  NAND U5863 ( .A(n5595), .B(n5594), .Z(n5596) );
  AND U5864 ( .A(n5597), .B(n5596), .Z(n5729) );
  XNOR U5865 ( .A(n5730), .B(n5729), .Z(n5732) );
  NANDN U5866 ( .A(n5599), .B(n5598), .Z(n5603) );
  NANDN U5867 ( .A(n5601), .B(n5600), .Z(n5602) );
  AND U5868 ( .A(n5603), .B(n5602), .Z(n5809) );
  NANDN U5869 ( .A(n19237), .B(n5604), .Z(n5606) );
  XOR U5870 ( .A(b[27]), .B(a[27]), .Z(n5753) );
  NANDN U5871 ( .A(n19277), .B(n5753), .Z(n5605) );
  AND U5872 ( .A(n5606), .B(n5605), .Z(n5816) );
  NANDN U5873 ( .A(n17072), .B(n5607), .Z(n5609) );
  XOR U5874 ( .A(b[5]), .B(a[49]), .Z(n5756) );
  NANDN U5875 ( .A(n17223), .B(n5756), .Z(n5608) );
  AND U5876 ( .A(n5609), .B(n5608), .Z(n5814) );
  NANDN U5877 ( .A(n18673), .B(n5610), .Z(n5612) );
  XOR U5878 ( .A(b[19]), .B(a[35]), .Z(n5759) );
  NANDN U5879 ( .A(n18758), .B(n5759), .Z(n5611) );
  NAND U5880 ( .A(n5612), .B(n5611), .Z(n5813) );
  XNOR U5881 ( .A(n5814), .B(n5813), .Z(n5815) );
  XNOR U5882 ( .A(n5816), .B(n5815), .Z(n5807) );
  NANDN U5883 ( .A(n19425), .B(n5613), .Z(n5615) );
  XOR U5884 ( .A(b[31]), .B(a[23]), .Z(n5762) );
  NANDN U5885 ( .A(n19426), .B(n5762), .Z(n5614) );
  AND U5886 ( .A(n5615), .B(n5614), .Z(n5774) );
  NANDN U5887 ( .A(n17067), .B(n5616), .Z(n5618) );
  XOR U5888 ( .A(b[3]), .B(a[51]), .Z(n5765) );
  NANDN U5889 ( .A(n17068), .B(n5765), .Z(n5617) );
  AND U5890 ( .A(n5618), .B(n5617), .Z(n5772) );
  NANDN U5891 ( .A(n18514), .B(n5619), .Z(n5621) );
  XOR U5892 ( .A(b[17]), .B(a[37]), .Z(n5768) );
  NANDN U5893 ( .A(n18585), .B(n5768), .Z(n5620) );
  NAND U5894 ( .A(n5621), .B(n5620), .Z(n5771) );
  XNOR U5895 ( .A(n5772), .B(n5771), .Z(n5773) );
  XOR U5896 ( .A(n5774), .B(n5773), .Z(n5808) );
  XOR U5897 ( .A(n5807), .B(n5808), .Z(n5810) );
  XOR U5898 ( .A(n5809), .B(n5810), .Z(n5742) );
  NANDN U5899 ( .A(n5623), .B(n5622), .Z(n5627) );
  NANDN U5900 ( .A(n5625), .B(n5624), .Z(n5626) );
  AND U5901 ( .A(n5627), .B(n5626), .Z(n5795) );
  NANDN U5902 ( .A(n5629), .B(n5628), .Z(n5633) );
  NANDN U5903 ( .A(n5631), .B(n5630), .Z(n5632) );
  NAND U5904 ( .A(n5633), .B(n5632), .Z(n5796) );
  XNOR U5905 ( .A(n5795), .B(n5796), .Z(n5797) );
  NANDN U5906 ( .A(n5635), .B(n5634), .Z(n5639) );
  NANDN U5907 ( .A(n5637), .B(n5636), .Z(n5638) );
  NAND U5908 ( .A(n5639), .B(n5638), .Z(n5798) );
  XNOR U5909 ( .A(n5797), .B(n5798), .Z(n5741) );
  XNOR U5910 ( .A(n5742), .B(n5741), .Z(n5744) );
  NANDN U5911 ( .A(n5641), .B(n5640), .Z(n5645) );
  NANDN U5912 ( .A(n5643), .B(n5642), .Z(n5644) );
  AND U5913 ( .A(n5645), .B(n5644), .Z(n5743) );
  XOR U5914 ( .A(n5744), .B(n5743), .Z(n5858) );
  NANDN U5915 ( .A(n5647), .B(n5646), .Z(n5651) );
  NANDN U5916 ( .A(n5649), .B(n5648), .Z(n5650) );
  AND U5917 ( .A(n5651), .B(n5650), .Z(n5855) );
  NANDN U5918 ( .A(n5653), .B(n5652), .Z(n5657) );
  NANDN U5919 ( .A(n5655), .B(n5654), .Z(n5656) );
  AND U5920 ( .A(n5657), .B(n5656), .Z(n5738) );
  NANDN U5921 ( .A(n5659), .B(n5658), .Z(n5663) );
  OR U5922 ( .A(n5661), .B(n5660), .Z(n5662) );
  AND U5923 ( .A(n5663), .B(n5662), .Z(n5736) );
  NANDN U5924 ( .A(n5665), .B(n5664), .Z(n5669) );
  NANDN U5925 ( .A(n5667), .B(n5666), .Z(n5668) );
  AND U5926 ( .A(n5669), .B(n5668), .Z(n5802) );
  NANDN U5927 ( .A(n5671), .B(n5670), .Z(n5675) );
  NANDN U5928 ( .A(n5673), .B(n5672), .Z(n5674) );
  NAND U5929 ( .A(n5675), .B(n5674), .Z(n5801) );
  XNOR U5930 ( .A(n5802), .B(n5801), .Z(n5803) );
  NAND U5931 ( .A(b[0]), .B(a[53]), .Z(n5676) );
  XNOR U5932 ( .A(b[1]), .B(n5676), .Z(n5678) );
  NANDN U5933 ( .A(b[0]), .B(a[52]), .Z(n5677) );
  NAND U5934 ( .A(n5678), .B(n5677), .Z(n5750) );
  NANDN U5935 ( .A(n19394), .B(n5679), .Z(n5681) );
  XOR U5936 ( .A(b[29]), .B(a[25]), .Z(n5828) );
  NANDN U5937 ( .A(n19395), .B(n5828), .Z(n5680) );
  AND U5938 ( .A(n5681), .B(n5680), .Z(n5748) );
  AND U5939 ( .A(b[31]), .B(a[21]), .Z(n5747) );
  XNOR U5940 ( .A(n5748), .B(n5747), .Z(n5749) );
  XNOR U5941 ( .A(n5750), .B(n5749), .Z(n5789) );
  NANDN U5942 ( .A(n19005), .B(n5682), .Z(n5684) );
  XOR U5943 ( .A(b[23]), .B(a[31]), .Z(n5831) );
  NANDN U5944 ( .A(n19055), .B(n5831), .Z(n5683) );
  AND U5945 ( .A(n5684), .B(n5683), .Z(n5822) );
  NANDN U5946 ( .A(n17362), .B(n5685), .Z(n5687) );
  XOR U5947 ( .A(b[7]), .B(a[47]), .Z(n5834) );
  NANDN U5948 ( .A(n17522), .B(n5834), .Z(n5686) );
  AND U5949 ( .A(n5687), .B(n5686), .Z(n5820) );
  NANDN U5950 ( .A(n19116), .B(n5688), .Z(n5690) );
  XOR U5951 ( .A(b[25]), .B(a[29]), .Z(n5837) );
  NANDN U5952 ( .A(n19179), .B(n5837), .Z(n5689) );
  NAND U5953 ( .A(n5690), .B(n5689), .Z(n5819) );
  XNOR U5954 ( .A(n5820), .B(n5819), .Z(n5821) );
  XOR U5955 ( .A(n5822), .B(n5821), .Z(n5790) );
  XNOR U5956 ( .A(n5789), .B(n5790), .Z(n5791) );
  NANDN U5957 ( .A(n18113), .B(n5691), .Z(n5693) );
  XOR U5958 ( .A(b[13]), .B(a[41]), .Z(n5840) );
  NANDN U5959 ( .A(n18229), .B(n5840), .Z(n5692) );
  AND U5960 ( .A(n5693), .B(n5692), .Z(n5784) );
  NANDN U5961 ( .A(n17888), .B(n5694), .Z(n5696) );
  XOR U5962 ( .A(b[11]), .B(a[43]), .Z(n5843) );
  NANDN U5963 ( .A(n18025), .B(n5843), .Z(n5695) );
  NAND U5964 ( .A(n5696), .B(n5695), .Z(n5783) );
  XNOR U5965 ( .A(n5784), .B(n5783), .Z(n5785) );
  NANDN U5966 ( .A(n18487), .B(n5697), .Z(n5699) );
  XOR U5967 ( .A(b[15]), .B(a[39]), .Z(n5846) );
  NANDN U5968 ( .A(n18311), .B(n5846), .Z(n5698) );
  AND U5969 ( .A(n5699), .B(n5698), .Z(n5780) );
  NANDN U5970 ( .A(n18853), .B(n5700), .Z(n5702) );
  XOR U5971 ( .A(b[21]), .B(a[33]), .Z(n5849) );
  NANDN U5972 ( .A(n18926), .B(n5849), .Z(n5701) );
  AND U5973 ( .A(n5702), .B(n5701), .Z(n5778) );
  NANDN U5974 ( .A(n17613), .B(n5703), .Z(n5705) );
  XOR U5975 ( .A(b[9]), .B(a[45]), .Z(n5852) );
  NANDN U5976 ( .A(n17739), .B(n5852), .Z(n5704) );
  NAND U5977 ( .A(n5705), .B(n5704), .Z(n5777) );
  XNOR U5978 ( .A(n5778), .B(n5777), .Z(n5779) );
  XOR U5979 ( .A(n5780), .B(n5779), .Z(n5786) );
  XOR U5980 ( .A(n5785), .B(n5786), .Z(n5792) );
  XOR U5981 ( .A(n5791), .B(n5792), .Z(n5804) );
  XNOR U5982 ( .A(n5803), .B(n5804), .Z(n5735) );
  XNOR U5983 ( .A(n5736), .B(n5735), .Z(n5737) );
  XOR U5984 ( .A(n5738), .B(n5737), .Z(n5856) );
  XNOR U5985 ( .A(n5855), .B(n5856), .Z(n5857) );
  XNOR U5986 ( .A(n5858), .B(n5857), .Z(n5731) );
  XOR U5987 ( .A(n5732), .B(n5731), .Z(n5724) );
  NANDN U5988 ( .A(n5707), .B(n5706), .Z(n5711) );
  OR U5989 ( .A(n5709), .B(n5708), .Z(n5710) );
  AND U5990 ( .A(n5711), .B(n5710), .Z(n5723) );
  XNOR U5991 ( .A(n5724), .B(n5723), .Z(n5725) );
  XNOR U5992 ( .A(n5726), .B(n5725), .Z(n5717) );
  XNOR U5993 ( .A(n5718), .B(n5717), .Z(n5719) );
  XNOR U5994 ( .A(n5720), .B(n5719), .Z(n5861) );
  XNOR U5995 ( .A(sreg[149]), .B(n5861), .Z(n5863) );
  NANDN U5996 ( .A(sreg[148]), .B(n5712), .Z(n5716) );
  NAND U5997 ( .A(n5714), .B(n5713), .Z(n5715) );
  NAND U5998 ( .A(n5716), .B(n5715), .Z(n5862) );
  XNOR U5999 ( .A(n5863), .B(n5862), .Z(c[149]) );
  NANDN U6000 ( .A(n5718), .B(n5717), .Z(n5722) );
  NANDN U6001 ( .A(n5720), .B(n5719), .Z(n5721) );
  AND U6002 ( .A(n5722), .B(n5721), .Z(n5869) );
  NANDN U6003 ( .A(n5724), .B(n5723), .Z(n5728) );
  NANDN U6004 ( .A(n5726), .B(n5725), .Z(n5727) );
  AND U6005 ( .A(n5728), .B(n5727), .Z(n5867) );
  NANDN U6006 ( .A(n5730), .B(n5729), .Z(n5734) );
  NAND U6007 ( .A(n5732), .B(n5731), .Z(n5733) );
  AND U6008 ( .A(n5734), .B(n5733), .Z(n5874) );
  NANDN U6009 ( .A(n5736), .B(n5735), .Z(n5740) );
  NANDN U6010 ( .A(n5738), .B(n5737), .Z(n5739) );
  AND U6011 ( .A(n5740), .B(n5739), .Z(n5879) );
  NANDN U6012 ( .A(n5742), .B(n5741), .Z(n5746) );
  NAND U6013 ( .A(n5744), .B(n5743), .Z(n5745) );
  AND U6014 ( .A(n5746), .B(n5745), .Z(n5878) );
  XNOR U6015 ( .A(n5879), .B(n5878), .Z(n5881) );
  NANDN U6016 ( .A(n5748), .B(n5747), .Z(n5752) );
  NANDN U6017 ( .A(n5750), .B(n5749), .Z(n5751) );
  AND U6018 ( .A(n5752), .B(n5751), .Z(n5958) );
  NANDN U6019 ( .A(n19237), .B(n5753), .Z(n5755) );
  XOR U6020 ( .A(b[27]), .B(a[28]), .Z(n5902) );
  NANDN U6021 ( .A(n19277), .B(n5902), .Z(n5754) );
  AND U6022 ( .A(n5755), .B(n5754), .Z(n5965) );
  NANDN U6023 ( .A(n17072), .B(n5756), .Z(n5758) );
  XOR U6024 ( .A(b[5]), .B(a[50]), .Z(n5905) );
  NANDN U6025 ( .A(n17223), .B(n5905), .Z(n5757) );
  AND U6026 ( .A(n5758), .B(n5757), .Z(n5963) );
  NANDN U6027 ( .A(n18673), .B(n5759), .Z(n5761) );
  XOR U6028 ( .A(b[19]), .B(a[36]), .Z(n5908) );
  NANDN U6029 ( .A(n18758), .B(n5908), .Z(n5760) );
  NAND U6030 ( .A(n5761), .B(n5760), .Z(n5962) );
  XNOR U6031 ( .A(n5963), .B(n5962), .Z(n5964) );
  XNOR U6032 ( .A(n5965), .B(n5964), .Z(n5956) );
  NANDN U6033 ( .A(n19425), .B(n5762), .Z(n5764) );
  XOR U6034 ( .A(b[31]), .B(a[24]), .Z(n5911) );
  NANDN U6035 ( .A(n19426), .B(n5911), .Z(n5763) );
  AND U6036 ( .A(n5764), .B(n5763), .Z(n5923) );
  NANDN U6037 ( .A(n17067), .B(n5765), .Z(n5767) );
  XOR U6038 ( .A(b[3]), .B(a[52]), .Z(n5914) );
  NANDN U6039 ( .A(n17068), .B(n5914), .Z(n5766) );
  AND U6040 ( .A(n5767), .B(n5766), .Z(n5921) );
  NANDN U6041 ( .A(n18514), .B(n5768), .Z(n5770) );
  XOR U6042 ( .A(b[17]), .B(a[38]), .Z(n5917) );
  NANDN U6043 ( .A(n18585), .B(n5917), .Z(n5769) );
  NAND U6044 ( .A(n5770), .B(n5769), .Z(n5920) );
  XNOR U6045 ( .A(n5921), .B(n5920), .Z(n5922) );
  XOR U6046 ( .A(n5923), .B(n5922), .Z(n5957) );
  XOR U6047 ( .A(n5956), .B(n5957), .Z(n5959) );
  XOR U6048 ( .A(n5958), .B(n5959), .Z(n5891) );
  NANDN U6049 ( .A(n5772), .B(n5771), .Z(n5776) );
  NANDN U6050 ( .A(n5774), .B(n5773), .Z(n5775) );
  AND U6051 ( .A(n5776), .B(n5775), .Z(n5944) );
  NANDN U6052 ( .A(n5778), .B(n5777), .Z(n5782) );
  NANDN U6053 ( .A(n5780), .B(n5779), .Z(n5781) );
  NAND U6054 ( .A(n5782), .B(n5781), .Z(n5945) );
  XNOR U6055 ( .A(n5944), .B(n5945), .Z(n5946) );
  NANDN U6056 ( .A(n5784), .B(n5783), .Z(n5788) );
  NANDN U6057 ( .A(n5786), .B(n5785), .Z(n5787) );
  NAND U6058 ( .A(n5788), .B(n5787), .Z(n5947) );
  XNOR U6059 ( .A(n5946), .B(n5947), .Z(n5890) );
  XNOR U6060 ( .A(n5891), .B(n5890), .Z(n5893) );
  NANDN U6061 ( .A(n5790), .B(n5789), .Z(n5794) );
  NANDN U6062 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U6063 ( .A(n5794), .B(n5793), .Z(n5892) );
  XOR U6064 ( .A(n5893), .B(n5892), .Z(n6007) );
  NANDN U6065 ( .A(n5796), .B(n5795), .Z(n5800) );
  NANDN U6066 ( .A(n5798), .B(n5797), .Z(n5799) );
  AND U6067 ( .A(n5800), .B(n5799), .Z(n6004) );
  NANDN U6068 ( .A(n5802), .B(n5801), .Z(n5806) );
  NANDN U6069 ( .A(n5804), .B(n5803), .Z(n5805) );
  AND U6070 ( .A(n5806), .B(n5805), .Z(n5887) );
  NANDN U6071 ( .A(n5808), .B(n5807), .Z(n5812) );
  OR U6072 ( .A(n5810), .B(n5809), .Z(n5811) );
  AND U6073 ( .A(n5812), .B(n5811), .Z(n5885) );
  NANDN U6074 ( .A(n5814), .B(n5813), .Z(n5818) );
  NANDN U6075 ( .A(n5816), .B(n5815), .Z(n5817) );
  AND U6076 ( .A(n5818), .B(n5817), .Z(n5951) );
  NANDN U6077 ( .A(n5820), .B(n5819), .Z(n5824) );
  NANDN U6078 ( .A(n5822), .B(n5821), .Z(n5823) );
  NAND U6079 ( .A(n5824), .B(n5823), .Z(n5950) );
  XNOR U6080 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U6081 ( .A(b[0]), .B(a[54]), .Z(n5825) );
  XNOR U6082 ( .A(b[1]), .B(n5825), .Z(n5827) );
  NANDN U6083 ( .A(b[0]), .B(a[53]), .Z(n5826) );
  NAND U6084 ( .A(n5827), .B(n5826), .Z(n5899) );
  NANDN U6085 ( .A(n19394), .B(n5828), .Z(n5830) );
  XOR U6086 ( .A(b[29]), .B(a[26]), .Z(n5977) );
  NANDN U6087 ( .A(n19395), .B(n5977), .Z(n5829) );
  AND U6088 ( .A(n5830), .B(n5829), .Z(n5897) );
  AND U6089 ( .A(b[31]), .B(a[22]), .Z(n5896) );
  XNOR U6090 ( .A(n5897), .B(n5896), .Z(n5898) );
  XNOR U6091 ( .A(n5899), .B(n5898), .Z(n5938) );
  NANDN U6092 ( .A(n19005), .B(n5831), .Z(n5833) );
  XOR U6093 ( .A(b[23]), .B(a[32]), .Z(n5980) );
  NANDN U6094 ( .A(n19055), .B(n5980), .Z(n5832) );
  AND U6095 ( .A(n5833), .B(n5832), .Z(n5971) );
  NANDN U6096 ( .A(n17362), .B(n5834), .Z(n5836) );
  XOR U6097 ( .A(b[7]), .B(a[48]), .Z(n5983) );
  NANDN U6098 ( .A(n17522), .B(n5983), .Z(n5835) );
  AND U6099 ( .A(n5836), .B(n5835), .Z(n5969) );
  NANDN U6100 ( .A(n19116), .B(n5837), .Z(n5839) );
  XOR U6101 ( .A(b[25]), .B(a[30]), .Z(n5986) );
  NANDN U6102 ( .A(n19179), .B(n5986), .Z(n5838) );
  NAND U6103 ( .A(n5839), .B(n5838), .Z(n5968) );
  XNOR U6104 ( .A(n5969), .B(n5968), .Z(n5970) );
  XOR U6105 ( .A(n5971), .B(n5970), .Z(n5939) );
  XNOR U6106 ( .A(n5938), .B(n5939), .Z(n5940) );
  NANDN U6107 ( .A(n18113), .B(n5840), .Z(n5842) );
  XOR U6108 ( .A(b[13]), .B(a[42]), .Z(n5989) );
  NANDN U6109 ( .A(n18229), .B(n5989), .Z(n5841) );
  AND U6110 ( .A(n5842), .B(n5841), .Z(n5933) );
  NANDN U6111 ( .A(n17888), .B(n5843), .Z(n5845) );
  XOR U6112 ( .A(b[11]), .B(a[44]), .Z(n5992) );
  NANDN U6113 ( .A(n18025), .B(n5992), .Z(n5844) );
  NAND U6114 ( .A(n5845), .B(n5844), .Z(n5932) );
  XNOR U6115 ( .A(n5933), .B(n5932), .Z(n5934) );
  NANDN U6116 ( .A(n18487), .B(n5846), .Z(n5848) );
  XOR U6117 ( .A(b[15]), .B(a[40]), .Z(n5995) );
  NANDN U6118 ( .A(n18311), .B(n5995), .Z(n5847) );
  AND U6119 ( .A(n5848), .B(n5847), .Z(n5929) );
  NANDN U6120 ( .A(n18853), .B(n5849), .Z(n5851) );
  XOR U6121 ( .A(b[21]), .B(a[34]), .Z(n5998) );
  NANDN U6122 ( .A(n18926), .B(n5998), .Z(n5850) );
  AND U6123 ( .A(n5851), .B(n5850), .Z(n5927) );
  NANDN U6124 ( .A(n17613), .B(n5852), .Z(n5854) );
  XOR U6125 ( .A(b[9]), .B(a[46]), .Z(n6001) );
  NANDN U6126 ( .A(n17739), .B(n6001), .Z(n5853) );
  NAND U6127 ( .A(n5854), .B(n5853), .Z(n5926) );
  XNOR U6128 ( .A(n5927), .B(n5926), .Z(n5928) );
  XOR U6129 ( .A(n5929), .B(n5928), .Z(n5935) );
  XOR U6130 ( .A(n5934), .B(n5935), .Z(n5941) );
  XOR U6131 ( .A(n5940), .B(n5941), .Z(n5953) );
  XNOR U6132 ( .A(n5952), .B(n5953), .Z(n5884) );
  XNOR U6133 ( .A(n5885), .B(n5884), .Z(n5886) );
  XOR U6134 ( .A(n5887), .B(n5886), .Z(n6005) );
  XNOR U6135 ( .A(n6004), .B(n6005), .Z(n6006) );
  XNOR U6136 ( .A(n6007), .B(n6006), .Z(n5880) );
  XOR U6137 ( .A(n5881), .B(n5880), .Z(n5873) );
  NANDN U6138 ( .A(n5856), .B(n5855), .Z(n5860) );
  NANDN U6139 ( .A(n5858), .B(n5857), .Z(n5859) );
  AND U6140 ( .A(n5860), .B(n5859), .Z(n5872) );
  XOR U6141 ( .A(n5873), .B(n5872), .Z(n5875) );
  XNOR U6142 ( .A(n5874), .B(n5875), .Z(n5866) );
  XNOR U6143 ( .A(n5867), .B(n5866), .Z(n5868) );
  XNOR U6144 ( .A(n5869), .B(n5868), .Z(n6010) );
  XNOR U6145 ( .A(sreg[150]), .B(n6010), .Z(n6012) );
  NANDN U6146 ( .A(sreg[149]), .B(n5861), .Z(n5865) );
  NAND U6147 ( .A(n5863), .B(n5862), .Z(n5864) );
  NAND U6148 ( .A(n5865), .B(n5864), .Z(n6011) );
  XNOR U6149 ( .A(n6012), .B(n6011), .Z(c[150]) );
  NANDN U6150 ( .A(n5867), .B(n5866), .Z(n5871) );
  NANDN U6151 ( .A(n5869), .B(n5868), .Z(n5870) );
  AND U6152 ( .A(n5871), .B(n5870), .Z(n6018) );
  NANDN U6153 ( .A(n5873), .B(n5872), .Z(n5877) );
  NANDN U6154 ( .A(n5875), .B(n5874), .Z(n5876) );
  AND U6155 ( .A(n5877), .B(n5876), .Z(n6016) );
  NANDN U6156 ( .A(n5879), .B(n5878), .Z(n5883) );
  NAND U6157 ( .A(n5881), .B(n5880), .Z(n5882) );
  AND U6158 ( .A(n5883), .B(n5882), .Z(n6023) );
  NANDN U6159 ( .A(n5885), .B(n5884), .Z(n5889) );
  NANDN U6160 ( .A(n5887), .B(n5886), .Z(n5888) );
  AND U6161 ( .A(n5889), .B(n5888), .Z(n6028) );
  NANDN U6162 ( .A(n5891), .B(n5890), .Z(n5895) );
  NAND U6163 ( .A(n5893), .B(n5892), .Z(n5894) );
  AND U6164 ( .A(n5895), .B(n5894), .Z(n6027) );
  XNOR U6165 ( .A(n6028), .B(n6027), .Z(n6030) );
  NANDN U6166 ( .A(n5897), .B(n5896), .Z(n5901) );
  NANDN U6167 ( .A(n5899), .B(n5898), .Z(n5900) );
  AND U6168 ( .A(n5901), .B(n5900), .Z(n6107) );
  NANDN U6169 ( .A(n19237), .B(n5902), .Z(n5904) );
  XOR U6170 ( .A(b[27]), .B(a[29]), .Z(n6051) );
  NANDN U6171 ( .A(n19277), .B(n6051), .Z(n5903) );
  AND U6172 ( .A(n5904), .B(n5903), .Z(n6114) );
  NANDN U6173 ( .A(n17072), .B(n5905), .Z(n5907) );
  XOR U6174 ( .A(b[5]), .B(a[51]), .Z(n6054) );
  NANDN U6175 ( .A(n17223), .B(n6054), .Z(n5906) );
  AND U6176 ( .A(n5907), .B(n5906), .Z(n6112) );
  NANDN U6177 ( .A(n18673), .B(n5908), .Z(n5910) );
  XOR U6178 ( .A(b[19]), .B(a[37]), .Z(n6057) );
  NANDN U6179 ( .A(n18758), .B(n6057), .Z(n5909) );
  NAND U6180 ( .A(n5910), .B(n5909), .Z(n6111) );
  XNOR U6181 ( .A(n6112), .B(n6111), .Z(n6113) );
  XNOR U6182 ( .A(n6114), .B(n6113), .Z(n6105) );
  NANDN U6183 ( .A(n19425), .B(n5911), .Z(n5913) );
  XOR U6184 ( .A(b[31]), .B(a[25]), .Z(n6060) );
  NANDN U6185 ( .A(n19426), .B(n6060), .Z(n5912) );
  AND U6186 ( .A(n5913), .B(n5912), .Z(n6072) );
  NANDN U6187 ( .A(n17067), .B(n5914), .Z(n5916) );
  XOR U6188 ( .A(b[3]), .B(a[53]), .Z(n6063) );
  NANDN U6189 ( .A(n17068), .B(n6063), .Z(n5915) );
  AND U6190 ( .A(n5916), .B(n5915), .Z(n6070) );
  NANDN U6191 ( .A(n18514), .B(n5917), .Z(n5919) );
  XOR U6192 ( .A(b[17]), .B(a[39]), .Z(n6066) );
  NANDN U6193 ( .A(n18585), .B(n6066), .Z(n5918) );
  NAND U6194 ( .A(n5919), .B(n5918), .Z(n6069) );
  XNOR U6195 ( .A(n6070), .B(n6069), .Z(n6071) );
  XOR U6196 ( .A(n6072), .B(n6071), .Z(n6106) );
  XOR U6197 ( .A(n6105), .B(n6106), .Z(n6108) );
  XOR U6198 ( .A(n6107), .B(n6108), .Z(n6040) );
  NANDN U6199 ( .A(n5921), .B(n5920), .Z(n5925) );
  NANDN U6200 ( .A(n5923), .B(n5922), .Z(n5924) );
  AND U6201 ( .A(n5925), .B(n5924), .Z(n6093) );
  NANDN U6202 ( .A(n5927), .B(n5926), .Z(n5931) );
  NANDN U6203 ( .A(n5929), .B(n5928), .Z(n5930) );
  NAND U6204 ( .A(n5931), .B(n5930), .Z(n6094) );
  XNOR U6205 ( .A(n6093), .B(n6094), .Z(n6095) );
  NANDN U6206 ( .A(n5933), .B(n5932), .Z(n5937) );
  NANDN U6207 ( .A(n5935), .B(n5934), .Z(n5936) );
  NAND U6208 ( .A(n5937), .B(n5936), .Z(n6096) );
  XNOR U6209 ( .A(n6095), .B(n6096), .Z(n6039) );
  XNOR U6210 ( .A(n6040), .B(n6039), .Z(n6042) );
  NANDN U6211 ( .A(n5939), .B(n5938), .Z(n5943) );
  NANDN U6212 ( .A(n5941), .B(n5940), .Z(n5942) );
  AND U6213 ( .A(n5943), .B(n5942), .Z(n6041) );
  XOR U6214 ( .A(n6042), .B(n6041), .Z(n6156) );
  NANDN U6215 ( .A(n5945), .B(n5944), .Z(n5949) );
  NANDN U6216 ( .A(n5947), .B(n5946), .Z(n5948) );
  AND U6217 ( .A(n5949), .B(n5948), .Z(n6153) );
  NANDN U6218 ( .A(n5951), .B(n5950), .Z(n5955) );
  NANDN U6219 ( .A(n5953), .B(n5952), .Z(n5954) );
  AND U6220 ( .A(n5955), .B(n5954), .Z(n6036) );
  NANDN U6221 ( .A(n5957), .B(n5956), .Z(n5961) );
  OR U6222 ( .A(n5959), .B(n5958), .Z(n5960) );
  AND U6223 ( .A(n5961), .B(n5960), .Z(n6034) );
  NANDN U6224 ( .A(n5963), .B(n5962), .Z(n5967) );
  NANDN U6225 ( .A(n5965), .B(n5964), .Z(n5966) );
  AND U6226 ( .A(n5967), .B(n5966), .Z(n6100) );
  NANDN U6227 ( .A(n5969), .B(n5968), .Z(n5973) );
  NANDN U6228 ( .A(n5971), .B(n5970), .Z(n5972) );
  NAND U6229 ( .A(n5973), .B(n5972), .Z(n6099) );
  XNOR U6230 ( .A(n6100), .B(n6099), .Z(n6101) );
  NAND U6231 ( .A(b[0]), .B(a[55]), .Z(n5974) );
  XNOR U6232 ( .A(b[1]), .B(n5974), .Z(n5976) );
  NANDN U6233 ( .A(b[0]), .B(a[54]), .Z(n5975) );
  NAND U6234 ( .A(n5976), .B(n5975), .Z(n6048) );
  NANDN U6235 ( .A(n19394), .B(n5977), .Z(n5979) );
  XOR U6236 ( .A(b[29]), .B(a[27]), .Z(n6126) );
  NANDN U6237 ( .A(n19395), .B(n6126), .Z(n5978) );
  AND U6238 ( .A(n5979), .B(n5978), .Z(n6046) );
  AND U6239 ( .A(b[31]), .B(a[23]), .Z(n6045) );
  XNOR U6240 ( .A(n6046), .B(n6045), .Z(n6047) );
  XNOR U6241 ( .A(n6048), .B(n6047), .Z(n6087) );
  NANDN U6242 ( .A(n19005), .B(n5980), .Z(n5982) );
  XOR U6243 ( .A(b[23]), .B(a[33]), .Z(n6129) );
  NANDN U6244 ( .A(n19055), .B(n6129), .Z(n5981) );
  AND U6245 ( .A(n5982), .B(n5981), .Z(n6120) );
  NANDN U6246 ( .A(n17362), .B(n5983), .Z(n5985) );
  XOR U6247 ( .A(b[7]), .B(a[49]), .Z(n6132) );
  NANDN U6248 ( .A(n17522), .B(n6132), .Z(n5984) );
  AND U6249 ( .A(n5985), .B(n5984), .Z(n6118) );
  NANDN U6250 ( .A(n19116), .B(n5986), .Z(n5988) );
  XOR U6251 ( .A(b[25]), .B(a[31]), .Z(n6135) );
  NANDN U6252 ( .A(n19179), .B(n6135), .Z(n5987) );
  NAND U6253 ( .A(n5988), .B(n5987), .Z(n6117) );
  XNOR U6254 ( .A(n6118), .B(n6117), .Z(n6119) );
  XOR U6255 ( .A(n6120), .B(n6119), .Z(n6088) );
  XNOR U6256 ( .A(n6087), .B(n6088), .Z(n6089) );
  NANDN U6257 ( .A(n18113), .B(n5989), .Z(n5991) );
  XOR U6258 ( .A(b[13]), .B(a[43]), .Z(n6138) );
  NANDN U6259 ( .A(n18229), .B(n6138), .Z(n5990) );
  AND U6260 ( .A(n5991), .B(n5990), .Z(n6082) );
  NANDN U6261 ( .A(n17888), .B(n5992), .Z(n5994) );
  XOR U6262 ( .A(b[11]), .B(a[45]), .Z(n6141) );
  NANDN U6263 ( .A(n18025), .B(n6141), .Z(n5993) );
  NAND U6264 ( .A(n5994), .B(n5993), .Z(n6081) );
  XNOR U6265 ( .A(n6082), .B(n6081), .Z(n6083) );
  NANDN U6266 ( .A(n18487), .B(n5995), .Z(n5997) );
  XOR U6267 ( .A(b[15]), .B(a[41]), .Z(n6144) );
  NANDN U6268 ( .A(n18311), .B(n6144), .Z(n5996) );
  AND U6269 ( .A(n5997), .B(n5996), .Z(n6078) );
  NANDN U6270 ( .A(n18853), .B(n5998), .Z(n6000) );
  XOR U6271 ( .A(b[21]), .B(a[35]), .Z(n6147) );
  NANDN U6272 ( .A(n18926), .B(n6147), .Z(n5999) );
  AND U6273 ( .A(n6000), .B(n5999), .Z(n6076) );
  NANDN U6274 ( .A(n17613), .B(n6001), .Z(n6003) );
  XOR U6275 ( .A(b[9]), .B(a[47]), .Z(n6150) );
  NANDN U6276 ( .A(n17739), .B(n6150), .Z(n6002) );
  NAND U6277 ( .A(n6003), .B(n6002), .Z(n6075) );
  XNOR U6278 ( .A(n6076), .B(n6075), .Z(n6077) );
  XOR U6279 ( .A(n6078), .B(n6077), .Z(n6084) );
  XOR U6280 ( .A(n6083), .B(n6084), .Z(n6090) );
  XOR U6281 ( .A(n6089), .B(n6090), .Z(n6102) );
  XNOR U6282 ( .A(n6101), .B(n6102), .Z(n6033) );
  XNOR U6283 ( .A(n6034), .B(n6033), .Z(n6035) );
  XOR U6284 ( .A(n6036), .B(n6035), .Z(n6154) );
  XNOR U6285 ( .A(n6153), .B(n6154), .Z(n6155) );
  XNOR U6286 ( .A(n6156), .B(n6155), .Z(n6029) );
  XOR U6287 ( .A(n6030), .B(n6029), .Z(n6022) );
  NANDN U6288 ( .A(n6005), .B(n6004), .Z(n6009) );
  NANDN U6289 ( .A(n6007), .B(n6006), .Z(n6008) );
  AND U6290 ( .A(n6009), .B(n6008), .Z(n6021) );
  XOR U6291 ( .A(n6022), .B(n6021), .Z(n6024) );
  XNOR U6292 ( .A(n6023), .B(n6024), .Z(n6015) );
  XNOR U6293 ( .A(n6016), .B(n6015), .Z(n6017) );
  XNOR U6294 ( .A(n6018), .B(n6017), .Z(n6159) );
  XNOR U6295 ( .A(sreg[151]), .B(n6159), .Z(n6161) );
  NANDN U6296 ( .A(sreg[150]), .B(n6010), .Z(n6014) );
  NAND U6297 ( .A(n6012), .B(n6011), .Z(n6013) );
  NAND U6298 ( .A(n6014), .B(n6013), .Z(n6160) );
  XNOR U6299 ( .A(n6161), .B(n6160), .Z(c[151]) );
  NANDN U6300 ( .A(n6016), .B(n6015), .Z(n6020) );
  NANDN U6301 ( .A(n6018), .B(n6017), .Z(n6019) );
  AND U6302 ( .A(n6020), .B(n6019), .Z(n6167) );
  NANDN U6303 ( .A(n6022), .B(n6021), .Z(n6026) );
  NANDN U6304 ( .A(n6024), .B(n6023), .Z(n6025) );
  AND U6305 ( .A(n6026), .B(n6025), .Z(n6165) );
  NANDN U6306 ( .A(n6028), .B(n6027), .Z(n6032) );
  NAND U6307 ( .A(n6030), .B(n6029), .Z(n6031) );
  AND U6308 ( .A(n6032), .B(n6031), .Z(n6172) );
  NANDN U6309 ( .A(n6034), .B(n6033), .Z(n6038) );
  NANDN U6310 ( .A(n6036), .B(n6035), .Z(n6037) );
  AND U6311 ( .A(n6038), .B(n6037), .Z(n6177) );
  NANDN U6312 ( .A(n6040), .B(n6039), .Z(n6044) );
  NAND U6313 ( .A(n6042), .B(n6041), .Z(n6043) );
  AND U6314 ( .A(n6044), .B(n6043), .Z(n6176) );
  XNOR U6315 ( .A(n6177), .B(n6176), .Z(n6179) );
  NANDN U6316 ( .A(n6046), .B(n6045), .Z(n6050) );
  NANDN U6317 ( .A(n6048), .B(n6047), .Z(n6049) );
  AND U6318 ( .A(n6050), .B(n6049), .Z(n6254) );
  NANDN U6319 ( .A(n19237), .B(n6051), .Z(n6053) );
  XOR U6320 ( .A(b[27]), .B(a[30]), .Z(n6200) );
  NANDN U6321 ( .A(n19277), .B(n6200), .Z(n6052) );
  AND U6322 ( .A(n6053), .B(n6052), .Z(n6261) );
  NANDN U6323 ( .A(n17072), .B(n6054), .Z(n6056) );
  XOR U6324 ( .A(b[5]), .B(a[52]), .Z(n6203) );
  NANDN U6325 ( .A(n17223), .B(n6203), .Z(n6055) );
  AND U6326 ( .A(n6056), .B(n6055), .Z(n6259) );
  NANDN U6327 ( .A(n18673), .B(n6057), .Z(n6059) );
  XOR U6328 ( .A(b[19]), .B(a[38]), .Z(n6206) );
  NANDN U6329 ( .A(n18758), .B(n6206), .Z(n6058) );
  NAND U6330 ( .A(n6059), .B(n6058), .Z(n6258) );
  XNOR U6331 ( .A(n6259), .B(n6258), .Z(n6260) );
  XNOR U6332 ( .A(n6261), .B(n6260), .Z(n6252) );
  NANDN U6333 ( .A(n19425), .B(n6060), .Z(n6062) );
  XOR U6334 ( .A(b[31]), .B(a[26]), .Z(n6209) );
  NANDN U6335 ( .A(n19426), .B(n6209), .Z(n6061) );
  AND U6336 ( .A(n6062), .B(n6061), .Z(n6221) );
  NANDN U6337 ( .A(n17067), .B(n6063), .Z(n6065) );
  XOR U6338 ( .A(b[3]), .B(a[54]), .Z(n6212) );
  NANDN U6339 ( .A(n17068), .B(n6212), .Z(n6064) );
  AND U6340 ( .A(n6065), .B(n6064), .Z(n6219) );
  NANDN U6341 ( .A(n18514), .B(n6066), .Z(n6068) );
  XOR U6342 ( .A(b[17]), .B(a[40]), .Z(n6215) );
  NANDN U6343 ( .A(n18585), .B(n6215), .Z(n6067) );
  NAND U6344 ( .A(n6068), .B(n6067), .Z(n6218) );
  XNOR U6345 ( .A(n6219), .B(n6218), .Z(n6220) );
  XOR U6346 ( .A(n6221), .B(n6220), .Z(n6253) );
  XOR U6347 ( .A(n6252), .B(n6253), .Z(n6255) );
  XOR U6348 ( .A(n6254), .B(n6255), .Z(n6189) );
  NANDN U6349 ( .A(n6070), .B(n6069), .Z(n6074) );
  NANDN U6350 ( .A(n6072), .B(n6071), .Z(n6073) );
  AND U6351 ( .A(n6074), .B(n6073), .Z(n6242) );
  NANDN U6352 ( .A(n6076), .B(n6075), .Z(n6080) );
  NANDN U6353 ( .A(n6078), .B(n6077), .Z(n6079) );
  NAND U6354 ( .A(n6080), .B(n6079), .Z(n6243) );
  XNOR U6355 ( .A(n6242), .B(n6243), .Z(n6244) );
  NANDN U6356 ( .A(n6082), .B(n6081), .Z(n6086) );
  NANDN U6357 ( .A(n6084), .B(n6083), .Z(n6085) );
  NAND U6358 ( .A(n6086), .B(n6085), .Z(n6245) );
  XNOR U6359 ( .A(n6244), .B(n6245), .Z(n6188) );
  XNOR U6360 ( .A(n6189), .B(n6188), .Z(n6191) );
  NANDN U6361 ( .A(n6088), .B(n6087), .Z(n6092) );
  NANDN U6362 ( .A(n6090), .B(n6089), .Z(n6091) );
  AND U6363 ( .A(n6092), .B(n6091), .Z(n6190) );
  XOR U6364 ( .A(n6191), .B(n6190), .Z(n6303) );
  NANDN U6365 ( .A(n6094), .B(n6093), .Z(n6098) );
  NANDN U6366 ( .A(n6096), .B(n6095), .Z(n6097) );
  AND U6367 ( .A(n6098), .B(n6097), .Z(n6300) );
  NANDN U6368 ( .A(n6100), .B(n6099), .Z(n6104) );
  NANDN U6369 ( .A(n6102), .B(n6101), .Z(n6103) );
  AND U6370 ( .A(n6104), .B(n6103), .Z(n6185) );
  NANDN U6371 ( .A(n6106), .B(n6105), .Z(n6110) );
  OR U6372 ( .A(n6108), .B(n6107), .Z(n6109) );
  AND U6373 ( .A(n6110), .B(n6109), .Z(n6183) );
  NANDN U6374 ( .A(n6112), .B(n6111), .Z(n6116) );
  NANDN U6375 ( .A(n6114), .B(n6113), .Z(n6115) );
  AND U6376 ( .A(n6116), .B(n6115), .Z(n6249) );
  NANDN U6377 ( .A(n6118), .B(n6117), .Z(n6122) );
  NANDN U6378 ( .A(n6120), .B(n6119), .Z(n6121) );
  NAND U6379 ( .A(n6122), .B(n6121), .Z(n6248) );
  XNOR U6380 ( .A(n6249), .B(n6248), .Z(n6251) );
  NAND U6381 ( .A(b[0]), .B(a[56]), .Z(n6123) );
  XNOR U6382 ( .A(b[1]), .B(n6123), .Z(n6125) );
  NANDN U6383 ( .A(b[0]), .B(a[55]), .Z(n6124) );
  NAND U6384 ( .A(n6125), .B(n6124), .Z(n6197) );
  NANDN U6385 ( .A(n19394), .B(n6126), .Z(n6128) );
  XOR U6386 ( .A(b[29]), .B(a[28]), .Z(n6270) );
  NANDN U6387 ( .A(n19395), .B(n6270), .Z(n6127) );
  AND U6388 ( .A(n6128), .B(n6127), .Z(n6195) );
  AND U6389 ( .A(b[31]), .B(a[24]), .Z(n6194) );
  XNOR U6390 ( .A(n6195), .B(n6194), .Z(n6196) );
  XNOR U6391 ( .A(n6197), .B(n6196), .Z(n6237) );
  NANDN U6392 ( .A(n19005), .B(n6129), .Z(n6131) );
  XOR U6393 ( .A(b[23]), .B(a[34]), .Z(n6276) );
  NANDN U6394 ( .A(n19055), .B(n6276), .Z(n6130) );
  AND U6395 ( .A(n6131), .B(n6130), .Z(n6266) );
  NANDN U6396 ( .A(n17362), .B(n6132), .Z(n6134) );
  XOR U6397 ( .A(b[7]), .B(a[50]), .Z(n6279) );
  NANDN U6398 ( .A(n17522), .B(n6279), .Z(n6133) );
  AND U6399 ( .A(n6134), .B(n6133), .Z(n6265) );
  NANDN U6400 ( .A(n19116), .B(n6135), .Z(n6137) );
  XOR U6401 ( .A(b[25]), .B(a[32]), .Z(n6282) );
  NANDN U6402 ( .A(n19179), .B(n6282), .Z(n6136) );
  NAND U6403 ( .A(n6137), .B(n6136), .Z(n6264) );
  XOR U6404 ( .A(n6265), .B(n6264), .Z(n6267) );
  XOR U6405 ( .A(n6266), .B(n6267), .Z(n6236) );
  XOR U6406 ( .A(n6237), .B(n6236), .Z(n6239) );
  NANDN U6407 ( .A(n18113), .B(n6138), .Z(n6140) );
  XOR U6408 ( .A(b[13]), .B(a[44]), .Z(n6285) );
  NANDN U6409 ( .A(n18229), .B(n6285), .Z(n6139) );
  AND U6410 ( .A(n6140), .B(n6139), .Z(n6231) );
  NANDN U6411 ( .A(n17888), .B(n6141), .Z(n6143) );
  XOR U6412 ( .A(b[11]), .B(a[46]), .Z(n6288) );
  NANDN U6413 ( .A(n18025), .B(n6288), .Z(n6142) );
  NAND U6414 ( .A(n6143), .B(n6142), .Z(n6230) );
  XNOR U6415 ( .A(n6231), .B(n6230), .Z(n6233) );
  NANDN U6416 ( .A(n18487), .B(n6144), .Z(n6146) );
  XOR U6417 ( .A(b[15]), .B(a[42]), .Z(n6291) );
  NANDN U6418 ( .A(n18311), .B(n6291), .Z(n6145) );
  AND U6419 ( .A(n6146), .B(n6145), .Z(n6227) );
  NANDN U6420 ( .A(n18853), .B(n6147), .Z(n6149) );
  XOR U6421 ( .A(b[21]), .B(a[36]), .Z(n6294) );
  NANDN U6422 ( .A(n18926), .B(n6294), .Z(n6148) );
  AND U6423 ( .A(n6149), .B(n6148), .Z(n6225) );
  NANDN U6424 ( .A(n17613), .B(n6150), .Z(n6152) );
  XOR U6425 ( .A(b[9]), .B(a[48]), .Z(n6297) );
  NANDN U6426 ( .A(n17739), .B(n6297), .Z(n6151) );
  NAND U6427 ( .A(n6152), .B(n6151), .Z(n6224) );
  XNOR U6428 ( .A(n6225), .B(n6224), .Z(n6226) );
  XNOR U6429 ( .A(n6227), .B(n6226), .Z(n6232) );
  XOR U6430 ( .A(n6233), .B(n6232), .Z(n6238) );
  XOR U6431 ( .A(n6239), .B(n6238), .Z(n6250) );
  XOR U6432 ( .A(n6251), .B(n6250), .Z(n6182) );
  XNOR U6433 ( .A(n6183), .B(n6182), .Z(n6184) );
  XOR U6434 ( .A(n6185), .B(n6184), .Z(n6301) );
  XNOR U6435 ( .A(n6300), .B(n6301), .Z(n6302) );
  XNOR U6436 ( .A(n6303), .B(n6302), .Z(n6178) );
  XOR U6437 ( .A(n6179), .B(n6178), .Z(n6171) );
  NANDN U6438 ( .A(n6154), .B(n6153), .Z(n6158) );
  NANDN U6439 ( .A(n6156), .B(n6155), .Z(n6157) );
  AND U6440 ( .A(n6158), .B(n6157), .Z(n6170) );
  XOR U6441 ( .A(n6171), .B(n6170), .Z(n6173) );
  XNOR U6442 ( .A(n6172), .B(n6173), .Z(n6164) );
  XNOR U6443 ( .A(n6165), .B(n6164), .Z(n6166) );
  XNOR U6444 ( .A(n6167), .B(n6166), .Z(n6306) );
  XNOR U6445 ( .A(sreg[152]), .B(n6306), .Z(n6308) );
  NANDN U6446 ( .A(sreg[151]), .B(n6159), .Z(n6163) );
  NAND U6447 ( .A(n6161), .B(n6160), .Z(n6162) );
  NAND U6448 ( .A(n6163), .B(n6162), .Z(n6307) );
  XNOR U6449 ( .A(n6308), .B(n6307), .Z(c[152]) );
  NANDN U6450 ( .A(n6165), .B(n6164), .Z(n6169) );
  NANDN U6451 ( .A(n6167), .B(n6166), .Z(n6168) );
  AND U6452 ( .A(n6169), .B(n6168), .Z(n6314) );
  NANDN U6453 ( .A(n6171), .B(n6170), .Z(n6175) );
  NANDN U6454 ( .A(n6173), .B(n6172), .Z(n6174) );
  AND U6455 ( .A(n6175), .B(n6174), .Z(n6312) );
  NANDN U6456 ( .A(n6177), .B(n6176), .Z(n6181) );
  NAND U6457 ( .A(n6179), .B(n6178), .Z(n6180) );
  AND U6458 ( .A(n6181), .B(n6180), .Z(n6319) );
  NANDN U6459 ( .A(n6183), .B(n6182), .Z(n6187) );
  NANDN U6460 ( .A(n6185), .B(n6184), .Z(n6186) );
  AND U6461 ( .A(n6187), .B(n6186), .Z(n6450) );
  NANDN U6462 ( .A(n6189), .B(n6188), .Z(n6193) );
  NAND U6463 ( .A(n6191), .B(n6190), .Z(n6192) );
  AND U6464 ( .A(n6193), .B(n6192), .Z(n6449) );
  XNOR U6465 ( .A(n6450), .B(n6449), .Z(n6452) );
  NANDN U6466 ( .A(n6195), .B(n6194), .Z(n6199) );
  NANDN U6467 ( .A(n6197), .B(n6196), .Z(n6198) );
  AND U6468 ( .A(n6199), .B(n6198), .Z(n6385) );
  NANDN U6469 ( .A(n19237), .B(n6200), .Z(n6202) );
  XOR U6470 ( .A(b[27]), .B(a[31]), .Z(n6329) );
  NANDN U6471 ( .A(n19277), .B(n6329), .Z(n6201) );
  AND U6472 ( .A(n6202), .B(n6201), .Z(n6392) );
  NANDN U6473 ( .A(n17072), .B(n6203), .Z(n6205) );
  XOR U6474 ( .A(b[5]), .B(a[53]), .Z(n6332) );
  NANDN U6475 ( .A(n17223), .B(n6332), .Z(n6204) );
  AND U6476 ( .A(n6205), .B(n6204), .Z(n6390) );
  NANDN U6477 ( .A(n18673), .B(n6206), .Z(n6208) );
  XOR U6478 ( .A(b[19]), .B(a[39]), .Z(n6335) );
  NANDN U6479 ( .A(n18758), .B(n6335), .Z(n6207) );
  NAND U6480 ( .A(n6208), .B(n6207), .Z(n6389) );
  XNOR U6481 ( .A(n6390), .B(n6389), .Z(n6391) );
  XNOR U6482 ( .A(n6392), .B(n6391), .Z(n6383) );
  NANDN U6483 ( .A(n19425), .B(n6209), .Z(n6211) );
  XOR U6484 ( .A(b[31]), .B(a[27]), .Z(n6338) );
  NANDN U6485 ( .A(n19426), .B(n6338), .Z(n6210) );
  AND U6486 ( .A(n6211), .B(n6210), .Z(n6350) );
  NANDN U6487 ( .A(n17067), .B(n6212), .Z(n6214) );
  XOR U6488 ( .A(b[3]), .B(a[55]), .Z(n6341) );
  NANDN U6489 ( .A(n17068), .B(n6341), .Z(n6213) );
  AND U6490 ( .A(n6214), .B(n6213), .Z(n6348) );
  NANDN U6491 ( .A(n18514), .B(n6215), .Z(n6217) );
  XOR U6492 ( .A(b[17]), .B(a[41]), .Z(n6344) );
  NANDN U6493 ( .A(n18585), .B(n6344), .Z(n6216) );
  NAND U6494 ( .A(n6217), .B(n6216), .Z(n6347) );
  XNOR U6495 ( .A(n6348), .B(n6347), .Z(n6349) );
  XOR U6496 ( .A(n6350), .B(n6349), .Z(n6384) );
  XOR U6497 ( .A(n6383), .B(n6384), .Z(n6386) );
  XOR U6498 ( .A(n6385), .B(n6386), .Z(n6432) );
  NANDN U6499 ( .A(n6219), .B(n6218), .Z(n6223) );
  NANDN U6500 ( .A(n6221), .B(n6220), .Z(n6222) );
  AND U6501 ( .A(n6223), .B(n6222), .Z(n6371) );
  NANDN U6502 ( .A(n6225), .B(n6224), .Z(n6229) );
  NANDN U6503 ( .A(n6227), .B(n6226), .Z(n6228) );
  NAND U6504 ( .A(n6229), .B(n6228), .Z(n6372) );
  XNOR U6505 ( .A(n6371), .B(n6372), .Z(n6373) );
  NANDN U6506 ( .A(n6231), .B(n6230), .Z(n6235) );
  NAND U6507 ( .A(n6233), .B(n6232), .Z(n6234) );
  NAND U6508 ( .A(n6235), .B(n6234), .Z(n6374) );
  XNOR U6509 ( .A(n6373), .B(n6374), .Z(n6431) );
  XNOR U6510 ( .A(n6432), .B(n6431), .Z(n6434) );
  NAND U6511 ( .A(n6237), .B(n6236), .Z(n6241) );
  NAND U6512 ( .A(n6239), .B(n6238), .Z(n6240) );
  AND U6513 ( .A(n6241), .B(n6240), .Z(n6433) );
  XOR U6514 ( .A(n6434), .B(n6433), .Z(n6446) );
  NANDN U6515 ( .A(n6243), .B(n6242), .Z(n6247) );
  NANDN U6516 ( .A(n6245), .B(n6244), .Z(n6246) );
  AND U6517 ( .A(n6247), .B(n6246), .Z(n6443) );
  NANDN U6518 ( .A(n6253), .B(n6252), .Z(n6257) );
  OR U6519 ( .A(n6255), .B(n6254), .Z(n6256) );
  AND U6520 ( .A(n6257), .B(n6256), .Z(n6438) );
  NANDN U6521 ( .A(n6259), .B(n6258), .Z(n6263) );
  NANDN U6522 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U6523 ( .A(n6263), .B(n6262), .Z(n6378) );
  NANDN U6524 ( .A(n6265), .B(n6264), .Z(n6269) );
  OR U6525 ( .A(n6267), .B(n6266), .Z(n6268) );
  NAND U6526 ( .A(n6269), .B(n6268), .Z(n6377) );
  XNOR U6527 ( .A(n6378), .B(n6377), .Z(n6379) );
  NANDN U6528 ( .A(n19394), .B(n6270), .Z(n6272) );
  XOR U6529 ( .A(b[29]), .B(a[29]), .Z(n6404) );
  NANDN U6530 ( .A(n19395), .B(n6404), .Z(n6271) );
  AND U6531 ( .A(n6272), .B(n6271), .Z(n6324) );
  AND U6532 ( .A(b[31]), .B(a[25]), .Z(n6323) );
  XNOR U6533 ( .A(n6324), .B(n6323), .Z(n6325) );
  NAND U6534 ( .A(b[0]), .B(a[57]), .Z(n6273) );
  XNOR U6535 ( .A(b[1]), .B(n6273), .Z(n6275) );
  NANDN U6536 ( .A(b[0]), .B(a[56]), .Z(n6274) );
  NAND U6537 ( .A(n6275), .B(n6274), .Z(n6326) );
  XNOR U6538 ( .A(n6325), .B(n6326), .Z(n6365) );
  NANDN U6539 ( .A(n19005), .B(n6276), .Z(n6278) );
  XOR U6540 ( .A(b[23]), .B(a[35]), .Z(n6407) );
  NANDN U6541 ( .A(n19055), .B(n6407), .Z(n6277) );
  AND U6542 ( .A(n6278), .B(n6277), .Z(n6398) );
  NANDN U6543 ( .A(n17362), .B(n6279), .Z(n6281) );
  XOR U6544 ( .A(b[7]), .B(a[51]), .Z(n6410) );
  NANDN U6545 ( .A(n17522), .B(n6410), .Z(n6280) );
  AND U6546 ( .A(n6281), .B(n6280), .Z(n6396) );
  NANDN U6547 ( .A(n19116), .B(n6282), .Z(n6284) );
  XOR U6548 ( .A(b[25]), .B(a[33]), .Z(n6413) );
  NANDN U6549 ( .A(n19179), .B(n6413), .Z(n6283) );
  NAND U6550 ( .A(n6284), .B(n6283), .Z(n6395) );
  XNOR U6551 ( .A(n6396), .B(n6395), .Z(n6397) );
  XOR U6552 ( .A(n6398), .B(n6397), .Z(n6366) );
  XNOR U6553 ( .A(n6365), .B(n6366), .Z(n6367) );
  NANDN U6554 ( .A(n18113), .B(n6285), .Z(n6287) );
  XOR U6555 ( .A(b[13]), .B(a[45]), .Z(n6416) );
  NANDN U6556 ( .A(n18229), .B(n6416), .Z(n6286) );
  AND U6557 ( .A(n6287), .B(n6286), .Z(n6360) );
  NANDN U6558 ( .A(n17888), .B(n6288), .Z(n6290) );
  XOR U6559 ( .A(b[11]), .B(a[47]), .Z(n6419) );
  NANDN U6560 ( .A(n18025), .B(n6419), .Z(n6289) );
  NAND U6561 ( .A(n6290), .B(n6289), .Z(n6359) );
  XNOR U6562 ( .A(n6360), .B(n6359), .Z(n6361) );
  NANDN U6563 ( .A(n18487), .B(n6291), .Z(n6293) );
  XOR U6564 ( .A(b[15]), .B(a[43]), .Z(n6422) );
  NANDN U6565 ( .A(n18311), .B(n6422), .Z(n6292) );
  AND U6566 ( .A(n6293), .B(n6292), .Z(n6356) );
  NANDN U6567 ( .A(n18853), .B(n6294), .Z(n6296) );
  XOR U6568 ( .A(b[21]), .B(a[37]), .Z(n6425) );
  NANDN U6569 ( .A(n18926), .B(n6425), .Z(n6295) );
  AND U6570 ( .A(n6296), .B(n6295), .Z(n6354) );
  NANDN U6571 ( .A(n17613), .B(n6297), .Z(n6299) );
  XOR U6572 ( .A(b[9]), .B(a[49]), .Z(n6428) );
  NANDN U6573 ( .A(n17739), .B(n6428), .Z(n6298) );
  NAND U6574 ( .A(n6299), .B(n6298), .Z(n6353) );
  XNOR U6575 ( .A(n6354), .B(n6353), .Z(n6355) );
  XOR U6576 ( .A(n6356), .B(n6355), .Z(n6362) );
  XOR U6577 ( .A(n6361), .B(n6362), .Z(n6368) );
  XOR U6578 ( .A(n6367), .B(n6368), .Z(n6380) );
  XNOR U6579 ( .A(n6379), .B(n6380), .Z(n6437) );
  XNOR U6580 ( .A(n6438), .B(n6437), .Z(n6439) );
  XOR U6581 ( .A(n6440), .B(n6439), .Z(n6444) );
  XNOR U6582 ( .A(n6443), .B(n6444), .Z(n6445) );
  XNOR U6583 ( .A(n6446), .B(n6445), .Z(n6451) );
  XOR U6584 ( .A(n6452), .B(n6451), .Z(n6318) );
  NANDN U6585 ( .A(n6301), .B(n6300), .Z(n6305) );
  NANDN U6586 ( .A(n6303), .B(n6302), .Z(n6304) );
  AND U6587 ( .A(n6305), .B(n6304), .Z(n6317) );
  XOR U6588 ( .A(n6318), .B(n6317), .Z(n6320) );
  XNOR U6589 ( .A(n6319), .B(n6320), .Z(n6311) );
  XNOR U6590 ( .A(n6312), .B(n6311), .Z(n6313) );
  XNOR U6591 ( .A(n6314), .B(n6313), .Z(n6455) );
  XNOR U6592 ( .A(sreg[153]), .B(n6455), .Z(n6457) );
  NANDN U6593 ( .A(sreg[152]), .B(n6306), .Z(n6310) );
  NAND U6594 ( .A(n6308), .B(n6307), .Z(n6309) );
  NAND U6595 ( .A(n6310), .B(n6309), .Z(n6456) );
  XNOR U6596 ( .A(n6457), .B(n6456), .Z(c[153]) );
  NANDN U6597 ( .A(n6312), .B(n6311), .Z(n6316) );
  NANDN U6598 ( .A(n6314), .B(n6313), .Z(n6315) );
  AND U6599 ( .A(n6316), .B(n6315), .Z(n6463) );
  NANDN U6600 ( .A(n6318), .B(n6317), .Z(n6322) );
  NANDN U6601 ( .A(n6320), .B(n6319), .Z(n6321) );
  AND U6602 ( .A(n6322), .B(n6321), .Z(n6461) );
  NANDN U6603 ( .A(n6324), .B(n6323), .Z(n6328) );
  NANDN U6604 ( .A(n6326), .B(n6325), .Z(n6327) );
  AND U6605 ( .A(n6328), .B(n6327), .Z(n6552) );
  NANDN U6606 ( .A(n19237), .B(n6329), .Z(n6331) );
  XOR U6607 ( .A(b[27]), .B(a[32]), .Z(n6496) );
  NANDN U6608 ( .A(n19277), .B(n6496), .Z(n6330) );
  AND U6609 ( .A(n6331), .B(n6330), .Z(n6559) );
  NANDN U6610 ( .A(n17072), .B(n6332), .Z(n6334) );
  XOR U6611 ( .A(b[5]), .B(a[54]), .Z(n6499) );
  NANDN U6612 ( .A(n17223), .B(n6499), .Z(n6333) );
  AND U6613 ( .A(n6334), .B(n6333), .Z(n6557) );
  NANDN U6614 ( .A(n18673), .B(n6335), .Z(n6337) );
  XOR U6615 ( .A(b[19]), .B(a[40]), .Z(n6502) );
  NANDN U6616 ( .A(n18758), .B(n6502), .Z(n6336) );
  NAND U6617 ( .A(n6337), .B(n6336), .Z(n6556) );
  XNOR U6618 ( .A(n6557), .B(n6556), .Z(n6558) );
  XNOR U6619 ( .A(n6559), .B(n6558), .Z(n6550) );
  NANDN U6620 ( .A(n19425), .B(n6338), .Z(n6340) );
  XOR U6621 ( .A(b[31]), .B(a[28]), .Z(n6505) );
  NANDN U6622 ( .A(n19426), .B(n6505), .Z(n6339) );
  AND U6623 ( .A(n6340), .B(n6339), .Z(n6517) );
  NANDN U6624 ( .A(n17067), .B(n6341), .Z(n6343) );
  XOR U6625 ( .A(b[3]), .B(a[56]), .Z(n6508) );
  NANDN U6626 ( .A(n17068), .B(n6508), .Z(n6342) );
  AND U6627 ( .A(n6343), .B(n6342), .Z(n6515) );
  NANDN U6628 ( .A(n18514), .B(n6344), .Z(n6346) );
  XOR U6629 ( .A(b[17]), .B(a[42]), .Z(n6511) );
  NANDN U6630 ( .A(n18585), .B(n6511), .Z(n6345) );
  NAND U6631 ( .A(n6346), .B(n6345), .Z(n6514) );
  XNOR U6632 ( .A(n6515), .B(n6514), .Z(n6516) );
  XOR U6633 ( .A(n6517), .B(n6516), .Z(n6551) );
  XOR U6634 ( .A(n6550), .B(n6551), .Z(n6553) );
  XOR U6635 ( .A(n6552), .B(n6553), .Z(n6485) );
  NANDN U6636 ( .A(n6348), .B(n6347), .Z(n6352) );
  NANDN U6637 ( .A(n6350), .B(n6349), .Z(n6351) );
  AND U6638 ( .A(n6352), .B(n6351), .Z(n6538) );
  NANDN U6639 ( .A(n6354), .B(n6353), .Z(n6358) );
  NANDN U6640 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U6641 ( .A(n6358), .B(n6357), .Z(n6539) );
  XNOR U6642 ( .A(n6538), .B(n6539), .Z(n6540) );
  NANDN U6643 ( .A(n6360), .B(n6359), .Z(n6364) );
  NANDN U6644 ( .A(n6362), .B(n6361), .Z(n6363) );
  NAND U6645 ( .A(n6364), .B(n6363), .Z(n6541) );
  XNOR U6646 ( .A(n6540), .B(n6541), .Z(n6484) );
  XNOR U6647 ( .A(n6485), .B(n6484), .Z(n6487) );
  NANDN U6648 ( .A(n6366), .B(n6365), .Z(n6370) );
  NANDN U6649 ( .A(n6368), .B(n6367), .Z(n6369) );
  AND U6650 ( .A(n6370), .B(n6369), .Z(n6486) );
  XOR U6651 ( .A(n6487), .B(n6486), .Z(n6600) );
  NANDN U6652 ( .A(n6372), .B(n6371), .Z(n6376) );
  NANDN U6653 ( .A(n6374), .B(n6373), .Z(n6375) );
  AND U6654 ( .A(n6376), .B(n6375), .Z(n6598) );
  NANDN U6655 ( .A(n6378), .B(n6377), .Z(n6382) );
  NANDN U6656 ( .A(n6380), .B(n6379), .Z(n6381) );
  AND U6657 ( .A(n6382), .B(n6381), .Z(n6481) );
  NANDN U6658 ( .A(n6384), .B(n6383), .Z(n6388) );
  OR U6659 ( .A(n6386), .B(n6385), .Z(n6387) );
  AND U6660 ( .A(n6388), .B(n6387), .Z(n6479) );
  NANDN U6661 ( .A(n6390), .B(n6389), .Z(n6394) );
  NANDN U6662 ( .A(n6392), .B(n6391), .Z(n6393) );
  AND U6663 ( .A(n6394), .B(n6393), .Z(n6545) );
  NANDN U6664 ( .A(n6396), .B(n6395), .Z(n6400) );
  NANDN U6665 ( .A(n6398), .B(n6397), .Z(n6399) );
  NAND U6666 ( .A(n6400), .B(n6399), .Z(n6544) );
  XNOR U6667 ( .A(n6545), .B(n6544), .Z(n6546) );
  NAND U6668 ( .A(b[0]), .B(a[58]), .Z(n6401) );
  XNOR U6669 ( .A(b[1]), .B(n6401), .Z(n6403) );
  NANDN U6670 ( .A(b[0]), .B(a[57]), .Z(n6402) );
  NAND U6671 ( .A(n6403), .B(n6402), .Z(n6493) );
  NANDN U6672 ( .A(n19394), .B(n6404), .Z(n6406) );
  XOR U6673 ( .A(b[29]), .B(a[30]), .Z(n6571) );
  NANDN U6674 ( .A(n19395), .B(n6571), .Z(n6405) );
  AND U6675 ( .A(n6406), .B(n6405), .Z(n6491) );
  AND U6676 ( .A(b[31]), .B(a[26]), .Z(n6490) );
  XNOR U6677 ( .A(n6491), .B(n6490), .Z(n6492) );
  XNOR U6678 ( .A(n6493), .B(n6492), .Z(n6532) );
  NANDN U6679 ( .A(n19005), .B(n6407), .Z(n6409) );
  XOR U6680 ( .A(b[23]), .B(a[36]), .Z(n6574) );
  NANDN U6681 ( .A(n19055), .B(n6574), .Z(n6408) );
  AND U6682 ( .A(n6409), .B(n6408), .Z(n6565) );
  NANDN U6683 ( .A(n17362), .B(n6410), .Z(n6412) );
  XOR U6684 ( .A(b[7]), .B(a[52]), .Z(n6577) );
  NANDN U6685 ( .A(n17522), .B(n6577), .Z(n6411) );
  AND U6686 ( .A(n6412), .B(n6411), .Z(n6563) );
  NANDN U6687 ( .A(n19116), .B(n6413), .Z(n6415) );
  XOR U6688 ( .A(b[25]), .B(a[34]), .Z(n6580) );
  NANDN U6689 ( .A(n19179), .B(n6580), .Z(n6414) );
  NAND U6690 ( .A(n6415), .B(n6414), .Z(n6562) );
  XNOR U6691 ( .A(n6563), .B(n6562), .Z(n6564) );
  XOR U6692 ( .A(n6565), .B(n6564), .Z(n6533) );
  XNOR U6693 ( .A(n6532), .B(n6533), .Z(n6534) );
  NANDN U6694 ( .A(n18113), .B(n6416), .Z(n6418) );
  XOR U6695 ( .A(b[13]), .B(a[46]), .Z(n6583) );
  NANDN U6696 ( .A(n18229), .B(n6583), .Z(n6417) );
  AND U6697 ( .A(n6418), .B(n6417), .Z(n6527) );
  NANDN U6698 ( .A(n17888), .B(n6419), .Z(n6421) );
  XOR U6699 ( .A(b[11]), .B(a[48]), .Z(n6586) );
  NANDN U6700 ( .A(n18025), .B(n6586), .Z(n6420) );
  NAND U6701 ( .A(n6421), .B(n6420), .Z(n6526) );
  XNOR U6702 ( .A(n6527), .B(n6526), .Z(n6528) );
  NANDN U6703 ( .A(n18487), .B(n6422), .Z(n6424) );
  XOR U6704 ( .A(b[15]), .B(a[44]), .Z(n6589) );
  NANDN U6705 ( .A(n18311), .B(n6589), .Z(n6423) );
  AND U6706 ( .A(n6424), .B(n6423), .Z(n6523) );
  NANDN U6707 ( .A(n18853), .B(n6425), .Z(n6427) );
  XOR U6708 ( .A(b[21]), .B(a[38]), .Z(n6592) );
  NANDN U6709 ( .A(n18926), .B(n6592), .Z(n6426) );
  AND U6710 ( .A(n6427), .B(n6426), .Z(n6521) );
  NANDN U6711 ( .A(n17613), .B(n6428), .Z(n6430) );
  XOR U6712 ( .A(b[9]), .B(a[50]), .Z(n6595) );
  NANDN U6713 ( .A(n17739), .B(n6595), .Z(n6429) );
  NAND U6714 ( .A(n6430), .B(n6429), .Z(n6520) );
  XNOR U6715 ( .A(n6521), .B(n6520), .Z(n6522) );
  XOR U6716 ( .A(n6523), .B(n6522), .Z(n6529) );
  XOR U6717 ( .A(n6528), .B(n6529), .Z(n6535) );
  XOR U6718 ( .A(n6534), .B(n6535), .Z(n6547) );
  XNOR U6719 ( .A(n6546), .B(n6547), .Z(n6478) );
  XNOR U6720 ( .A(n6479), .B(n6478), .Z(n6480) );
  XOR U6721 ( .A(n6481), .B(n6480), .Z(n6599) );
  XOR U6722 ( .A(n6598), .B(n6599), .Z(n6601) );
  XOR U6723 ( .A(n6600), .B(n6601), .Z(n6475) );
  NANDN U6724 ( .A(n6432), .B(n6431), .Z(n6436) );
  NAND U6725 ( .A(n6434), .B(n6433), .Z(n6435) );
  AND U6726 ( .A(n6436), .B(n6435), .Z(n6473) );
  NANDN U6727 ( .A(n6438), .B(n6437), .Z(n6442) );
  NANDN U6728 ( .A(n6440), .B(n6439), .Z(n6441) );
  AND U6729 ( .A(n6442), .B(n6441), .Z(n6472) );
  XNOR U6730 ( .A(n6473), .B(n6472), .Z(n6474) );
  XNOR U6731 ( .A(n6475), .B(n6474), .Z(n6466) );
  NANDN U6732 ( .A(n6444), .B(n6443), .Z(n6448) );
  NANDN U6733 ( .A(n6446), .B(n6445), .Z(n6447) );
  NAND U6734 ( .A(n6448), .B(n6447), .Z(n6467) );
  XNOR U6735 ( .A(n6466), .B(n6467), .Z(n6468) );
  NANDN U6736 ( .A(n6450), .B(n6449), .Z(n6454) );
  NAND U6737 ( .A(n6452), .B(n6451), .Z(n6453) );
  NAND U6738 ( .A(n6454), .B(n6453), .Z(n6469) );
  XNOR U6739 ( .A(n6468), .B(n6469), .Z(n6460) );
  XNOR U6740 ( .A(n6461), .B(n6460), .Z(n6462) );
  XNOR U6741 ( .A(n6463), .B(n6462), .Z(n6604) );
  XNOR U6742 ( .A(sreg[154]), .B(n6604), .Z(n6606) );
  NANDN U6743 ( .A(sreg[153]), .B(n6455), .Z(n6459) );
  NAND U6744 ( .A(n6457), .B(n6456), .Z(n6458) );
  NAND U6745 ( .A(n6459), .B(n6458), .Z(n6605) );
  XNOR U6746 ( .A(n6606), .B(n6605), .Z(c[154]) );
  NANDN U6747 ( .A(n6461), .B(n6460), .Z(n6465) );
  NANDN U6748 ( .A(n6463), .B(n6462), .Z(n6464) );
  AND U6749 ( .A(n6465), .B(n6464), .Z(n6612) );
  NANDN U6750 ( .A(n6467), .B(n6466), .Z(n6471) );
  NANDN U6751 ( .A(n6469), .B(n6468), .Z(n6470) );
  AND U6752 ( .A(n6471), .B(n6470), .Z(n6610) );
  NANDN U6753 ( .A(n6473), .B(n6472), .Z(n6477) );
  NANDN U6754 ( .A(n6475), .B(n6474), .Z(n6476) );
  AND U6755 ( .A(n6477), .B(n6476), .Z(n6618) );
  NANDN U6756 ( .A(n6479), .B(n6478), .Z(n6483) );
  NANDN U6757 ( .A(n6481), .B(n6480), .Z(n6482) );
  AND U6758 ( .A(n6483), .B(n6482), .Z(n6748) );
  NANDN U6759 ( .A(n6485), .B(n6484), .Z(n6489) );
  NAND U6760 ( .A(n6487), .B(n6486), .Z(n6488) );
  AND U6761 ( .A(n6489), .B(n6488), .Z(n6747) );
  XNOR U6762 ( .A(n6748), .B(n6747), .Z(n6750) );
  NANDN U6763 ( .A(n6491), .B(n6490), .Z(n6495) );
  NANDN U6764 ( .A(n6493), .B(n6492), .Z(n6494) );
  AND U6765 ( .A(n6495), .B(n6494), .Z(n6695) );
  NANDN U6766 ( .A(n19237), .B(n6496), .Z(n6498) );
  XOR U6767 ( .A(b[27]), .B(a[33]), .Z(n6639) );
  NANDN U6768 ( .A(n19277), .B(n6639), .Z(n6497) );
  AND U6769 ( .A(n6498), .B(n6497), .Z(n6702) );
  NANDN U6770 ( .A(n17072), .B(n6499), .Z(n6501) );
  XOR U6771 ( .A(b[5]), .B(a[55]), .Z(n6642) );
  NANDN U6772 ( .A(n17223), .B(n6642), .Z(n6500) );
  AND U6773 ( .A(n6501), .B(n6500), .Z(n6700) );
  NANDN U6774 ( .A(n18673), .B(n6502), .Z(n6504) );
  XOR U6775 ( .A(b[19]), .B(a[41]), .Z(n6645) );
  NANDN U6776 ( .A(n18758), .B(n6645), .Z(n6503) );
  NAND U6777 ( .A(n6504), .B(n6503), .Z(n6699) );
  XNOR U6778 ( .A(n6700), .B(n6699), .Z(n6701) );
  XNOR U6779 ( .A(n6702), .B(n6701), .Z(n6693) );
  NANDN U6780 ( .A(n19425), .B(n6505), .Z(n6507) );
  XOR U6781 ( .A(b[31]), .B(a[29]), .Z(n6648) );
  NANDN U6782 ( .A(n19426), .B(n6648), .Z(n6506) );
  AND U6783 ( .A(n6507), .B(n6506), .Z(n6660) );
  NANDN U6784 ( .A(n17067), .B(n6508), .Z(n6510) );
  XOR U6785 ( .A(b[3]), .B(a[57]), .Z(n6651) );
  NANDN U6786 ( .A(n17068), .B(n6651), .Z(n6509) );
  AND U6787 ( .A(n6510), .B(n6509), .Z(n6658) );
  NANDN U6788 ( .A(n18514), .B(n6511), .Z(n6513) );
  XOR U6789 ( .A(b[17]), .B(a[43]), .Z(n6654) );
  NANDN U6790 ( .A(n18585), .B(n6654), .Z(n6512) );
  NAND U6791 ( .A(n6513), .B(n6512), .Z(n6657) );
  XNOR U6792 ( .A(n6658), .B(n6657), .Z(n6659) );
  XOR U6793 ( .A(n6660), .B(n6659), .Z(n6694) );
  XOR U6794 ( .A(n6693), .B(n6694), .Z(n6696) );
  XOR U6795 ( .A(n6695), .B(n6696), .Z(n6628) );
  NANDN U6796 ( .A(n6515), .B(n6514), .Z(n6519) );
  NANDN U6797 ( .A(n6517), .B(n6516), .Z(n6518) );
  AND U6798 ( .A(n6519), .B(n6518), .Z(n6681) );
  NANDN U6799 ( .A(n6521), .B(n6520), .Z(n6525) );
  NANDN U6800 ( .A(n6523), .B(n6522), .Z(n6524) );
  NAND U6801 ( .A(n6525), .B(n6524), .Z(n6682) );
  XNOR U6802 ( .A(n6681), .B(n6682), .Z(n6683) );
  NANDN U6803 ( .A(n6527), .B(n6526), .Z(n6531) );
  NANDN U6804 ( .A(n6529), .B(n6528), .Z(n6530) );
  NAND U6805 ( .A(n6531), .B(n6530), .Z(n6684) );
  XNOR U6806 ( .A(n6683), .B(n6684), .Z(n6627) );
  XNOR U6807 ( .A(n6628), .B(n6627), .Z(n6630) );
  NANDN U6808 ( .A(n6533), .B(n6532), .Z(n6537) );
  NANDN U6809 ( .A(n6535), .B(n6534), .Z(n6536) );
  AND U6810 ( .A(n6537), .B(n6536), .Z(n6629) );
  XOR U6811 ( .A(n6630), .B(n6629), .Z(n6744) );
  NANDN U6812 ( .A(n6539), .B(n6538), .Z(n6543) );
  NANDN U6813 ( .A(n6541), .B(n6540), .Z(n6542) );
  AND U6814 ( .A(n6543), .B(n6542), .Z(n6741) );
  NANDN U6815 ( .A(n6545), .B(n6544), .Z(n6549) );
  NANDN U6816 ( .A(n6547), .B(n6546), .Z(n6548) );
  AND U6817 ( .A(n6549), .B(n6548), .Z(n6624) );
  NANDN U6818 ( .A(n6551), .B(n6550), .Z(n6555) );
  OR U6819 ( .A(n6553), .B(n6552), .Z(n6554) );
  AND U6820 ( .A(n6555), .B(n6554), .Z(n6622) );
  NANDN U6821 ( .A(n6557), .B(n6556), .Z(n6561) );
  NANDN U6822 ( .A(n6559), .B(n6558), .Z(n6560) );
  AND U6823 ( .A(n6561), .B(n6560), .Z(n6688) );
  NANDN U6824 ( .A(n6563), .B(n6562), .Z(n6567) );
  NANDN U6825 ( .A(n6565), .B(n6564), .Z(n6566) );
  NAND U6826 ( .A(n6567), .B(n6566), .Z(n6687) );
  XNOR U6827 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U6828 ( .A(b[0]), .B(a[59]), .Z(n6568) );
  XNOR U6829 ( .A(b[1]), .B(n6568), .Z(n6570) );
  NANDN U6830 ( .A(b[0]), .B(a[58]), .Z(n6569) );
  NAND U6831 ( .A(n6570), .B(n6569), .Z(n6636) );
  NANDN U6832 ( .A(n19394), .B(n6571), .Z(n6573) );
  XOR U6833 ( .A(b[29]), .B(a[31]), .Z(n6714) );
  NANDN U6834 ( .A(n19395), .B(n6714), .Z(n6572) );
  AND U6835 ( .A(n6573), .B(n6572), .Z(n6634) );
  AND U6836 ( .A(b[31]), .B(a[27]), .Z(n6633) );
  XNOR U6837 ( .A(n6634), .B(n6633), .Z(n6635) );
  XNOR U6838 ( .A(n6636), .B(n6635), .Z(n6675) );
  NANDN U6839 ( .A(n19005), .B(n6574), .Z(n6576) );
  XOR U6840 ( .A(b[23]), .B(a[37]), .Z(n6717) );
  NANDN U6841 ( .A(n19055), .B(n6717), .Z(n6575) );
  AND U6842 ( .A(n6576), .B(n6575), .Z(n6708) );
  NANDN U6843 ( .A(n17362), .B(n6577), .Z(n6579) );
  XOR U6844 ( .A(b[7]), .B(a[53]), .Z(n6720) );
  NANDN U6845 ( .A(n17522), .B(n6720), .Z(n6578) );
  AND U6846 ( .A(n6579), .B(n6578), .Z(n6706) );
  NANDN U6847 ( .A(n19116), .B(n6580), .Z(n6582) );
  XOR U6848 ( .A(b[25]), .B(a[35]), .Z(n6723) );
  NANDN U6849 ( .A(n19179), .B(n6723), .Z(n6581) );
  NAND U6850 ( .A(n6582), .B(n6581), .Z(n6705) );
  XNOR U6851 ( .A(n6706), .B(n6705), .Z(n6707) );
  XOR U6852 ( .A(n6708), .B(n6707), .Z(n6676) );
  XNOR U6853 ( .A(n6675), .B(n6676), .Z(n6677) );
  NANDN U6854 ( .A(n18113), .B(n6583), .Z(n6585) );
  XOR U6855 ( .A(b[13]), .B(a[47]), .Z(n6726) );
  NANDN U6856 ( .A(n18229), .B(n6726), .Z(n6584) );
  AND U6857 ( .A(n6585), .B(n6584), .Z(n6670) );
  NANDN U6858 ( .A(n17888), .B(n6586), .Z(n6588) );
  XOR U6859 ( .A(b[11]), .B(a[49]), .Z(n6729) );
  NANDN U6860 ( .A(n18025), .B(n6729), .Z(n6587) );
  NAND U6861 ( .A(n6588), .B(n6587), .Z(n6669) );
  XNOR U6862 ( .A(n6670), .B(n6669), .Z(n6671) );
  NANDN U6863 ( .A(n18487), .B(n6589), .Z(n6591) );
  XOR U6864 ( .A(b[15]), .B(a[45]), .Z(n6732) );
  NANDN U6865 ( .A(n18311), .B(n6732), .Z(n6590) );
  AND U6866 ( .A(n6591), .B(n6590), .Z(n6666) );
  NANDN U6867 ( .A(n18853), .B(n6592), .Z(n6594) );
  XOR U6868 ( .A(b[21]), .B(a[39]), .Z(n6735) );
  NANDN U6869 ( .A(n18926), .B(n6735), .Z(n6593) );
  AND U6870 ( .A(n6594), .B(n6593), .Z(n6664) );
  NANDN U6871 ( .A(n17613), .B(n6595), .Z(n6597) );
  XOR U6872 ( .A(b[9]), .B(a[51]), .Z(n6738) );
  NANDN U6873 ( .A(n17739), .B(n6738), .Z(n6596) );
  NAND U6874 ( .A(n6597), .B(n6596), .Z(n6663) );
  XNOR U6875 ( .A(n6664), .B(n6663), .Z(n6665) );
  XOR U6876 ( .A(n6666), .B(n6665), .Z(n6672) );
  XOR U6877 ( .A(n6671), .B(n6672), .Z(n6678) );
  XOR U6878 ( .A(n6677), .B(n6678), .Z(n6690) );
  XNOR U6879 ( .A(n6689), .B(n6690), .Z(n6621) );
  XNOR U6880 ( .A(n6622), .B(n6621), .Z(n6623) );
  XOR U6881 ( .A(n6624), .B(n6623), .Z(n6742) );
  XNOR U6882 ( .A(n6741), .B(n6742), .Z(n6743) );
  XNOR U6883 ( .A(n6744), .B(n6743), .Z(n6749) );
  XOR U6884 ( .A(n6750), .B(n6749), .Z(n6616) );
  NANDN U6885 ( .A(n6599), .B(n6598), .Z(n6603) );
  OR U6886 ( .A(n6601), .B(n6600), .Z(n6602) );
  AND U6887 ( .A(n6603), .B(n6602), .Z(n6615) );
  XNOR U6888 ( .A(n6616), .B(n6615), .Z(n6617) );
  XNOR U6889 ( .A(n6618), .B(n6617), .Z(n6609) );
  XNOR U6890 ( .A(n6610), .B(n6609), .Z(n6611) );
  XNOR U6891 ( .A(n6612), .B(n6611), .Z(n6753) );
  XNOR U6892 ( .A(sreg[155]), .B(n6753), .Z(n6755) );
  NANDN U6893 ( .A(sreg[154]), .B(n6604), .Z(n6608) );
  NAND U6894 ( .A(n6606), .B(n6605), .Z(n6607) );
  NAND U6895 ( .A(n6608), .B(n6607), .Z(n6754) );
  XNOR U6896 ( .A(n6755), .B(n6754), .Z(c[155]) );
  NANDN U6897 ( .A(n6610), .B(n6609), .Z(n6614) );
  NANDN U6898 ( .A(n6612), .B(n6611), .Z(n6613) );
  AND U6899 ( .A(n6614), .B(n6613), .Z(n6761) );
  NANDN U6900 ( .A(n6616), .B(n6615), .Z(n6620) );
  NANDN U6901 ( .A(n6618), .B(n6617), .Z(n6619) );
  AND U6902 ( .A(n6620), .B(n6619), .Z(n6759) );
  NANDN U6903 ( .A(n6622), .B(n6621), .Z(n6626) );
  NANDN U6904 ( .A(n6624), .B(n6623), .Z(n6625) );
  AND U6905 ( .A(n6626), .B(n6625), .Z(n6897) );
  NANDN U6906 ( .A(n6628), .B(n6627), .Z(n6632) );
  NAND U6907 ( .A(n6630), .B(n6629), .Z(n6631) );
  AND U6908 ( .A(n6632), .B(n6631), .Z(n6896) );
  XNOR U6909 ( .A(n6897), .B(n6896), .Z(n6899) );
  NANDN U6910 ( .A(n6634), .B(n6633), .Z(n6638) );
  NANDN U6911 ( .A(n6636), .B(n6635), .Z(n6637) );
  AND U6912 ( .A(n6638), .B(n6637), .Z(n6844) );
  NANDN U6913 ( .A(n19237), .B(n6639), .Z(n6641) );
  XOR U6914 ( .A(b[27]), .B(a[34]), .Z(n6788) );
  NANDN U6915 ( .A(n19277), .B(n6788), .Z(n6640) );
  AND U6916 ( .A(n6641), .B(n6640), .Z(n6851) );
  NANDN U6917 ( .A(n17072), .B(n6642), .Z(n6644) );
  XOR U6918 ( .A(b[5]), .B(a[56]), .Z(n6791) );
  NANDN U6919 ( .A(n17223), .B(n6791), .Z(n6643) );
  AND U6920 ( .A(n6644), .B(n6643), .Z(n6849) );
  NANDN U6921 ( .A(n18673), .B(n6645), .Z(n6647) );
  XOR U6922 ( .A(b[19]), .B(a[42]), .Z(n6794) );
  NANDN U6923 ( .A(n18758), .B(n6794), .Z(n6646) );
  NAND U6924 ( .A(n6647), .B(n6646), .Z(n6848) );
  XNOR U6925 ( .A(n6849), .B(n6848), .Z(n6850) );
  XNOR U6926 ( .A(n6851), .B(n6850), .Z(n6842) );
  NANDN U6927 ( .A(n19425), .B(n6648), .Z(n6650) );
  XOR U6928 ( .A(b[31]), .B(a[30]), .Z(n6797) );
  NANDN U6929 ( .A(n19426), .B(n6797), .Z(n6649) );
  AND U6930 ( .A(n6650), .B(n6649), .Z(n6809) );
  NANDN U6931 ( .A(n17067), .B(n6651), .Z(n6653) );
  XOR U6932 ( .A(b[3]), .B(a[58]), .Z(n6800) );
  NANDN U6933 ( .A(n17068), .B(n6800), .Z(n6652) );
  AND U6934 ( .A(n6653), .B(n6652), .Z(n6807) );
  NANDN U6935 ( .A(n18514), .B(n6654), .Z(n6656) );
  XOR U6936 ( .A(b[17]), .B(a[44]), .Z(n6803) );
  NANDN U6937 ( .A(n18585), .B(n6803), .Z(n6655) );
  NAND U6938 ( .A(n6656), .B(n6655), .Z(n6806) );
  XNOR U6939 ( .A(n6807), .B(n6806), .Z(n6808) );
  XOR U6940 ( .A(n6809), .B(n6808), .Z(n6843) );
  XOR U6941 ( .A(n6842), .B(n6843), .Z(n6845) );
  XOR U6942 ( .A(n6844), .B(n6845), .Z(n6777) );
  NANDN U6943 ( .A(n6658), .B(n6657), .Z(n6662) );
  NANDN U6944 ( .A(n6660), .B(n6659), .Z(n6661) );
  AND U6945 ( .A(n6662), .B(n6661), .Z(n6830) );
  NANDN U6946 ( .A(n6664), .B(n6663), .Z(n6668) );
  NANDN U6947 ( .A(n6666), .B(n6665), .Z(n6667) );
  NAND U6948 ( .A(n6668), .B(n6667), .Z(n6831) );
  XNOR U6949 ( .A(n6830), .B(n6831), .Z(n6832) );
  NANDN U6950 ( .A(n6670), .B(n6669), .Z(n6674) );
  NANDN U6951 ( .A(n6672), .B(n6671), .Z(n6673) );
  NAND U6952 ( .A(n6674), .B(n6673), .Z(n6833) );
  XNOR U6953 ( .A(n6832), .B(n6833), .Z(n6776) );
  XNOR U6954 ( .A(n6777), .B(n6776), .Z(n6779) );
  NANDN U6955 ( .A(n6676), .B(n6675), .Z(n6680) );
  NANDN U6956 ( .A(n6678), .B(n6677), .Z(n6679) );
  AND U6957 ( .A(n6680), .B(n6679), .Z(n6778) );
  XOR U6958 ( .A(n6779), .B(n6778), .Z(n6893) );
  NANDN U6959 ( .A(n6682), .B(n6681), .Z(n6686) );
  NANDN U6960 ( .A(n6684), .B(n6683), .Z(n6685) );
  AND U6961 ( .A(n6686), .B(n6685), .Z(n6890) );
  NANDN U6962 ( .A(n6688), .B(n6687), .Z(n6692) );
  NANDN U6963 ( .A(n6690), .B(n6689), .Z(n6691) );
  AND U6964 ( .A(n6692), .B(n6691), .Z(n6773) );
  NANDN U6965 ( .A(n6694), .B(n6693), .Z(n6698) );
  OR U6966 ( .A(n6696), .B(n6695), .Z(n6697) );
  AND U6967 ( .A(n6698), .B(n6697), .Z(n6771) );
  NANDN U6968 ( .A(n6700), .B(n6699), .Z(n6704) );
  NANDN U6969 ( .A(n6702), .B(n6701), .Z(n6703) );
  AND U6970 ( .A(n6704), .B(n6703), .Z(n6837) );
  NANDN U6971 ( .A(n6706), .B(n6705), .Z(n6710) );
  NANDN U6972 ( .A(n6708), .B(n6707), .Z(n6709) );
  NAND U6973 ( .A(n6710), .B(n6709), .Z(n6836) );
  XNOR U6974 ( .A(n6837), .B(n6836), .Z(n6838) );
  NAND U6975 ( .A(b[0]), .B(a[60]), .Z(n6711) );
  XNOR U6976 ( .A(b[1]), .B(n6711), .Z(n6713) );
  NANDN U6977 ( .A(b[0]), .B(a[59]), .Z(n6712) );
  NAND U6978 ( .A(n6713), .B(n6712), .Z(n6785) );
  NANDN U6979 ( .A(n19394), .B(n6714), .Z(n6716) );
  XOR U6980 ( .A(b[29]), .B(a[32]), .Z(n6863) );
  NANDN U6981 ( .A(n19395), .B(n6863), .Z(n6715) );
  AND U6982 ( .A(n6716), .B(n6715), .Z(n6783) );
  AND U6983 ( .A(b[31]), .B(a[28]), .Z(n6782) );
  XNOR U6984 ( .A(n6783), .B(n6782), .Z(n6784) );
  XNOR U6985 ( .A(n6785), .B(n6784), .Z(n6824) );
  NANDN U6986 ( .A(n19005), .B(n6717), .Z(n6719) );
  XOR U6987 ( .A(b[23]), .B(a[38]), .Z(n6866) );
  NANDN U6988 ( .A(n19055), .B(n6866), .Z(n6718) );
  AND U6989 ( .A(n6719), .B(n6718), .Z(n6857) );
  NANDN U6990 ( .A(n17362), .B(n6720), .Z(n6722) );
  XOR U6991 ( .A(b[7]), .B(a[54]), .Z(n6869) );
  NANDN U6992 ( .A(n17522), .B(n6869), .Z(n6721) );
  AND U6993 ( .A(n6722), .B(n6721), .Z(n6855) );
  NANDN U6994 ( .A(n19116), .B(n6723), .Z(n6725) );
  XOR U6995 ( .A(b[25]), .B(a[36]), .Z(n6872) );
  NANDN U6996 ( .A(n19179), .B(n6872), .Z(n6724) );
  NAND U6997 ( .A(n6725), .B(n6724), .Z(n6854) );
  XNOR U6998 ( .A(n6855), .B(n6854), .Z(n6856) );
  XOR U6999 ( .A(n6857), .B(n6856), .Z(n6825) );
  XNOR U7000 ( .A(n6824), .B(n6825), .Z(n6826) );
  NANDN U7001 ( .A(n18113), .B(n6726), .Z(n6728) );
  XOR U7002 ( .A(b[13]), .B(a[48]), .Z(n6875) );
  NANDN U7003 ( .A(n18229), .B(n6875), .Z(n6727) );
  AND U7004 ( .A(n6728), .B(n6727), .Z(n6819) );
  NANDN U7005 ( .A(n17888), .B(n6729), .Z(n6731) );
  XOR U7006 ( .A(b[11]), .B(a[50]), .Z(n6878) );
  NANDN U7007 ( .A(n18025), .B(n6878), .Z(n6730) );
  NAND U7008 ( .A(n6731), .B(n6730), .Z(n6818) );
  XNOR U7009 ( .A(n6819), .B(n6818), .Z(n6820) );
  NANDN U7010 ( .A(n18487), .B(n6732), .Z(n6734) );
  XOR U7011 ( .A(b[15]), .B(a[46]), .Z(n6881) );
  NANDN U7012 ( .A(n18311), .B(n6881), .Z(n6733) );
  AND U7013 ( .A(n6734), .B(n6733), .Z(n6815) );
  NANDN U7014 ( .A(n18853), .B(n6735), .Z(n6737) );
  XOR U7015 ( .A(b[21]), .B(a[40]), .Z(n6884) );
  NANDN U7016 ( .A(n18926), .B(n6884), .Z(n6736) );
  AND U7017 ( .A(n6737), .B(n6736), .Z(n6813) );
  NANDN U7018 ( .A(n17613), .B(n6738), .Z(n6740) );
  XOR U7019 ( .A(b[9]), .B(a[52]), .Z(n6887) );
  NANDN U7020 ( .A(n17739), .B(n6887), .Z(n6739) );
  NAND U7021 ( .A(n6740), .B(n6739), .Z(n6812) );
  XNOR U7022 ( .A(n6813), .B(n6812), .Z(n6814) );
  XOR U7023 ( .A(n6815), .B(n6814), .Z(n6821) );
  XOR U7024 ( .A(n6820), .B(n6821), .Z(n6827) );
  XOR U7025 ( .A(n6826), .B(n6827), .Z(n6839) );
  XNOR U7026 ( .A(n6838), .B(n6839), .Z(n6770) );
  XNOR U7027 ( .A(n6771), .B(n6770), .Z(n6772) );
  XOR U7028 ( .A(n6773), .B(n6772), .Z(n6891) );
  XNOR U7029 ( .A(n6890), .B(n6891), .Z(n6892) );
  XNOR U7030 ( .A(n6893), .B(n6892), .Z(n6898) );
  XOR U7031 ( .A(n6899), .B(n6898), .Z(n6765) );
  NANDN U7032 ( .A(n6742), .B(n6741), .Z(n6746) );
  NANDN U7033 ( .A(n6744), .B(n6743), .Z(n6745) );
  AND U7034 ( .A(n6746), .B(n6745), .Z(n6764) );
  XNOR U7035 ( .A(n6765), .B(n6764), .Z(n6766) );
  NANDN U7036 ( .A(n6748), .B(n6747), .Z(n6752) );
  NAND U7037 ( .A(n6750), .B(n6749), .Z(n6751) );
  NAND U7038 ( .A(n6752), .B(n6751), .Z(n6767) );
  XNOR U7039 ( .A(n6766), .B(n6767), .Z(n6758) );
  XNOR U7040 ( .A(n6759), .B(n6758), .Z(n6760) );
  XNOR U7041 ( .A(n6761), .B(n6760), .Z(n6902) );
  XNOR U7042 ( .A(sreg[156]), .B(n6902), .Z(n6904) );
  NANDN U7043 ( .A(sreg[155]), .B(n6753), .Z(n6757) );
  NAND U7044 ( .A(n6755), .B(n6754), .Z(n6756) );
  NAND U7045 ( .A(n6757), .B(n6756), .Z(n6903) );
  XNOR U7046 ( .A(n6904), .B(n6903), .Z(c[156]) );
  NANDN U7047 ( .A(n6759), .B(n6758), .Z(n6763) );
  NANDN U7048 ( .A(n6761), .B(n6760), .Z(n6762) );
  AND U7049 ( .A(n6763), .B(n6762), .Z(n6910) );
  NANDN U7050 ( .A(n6765), .B(n6764), .Z(n6769) );
  NANDN U7051 ( .A(n6767), .B(n6766), .Z(n6768) );
  AND U7052 ( .A(n6769), .B(n6768), .Z(n6908) );
  NANDN U7053 ( .A(n6771), .B(n6770), .Z(n6775) );
  NANDN U7054 ( .A(n6773), .B(n6772), .Z(n6774) );
  AND U7055 ( .A(n6775), .B(n6774), .Z(n6920) );
  NANDN U7056 ( .A(n6777), .B(n6776), .Z(n6781) );
  NAND U7057 ( .A(n6779), .B(n6778), .Z(n6780) );
  AND U7058 ( .A(n6781), .B(n6780), .Z(n6919) );
  XNOR U7059 ( .A(n6920), .B(n6919), .Z(n6922) );
  NANDN U7060 ( .A(n6783), .B(n6782), .Z(n6787) );
  NANDN U7061 ( .A(n6785), .B(n6784), .Z(n6786) );
  AND U7062 ( .A(n6787), .B(n6786), .Z(n6999) );
  NANDN U7063 ( .A(n19237), .B(n6788), .Z(n6790) );
  XOR U7064 ( .A(b[27]), .B(a[35]), .Z(n6943) );
  NANDN U7065 ( .A(n19277), .B(n6943), .Z(n6789) );
  AND U7066 ( .A(n6790), .B(n6789), .Z(n7006) );
  NANDN U7067 ( .A(n17072), .B(n6791), .Z(n6793) );
  XOR U7068 ( .A(b[5]), .B(a[57]), .Z(n6946) );
  NANDN U7069 ( .A(n17223), .B(n6946), .Z(n6792) );
  AND U7070 ( .A(n6793), .B(n6792), .Z(n7004) );
  NANDN U7071 ( .A(n18673), .B(n6794), .Z(n6796) );
  XOR U7072 ( .A(b[19]), .B(a[43]), .Z(n6949) );
  NANDN U7073 ( .A(n18758), .B(n6949), .Z(n6795) );
  NAND U7074 ( .A(n6796), .B(n6795), .Z(n7003) );
  XNOR U7075 ( .A(n7004), .B(n7003), .Z(n7005) );
  XNOR U7076 ( .A(n7006), .B(n7005), .Z(n6997) );
  NANDN U7077 ( .A(n19425), .B(n6797), .Z(n6799) );
  XOR U7078 ( .A(b[31]), .B(a[31]), .Z(n6952) );
  NANDN U7079 ( .A(n19426), .B(n6952), .Z(n6798) );
  AND U7080 ( .A(n6799), .B(n6798), .Z(n6964) );
  NANDN U7081 ( .A(n17067), .B(n6800), .Z(n6802) );
  XOR U7082 ( .A(b[3]), .B(a[59]), .Z(n6955) );
  NANDN U7083 ( .A(n17068), .B(n6955), .Z(n6801) );
  AND U7084 ( .A(n6802), .B(n6801), .Z(n6962) );
  NANDN U7085 ( .A(n18514), .B(n6803), .Z(n6805) );
  XOR U7086 ( .A(b[17]), .B(a[45]), .Z(n6958) );
  NANDN U7087 ( .A(n18585), .B(n6958), .Z(n6804) );
  NAND U7088 ( .A(n6805), .B(n6804), .Z(n6961) );
  XNOR U7089 ( .A(n6962), .B(n6961), .Z(n6963) );
  XOR U7090 ( .A(n6964), .B(n6963), .Z(n6998) );
  XOR U7091 ( .A(n6997), .B(n6998), .Z(n7000) );
  XOR U7092 ( .A(n6999), .B(n7000), .Z(n6932) );
  NANDN U7093 ( .A(n6807), .B(n6806), .Z(n6811) );
  NANDN U7094 ( .A(n6809), .B(n6808), .Z(n6810) );
  AND U7095 ( .A(n6811), .B(n6810), .Z(n6985) );
  NANDN U7096 ( .A(n6813), .B(n6812), .Z(n6817) );
  NANDN U7097 ( .A(n6815), .B(n6814), .Z(n6816) );
  NAND U7098 ( .A(n6817), .B(n6816), .Z(n6986) );
  XNOR U7099 ( .A(n6985), .B(n6986), .Z(n6987) );
  NANDN U7100 ( .A(n6819), .B(n6818), .Z(n6823) );
  NANDN U7101 ( .A(n6821), .B(n6820), .Z(n6822) );
  NAND U7102 ( .A(n6823), .B(n6822), .Z(n6988) );
  XNOR U7103 ( .A(n6987), .B(n6988), .Z(n6931) );
  XNOR U7104 ( .A(n6932), .B(n6931), .Z(n6934) );
  NANDN U7105 ( .A(n6825), .B(n6824), .Z(n6829) );
  NANDN U7106 ( .A(n6827), .B(n6826), .Z(n6828) );
  AND U7107 ( .A(n6829), .B(n6828), .Z(n6933) );
  XOR U7108 ( .A(n6934), .B(n6933), .Z(n7048) );
  NANDN U7109 ( .A(n6831), .B(n6830), .Z(n6835) );
  NANDN U7110 ( .A(n6833), .B(n6832), .Z(n6834) );
  AND U7111 ( .A(n6835), .B(n6834), .Z(n7045) );
  NANDN U7112 ( .A(n6837), .B(n6836), .Z(n6841) );
  NANDN U7113 ( .A(n6839), .B(n6838), .Z(n6840) );
  AND U7114 ( .A(n6841), .B(n6840), .Z(n6928) );
  NANDN U7115 ( .A(n6843), .B(n6842), .Z(n6847) );
  OR U7116 ( .A(n6845), .B(n6844), .Z(n6846) );
  AND U7117 ( .A(n6847), .B(n6846), .Z(n6926) );
  NANDN U7118 ( .A(n6849), .B(n6848), .Z(n6853) );
  NANDN U7119 ( .A(n6851), .B(n6850), .Z(n6852) );
  AND U7120 ( .A(n6853), .B(n6852), .Z(n6992) );
  NANDN U7121 ( .A(n6855), .B(n6854), .Z(n6859) );
  NANDN U7122 ( .A(n6857), .B(n6856), .Z(n6858) );
  NAND U7123 ( .A(n6859), .B(n6858), .Z(n6991) );
  XNOR U7124 ( .A(n6992), .B(n6991), .Z(n6993) );
  NAND U7125 ( .A(b[0]), .B(a[61]), .Z(n6860) );
  XNOR U7126 ( .A(b[1]), .B(n6860), .Z(n6862) );
  NANDN U7127 ( .A(b[0]), .B(a[60]), .Z(n6861) );
  NAND U7128 ( .A(n6862), .B(n6861), .Z(n6940) );
  NANDN U7129 ( .A(n19394), .B(n6863), .Z(n6865) );
  XOR U7130 ( .A(b[29]), .B(a[33]), .Z(n7018) );
  NANDN U7131 ( .A(n19395), .B(n7018), .Z(n6864) );
  AND U7132 ( .A(n6865), .B(n6864), .Z(n6938) );
  AND U7133 ( .A(b[31]), .B(a[29]), .Z(n6937) );
  XNOR U7134 ( .A(n6938), .B(n6937), .Z(n6939) );
  XNOR U7135 ( .A(n6940), .B(n6939), .Z(n6979) );
  NANDN U7136 ( .A(n19005), .B(n6866), .Z(n6868) );
  XOR U7137 ( .A(b[23]), .B(a[39]), .Z(n7021) );
  NANDN U7138 ( .A(n19055), .B(n7021), .Z(n6867) );
  AND U7139 ( .A(n6868), .B(n6867), .Z(n7012) );
  NANDN U7140 ( .A(n17362), .B(n6869), .Z(n6871) );
  XOR U7141 ( .A(b[7]), .B(a[55]), .Z(n7024) );
  NANDN U7142 ( .A(n17522), .B(n7024), .Z(n6870) );
  AND U7143 ( .A(n6871), .B(n6870), .Z(n7010) );
  NANDN U7144 ( .A(n19116), .B(n6872), .Z(n6874) );
  XOR U7145 ( .A(b[25]), .B(a[37]), .Z(n7027) );
  NANDN U7146 ( .A(n19179), .B(n7027), .Z(n6873) );
  NAND U7147 ( .A(n6874), .B(n6873), .Z(n7009) );
  XNOR U7148 ( .A(n7010), .B(n7009), .Z(n7011) );
  XOR U7149 ( .A(n7012), .B(n7011), .Z(n6980) );
  XNOR U7150 ( .A(n6979), .B(n6980), .Z(n6981) );
  NANDN U7151 ( .A(n18113), .B(n6875), .Z(n6877) );
  XOR U7152 ( .A(b[13]), .B(a[49]), .Z(n7030) );
  NANDN U7153 ( .A(n18229), .B(n7030), .Z(n6876) );
  AND U7154 ( .A(n6877), .B(n6876), .Z(n6974) );
  NANDN U7155 ( .A(n17888), .B(n6878), .Z(n6880) );
  XOR U7156 ( .A(b[11]), .B(a[51]), .Z(n7033) );
  NANDN U7157 ( .A(n18025), .B(n7033), .Z(n6879) );
  NAND U7158 ( .A(n6880), .B(n6879), .Z(n6973) );
  XNOR U7159 ( .A(n6974), .B(n6973), .Z(n6975) );
  NANDN U7160 ( .A(n18487), .B(n6881), .Z(n6883) );
  XOR U7161 ( .A(b[15]), .B(a[47]), .Z(n7036) );
  NANDN U7162 ( .A(n18311), .B(n7036), .Z(n6882) );
  AND U7163 ( .A(n6883), .B(n6882), .Z(n6970) );
  NANDN U7164 ( .A(n18853), .B(n6884), .Z(n6886) );
  XOR U7165 ( .A(b[21]), .B(a[41]), .Z(n7039) );
  NANDN U7166 ( .A(n18926), .B(n7039), .Z(n6885) );
  AND U7167 ( .A(n6886), .B(n6885), .Z(n6968) );
  NANDN U7168 ( .A(n17613), .B(n6887), .Z(n6889) );
  XOR U7169 ( .A(b[9]), .B(a[53]), .Z(n7042) );
  NANDN U7170 ( .A(n17739), .B(n7042), .Z(n6888) );
  NAND U7171 ( .A(n6889), .B(n6888), .Z(n6967) );
  XNOR U7172 ( .A(n6968), .B(n6967), .Z(n6969) );
  XOR U7173 ( .A(n6970), .B(n6969), .Z(n6976) );
  XOR U7174 ( .A(n6975), .B(n6976), .Z(n6982) );
  XOR U7175 ( .A(n6981), .B(n6982), .Z(n6994) );
  XNOR U7176 ( .A(n6993), .B(n6994), .Z(n6925) );
  XNOR U7177 ( .A(n6926), .B(n6925), .Z(n6927) );
  XOR U7178 ( .A(n6928), .B(n6927), .Z(n7046) );
  XNOR U7179 ( .A(n7045), .B(n7046), .Z(n7047) );
  XNOR U7180 ( .A(n7048), .B(n7047), .Z(n6921) );
  XOR U7181 ( .A(n6922), .B(n6921), .Z(n6914) );
  NANDN U7182 ( .A(n6891), .B(n6890), .Z(n6895) );
  NANDN U7183 ( .A(n6893), .B(n6892), .Z(n6894) );
  AND U7184 ( .A(n6895), .B(n6894), .Z(n6913) );
  XNOR U7185 ( .A(n6914), .B(n6913), .Z(n6915) );
  NANDN U7186 ( .A(n6897), .B(n6896), .Z(n6901) );
  NAND U7187 ( .A(n6899), .B(n6898), .Z(n6900) );
  NAND U7188 ( .A(n6901), .B(n6900), .Z(n6916) );
  XNOR U7189 ( .A(n6915), .B(n6916), .Z(n6907) );
  XNOR U7190 ( .A(n6908), .B(n6907), .Z(n6909) );
  XNOR U7191 ( .A(n6910), .B(n6909), .Z(n7051) );
  XNOR U7192 ( .A(sreg[157]), .B(n7051), .Z(n7053) );
  NANDN U7193 ( .A(sreg[156]), .B(n6902), .Z(n6906) );
  NAND U7194 ( .A(n6904), .B(n6903), .Z(n6905) );
  NAND U7195 ( .A(n6906), .B(n6905), .Z(n7052) );
  XNOR U7196 ( .A(n7053), .B(n7052), .Z(c[157]) );
  NANDN U7197 ( .A(n6908), .B(n6907), .Z(n6912) );
  NANDN U7198 ( .A(n6910), .B(n6909), .Z(n6911) );
  AND U7199 ( .A(n6912), .B(n6911), .Z(n7059) );
  NANDN U7200 ( .A(n6914), .B(n6913), .Z(n6918) );
  NANDN U7201 ( .A(n6916), .B(n6915), .Z(n6917) );
  AND U7202 ( .A(n6918), .B(n6917), .Z(n7057) );
  NANDN U7203 ( .A(n6920), .B(n6919), .Z(n6924) );
  NAND U7204 ( .A(n6922), .B(n6921), .Z(n6923) );
  AND U7205 ( .A(n6924), .B(n6923), .Z(n7064) );
  NANDN U7206 ( .A(n6926), .B(n6925), .Z(n6930) );
  NANDN U7207 ( .A(n6928), .B(n6927), .Z(n6929) );
  AND U7208 ( .A(n6930), .B(n6929), .Z(n7069) );
  NANDN U7209 ( .A(n6932), .B(n6931), .Z(n6936) );
  NAND U7210 ( .A(n6934), .B(n6933), .Z(n6935) );
  AND U7211 ( .A(n6936), .B(n6935), .Z(n7068) );
  XNOR U7212 ( .A(n7069), .B(n7068), .Z(n7071) );
  NANDN U7213 ( .A(n6938), .B(n6937), .Z(n6942) );
  NANDN U7214 ( .A(n6940), .B(n6939), .Z(n6941) );
  AND U7215 ( .A(n6942), .B(n6941), .Z(n7148) );
  NANDN U7216 ( .A(n19237), .B(n6943), .Z(n6945) );
  XOR U7217 ( .A(b[27]), .B(a[36]), .Z(n7092) );
  NANDN U7218 ( .A(n19277), .B(n7092), .Z(n6944) );
  AND U7219 ( .A(n6945), .B(n6944), .Z(n7155) );
  NANDN U7220 ( .A(n17072), .B(n6946), .Z(n6948) );
  XOR U7221 ( .A(b[5]), .B(a[58]), .Z(n7095) );
  NANDN U7222 ( .A(n17223), .B(n7095), .Z(n6947) );
  AND U7223 ( .A(n6948), .B(n6947), .Z(n7153) );
  NANDN U7224 ( .A(n18673), .B(n6949), .Z(n6951) );
  XOR U7225 ( .A(b[19]), .B(a[44]), .Z(n7098) );
  NANDN U7226 ( .A(n18758), .B(n7098), .Z(n6950) );
  NAND U7227 ( .A(n6951), .B(n6950), .Z(n7152) );
  XNOR U7228 ( .A(n7153), .B(n7152), .Z(n7154) );
  XNOR U7229 ( .A(n7155), .B(n7154), .Z(n7146) );
  NANDN U7230 ( .A(n19425), .B(n6952), .Z(n6954) );
  XOR U7231 ( .A(b[31]), .B(a[32]), .Z(n7101) );
  NANDN U7232 ( .A(n19426), .B(n7101), .Z(n6953) );
  AND U7233 ( .A(n6954), .B(n6953), .Z(n7113) );
  NANDN U7234 ( .A(n17067), .B(n6955), .Z(n6957) );
  XOR U7235 ( .A(b[3]), .B(a[60]), .Z(n7104) );
  NANDN U7236 ( .A(n17068), .B(n7104), .Z(n6956) );
  AND U7237 ( .A(n6957), .B(n6956), .Z(n7111) );
  NANDN U7238 ( .A(n18514), .B(n6958), .Z(n6960) );
  XOR U7239 ( .A(b[17]), .B(a[46]), .Z(n7107) );
  NANDN U7240 ( .A(n18585), .B(n7107), .Z(n6959) );
  NAND U7241 ( .A(n6960), .B(n6959), .Z(n7110) );
  XNOR U7242 ( .A(n7111), .B(n7110), .Z(n7112) );
  XOR U7243 ( .A(n7113), .B(n7112), .Z(n7147) );
  XOR U7244 ( .A(n7146), .B(n7147), .Z(n7149) );
  XOR U7245 ( .A(n7148), .B(n7149), .Z(n7081) );
  NANDN U7246 ( .A(n6962), .B(n6961), .Z(n6966) );
  NANDN U7247 ( .A(n6964), .B(n6963), .Z(n6965) );
  AND U7248 ( .A(n6966), .B(n6965), .Z(n7134) );
  NANDN U7249 ( .A(n6968), .B(n6967), .Z(n6972) );
  NANDN U7250 ( .A(n6970), .B(n6969), .Z(n6971) );
  NAND U7251 ( .A(n6972), .B(n6971), .Z(n7135) );
  XNOR U7252 ( .A(n7134), .B(n7135), .Z(n7136) );
  NANDN U7253 ( .A(n6974), .B(n6973), .Z(n6978) );
  NANDN U7254 ( .A(n6976), .B(n6975), .Z(n6977) );
  NAND U7255 ( .A(n6978), .B(n6977), .Z(n7137) );
  XNOR U7256 ( .A(n7136), .B(n7137), .Z(n7080) );
  XNOR U7257 ( .A(n7081), .B(n7080), .Z(n7083) );
  NANDN U7258 ( .A(n6980), .B(n6979), .Z(n6984) );
  NANDN U7259 ( .A(n6982), .B(n6981), .Z(n6983) );
  AND U7260 ( .A(n6984), .B(n6983), .Z(n7082) );
  XOR U7261 ( .A(n7083), .B(n7082), .Z(n7197) );
  NANDN U7262 ( .A(n6986), .B(n6985), .Z(n6990) );
  NANDN U7263 ( .A(n6988), .B(n6987), .Z(n6989) );
  AND U7264 ( .A(n6990), .B(n6989), .Z(n7194) );
  NANDN U7265 ( .A(n6992), .B(n6991), .Z(n6996) );
  NANDN U7266 ( .A(n6994), .B(n6993), .Z(n6995) );
  AND U7267 ( .A(n6996), .B(n6995), .Z(n7077) );
  NANDN U7268 ( .A(n6998), .B(n6997), .Z(n7002) );
  OR U7269 ( .A(n7000), .B(n6999), .Z(n7001) );
  AND U7270 ( .A(n7002), .B(n7001), .Z(n7075) );
  NANDN U7271 ( .A(n7004), .B(n7003), .Z(n7008) );
  NANDN U7272 ( .A(n7006), .B(n7005), .Z(n7007) );
  AND U7273 ( .A(n7008), .B(n7007), .Z(n7141) );
  NANDN U7274 ( .A(n7010), .B(n7009), .Z(n7014) );
  NANDN U7275 ( .A(n7012), .B(n7011), .Z(n7013) );
  NAND U7276 ( .A(n7014), .B(n7013), .Z(n7140) );
  XNOR U7277 ( .A(n7141), .B(n7140), .Z(n7142) );
  NAND U7278 ( .A(b[0]), .B(a[62]), .Z(n7015) );
  XNOR U7279 ( .A(b[1]), .B(n7015), .Z(n7017) );
  NANDN U7280 ( .A(b[0]), .B(a[61]), .Z(n7016) );
  NAND U7281 ( .A(n7017), .B(n7016), .Z(n7089) );
  NANDN U7282 ( .A(n19394), .B(n7018), .Z(n7020) );
  XOR U7283 ( .A(b[29]), .B(a[34]), .Z(n7167) );
  NANDN U7284 ( .A(n19395), .B(n7167), .Z(n7019) );
  AND U7285 ( .A(n7020), .B(n7019), .Z(n7087) );
  AND U7286 ( .A(b[31]), .B(a[30]), .Z(n7086) );
  XNOR U7287 ( .A(n7087), .B(n7086), .Z(n7088) );
  XNOR U7288 ( .A(n7089), .B(n7088), .Z(n7128) );
  NANDN U7289 ( .A(n19005), .B(n7021), .Z(n7023) );
  XOR U7290 ( .A(b[23]), .B(a[40]), .Z(n7170) );
  NANDN U7291 ( .A(n19055), .B(n7170), .Z(n7022) );
  AND U7292 ( .A(n7023), .B(n7022), .Z(n7161) );
  NANDN U7293 ( .A(n17362), .B(n7024), .Z(n7026) );
  XOR U7294 ( .A(b[7]), .B(a[56]), .Z(n7173) );
  NANDN U7295 ( .A(n17522), .B(n7173), .Z(n7025) );
  AND U7296 ( .A(n7026), .B(n7025), .Z(n7159) );
  NANDN U7297 ( .A(n19116), .B(n7027), .Z(n7029) );
  XOR U7298 ( .A(b[25]), .B(a[38]), .Z(n7176) );
  NANDN U7299 ( .A(n19179), .B(n7176), .Z(n7028) );
  NAND U7300 ( .A(n7029), .B(n7028), .Z(n7158) );
  XNOR U7301 ( .A(n7159), .B(n7158), .Z(n7160) );
  XOR U7302 ( .A(n7161), .B(n7160), .Z(n7129) );
  XNOR U7303 ( .A(n7128), .B(n7129), .Z(n7130) );
  NANDN U7304 ( .A(n18113), .B(n7030), .Z(n7032) );
  XOR U7305 ( .A(b[13]), .B(a[50]), .Z(n7179) );
  NANDN U7306 ( .A(n18229), .B(n7179), .Z(n7031) );
  AND U7307 ( .A(n7032), .B(n7031), .Z(n7123) );
  NANDN U7308 ( .A(n17888), .B(n7033), .Z(n7035) );
  XOR U7309 ( .A(b[11]), .B(a[52]), .Z(n7182) );
  NANDN U7310 ( .A(n18025), .B(n7182), .Z(n7034) );
  NAND U7311 ( .A(n7035), .B(n7034), .Z(n7122) );
  XNOR U7312 ( .A(n7123), .B(n7122), .Z(n7124) );
  NANDN U7313 ( .A(n18487), .B(n7036), .Z(n7038) );
  XOR U7314 ( .A(b[15]), .B(a[48]), .Z(n7185) );
  NANDN U7315 ( .A(n18311), .B(n7185), .Z(n7037) );
  AND U7316 ( .A(n7038), .B(n7037), .Z(n7119) );
  NANDN U7317 ( .A(n18853), .B(n7039), .Z(n7041) );
  XOR U7318 ( .A(b[21]), .B(a[42]), .Z(n7188) );
  NANDN U7319 ( .A(n18926), .B(n7188), .Z(n7040) );
  AND U7320 ( .A(n7041), .B(n7040), .Z(n7117) );
  NANDN U7321 ( .A(n17613), .B(n7042), .Z(n7044) );
  XOR U7322 ( .A(b[9]), .B(a[54]), .Z(n7191) );
  NANDN U7323 ( .A(n17739), .B(n7191), .Z(n7043) );
  NAND U7324 ( .A(n7044), .B(n7043), .Z(n7116) );
  XNOR U7325 ( .A(n7117), .B(n7116), .Z(n7118) );
  XOR U7326 ( .A(n7119), .B(n7118), .Z(n7125) );
  XOR U7327 ( .A(n7124), .B(n7125), .Z(n7131) );
  XOR U7328 ( .A(n7130), .B(n7131), .Z(n7143) );
  XNOR U7329 ( .A(n7142), .B(n7143), .Z(n7074) );
  XNOR U7330 ( .A(n7075), .B(n7074), .Z(n7076) );
  XOR U7331 ( .A(n7077), .B(n7076), .Z(n7195) );
  XNOR U7332 ( .A(n7194), .B(n7195), .Z(n7196) );
  XNOR U7333 ( .A(n7197), .B(n7196), .Z(n7070) );
  XOR U7334 ( .A(n7071), .B(n7070), .Z(n7063) );
  NANDN U7335 ( .A(n7046), .B(n7045), .Z(n7050) );
  NANDN U7336 ( .A(n7048), .B(n7047), .Z(n7049) );
  AND U7337 ( .A(n7050), .B(n7049), .Z(n7062) );
  XOR U7338 ( .A(n7063), .B(n7062), .Z(n7065) );
  XNOR U7339 ( .A(n7064), .B(n7065), .Z(n7056) );
  XNOR U7340 ( .A(n7057), .B(n7056), .Z(n7058) );
  XNOR U7341 ( .A(n7059), .B(n7058), .Z(n7200) );
  XNOR U7342 ( .A(sreg[158]), .B(n7200), .Z(n7202) );
  NANDN U7343 ( .A(sreg[157]), .B(n7051), .Z(n7055) );
  NAND U7344 ( .A(n7053), .B(n7052), .Z(n7054) );
  NAND U7345 ( .A(n7055), .B(n7054), .Z(n7201) );
  XNOR U7346 ( .A(n7202), .B(n7201), .Z(c[158]) );
  NANDN U7347 ( .A(n7057), .B(n7056), .Z(n7061) );
  NANDN U7348 ( .A(n7059), .B(n7058), .Z(n7060) );
  AND U7349 ( .A(n7061), .B(n7060), .Z(n7208) );
  NANDN U7350 ( .A(n7063), .B(n7062), .Z(n7067) );
  NANDN U7351 ( .A(n7065), .B(n7064), .Z(n7066) );
  AND U7352 ( .A(n7067), .B(n7066), .Z(n7206) );
  NANDN U7353 ( .A(n7069), .B(n7068), .Z(n7073) );
  NAND U7354 ( .A(n7071), .B(n7070), .Z(n7072) );
  AND U7355 ( .A(n7073), .B(n7072), .Z(n7213) );
  NANDN U7356 ( .A(n7075), .B(n7074), .Z(n7079) );
  NANDN U7357 ( .A(n7077), .B(n7076), .Z(n7078) );
  AND U7358 ( .A(n7079), .B(n7078), .Z(n7218) );
  NANDN U7359 ( .A(n7081), .B(n7080), .Z(n7085) );
  NAND U7360 ( .A(n7083), .B(n7082), .Z(n7084) );
  AND U7361 ( .A(n7085), .B(n7084), .Z(n7217) );
  XNOR U7362 ( .A(n7218), .B(n7217), .Z(n7220) );
  NANDN U7363 ( .A(n7087), .B(n7086), .Z(n7091) );
  NANDN U7364 ( .A(n7089), .B(n7088), .Z(n7090) );
  AND U7365 ( .A(n7091), .B(n7090), .Z(n7297) );
  NANDN U7366 ( .A(n19237), .B(n7092), .Z(n7094) );
  XOR U7367 ( .A(b[27]), .B(a[37]), .Z(n7241) );
  NANDN U7368 ( .A(n19277), .B(n7241), .Z(n7093) );
  AND U7369 ( .A(n7094), .B(n7093), .Z(n7304) );
  NANDN U7370 ( .A(n17072), .B(n7095), .Z(n7097) );
  XOR U7371 ( .A(b[5]), .B(a[59]), .Z(n7244) );
  NANDN U7372 ( .A(n17223), .B(n7244), .Z(n7096) );
  AND U7373 ( .A(n7097), .B(n7096), .Z(n7302) );
  NANDN U7374 ( .A(n18673), .B(n7098), .Z(n7100) );
  XOR U7375 ( .A(b[19]), .B(a[45]), .Z(n7247) );
  NANDN U7376 ( .A(n18758), .B(n7247), .Z(n7099) );
  NAND U7377 ( .A(n7100), .B(n7099), .Z(n7301) );
  XNOR U7378 ( .A(n7302), .B(n7301), .Z(n7303) );
  XNOR U7379 ( .A(n7304), .B(n7303), .Z(n7295) );
  NANDN U7380 ( .A(n19425), .B(n7101), .Z(n7103) );
  XOR U7381 ( .A(b[31]), .B(a[33]), .Z(n7250) );
  NANDN U7382 ( .A(n19426), .B(n7250), .Z(n7102) );
  AND U7383 ( .A(n7103), .B(n7102), .Z(n7262) );
  NANDN U7384 ( .A(n17067), .B(n7104), .Z(n7106) );
  XOR U7385 ( .A(b[3]), .B(a[61]), .Z(n7253) );
  NANDN U7386 ( .A(n17068), .B(n7253), .Z(n7105) );
  AND U7387 ( .A(n7106), .B(n7105), .Z(n7260) );
  NANDN U7388 ( .A(n18514), .B(n7107), .Z(n7109) );
  XOR U7389 ( .A(b[17]), .B(a[47]), .Z(n7256) );
  NANDN U7390 ( .A(n18585), .B(n7256), .Z(n7108) );
  NAND U7391 ( .A(n7109), .B(n7108), .Z(n7259) );
  XNOR U7392 ( .A(n7260), .B(n7259), .Z(n7261) );
  XOR U7393 ( .A(n7262), .B(n7261), .Z(n7296) );
  XOR U7394 ( .A(n7295), .B(n7296), .Z(n7298) );
  XOR U7395 ( .A(n7297), .B(n7298), .Z(n7230) );
  NANDN U7396 ( .A(n7111), .B(n7110), .Z(n7115) );
  NANDN U7397 ( .A(n7113), .B(n7112), .Z(n7114) );
  AND U7398 ( .A(n7115), .B(n7114), .Z(n7283) );
  NANDN U7399 ( .A(n7117), .B(n7116), .Z(n7121) );
  NANDN U7400 ( .A(n7119), .B(n7118), .Z(n7120) );
  NAND U7401 ( .A(n7121), .B(n7120), .Z(n7284) );
  XNOR U7402 ( .A(n7283), .B(n7284), .Z(n7285) );
  NANDN U7403 ( .A(n7123), .B(n7122), .Z(n7127) );
  NANDN U7404 ( .A(n7125), .B(n7124), .Z(n7126) );
  NAND U7405 ( .A(n7127), .B(n7126), .Z(n7286) );
  XNOR U7406 ( .A(n7285), .B(n7286), .Z(n7229) );
  XNOR U7407 ( .A(n7230), .B(n7229), .Z(n7232) );
  NANDN U7408 ( .A(n7129), .B(n7128), .Z(n7133) );
  NANDN U7409 ( .A(n7131), .B(n7130), .Z(n7132) );
  AND U7410 ( .A(n7133), .B(n7132), .Z(n7231) );
  XOR U7411 ( .A(n7232), .B(n7231), .Z(n7346) );
  NANDN U7412 ( .A(n7135), .B(n7134), .Z(n7139) );
  NANDN U7413 ( .A(n7137), .B(n7136), .Z(n7138) );
  AND U7414 ( .A(n7139), .B(n7138), .Z(n7343) );
  NANDN U7415 ( .A(n7141), .B(n7140), .Z(n7145) );
  NANDN U7416 ( .A(n7143), .B(n7142), .Z(n7144) );
  AND U7417 ( .A(n7145), .B(n7144), .Z(n7226) );
  NANDN U7418 ( .A(n7147), .B(n7146), .Z(n7151) );
  OR U7419 ( .A(n7149), .B(n7148), .Z(n7150) );
  AND U7420 ( .A(n7151), .B(n7150), .Z(n7224) );
  NANDN U7421 ( .A(n7153), .B(n7152), .Z(n7157) );
  NANDN U7422 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U7423 ( .A(n7157), .B(n7156), .Z(n7290) );
  NANDN U7424 ( .A(n7159), .B(n7158), .Z(n7163) );
  NANDN U7425 ( .A(n7161), .B(n7160), .Z(n7162) );
  NAND U7426 ( .A(n7163), .B(n7162), .Z(n7289) );
  XNOR U7427 ( .A(n7290), .B(n7289), .Z(n7291) );
  NAND U7428 ( .A(b[0]), .B(a[63]), .Z(n7164) );
  XNOR U7429 ( .A(b[1]), .B(n7164), .Z(n7166) );
  NANDN U7430 ( .A(b[0]), .B(a[62]), .Z(n7165) );
  NAND U7431 ( .A(n7166), .B(n7165), .Z(n7238) );
  NANDN U7432 ( .A(n19394), .B(n7167), .Z(n7169) );
  XOR U7433 ( .A(b[29]), .B(a[35]), .Z(n7316) );
  NANDN U7434 ( .A(n19395), .B(n7316), .Z(n7168) );
  AND U7435 ( .A(n7169), .B(n7168), .Z(n7236) );
  AND U7436 ( .A(b[31]), .B(a[31]), .Z(n7235) );
  XNOR U7437 ( .A(n7236), .B(n7235), .Z(n7237) );
  XNOR U7438 ( .A(n7238), .B(n7237), .Z(n7277) );
  NANDN U7439 ( .A(n19005), .B(n7170), .Z(n7172) );
  XOR U7440 ( .A(b[23]), .B(a[41]), .Z(n7319) );
  NANDN U7441 ( .A(n19055), .B(n7319), .Z(n7171) );
  AND U7442 ( .A(n7172), .B(n7171), .Z(n7310) );
  NANDN U7443 ( .A(n17362), .B(n7173), .Z(n7175) );
  XOR U7444 ( .A(b[7]), .B(a[57]), .Z(n7322) );
  NANDN U7445 ( .A(n17522), .B(n7322), .Z(n7174) );
  AND U7446 ( .A(n7175), .B(n7174), .Z(n7308) );
  NANDN U7447 ( .A(n19116), .B(n7176), .Z(n7178) );
  XOR U7448 ( .A(b[25]), .B(a[39]), .Z(n7325) );
  NANDN U7449 ( .A(n19179), .B(n7325), .Z(n7177) );
  NAND U7450 ( .A(n7178), .B(n7177), .Z(n7307) );
  XNOR U7451 ( .A(n7308), .B(n7307), .Z(n7309) );
  XOR U7452 ( .A(n7310), .B(n7309), .Z(n7278) );
  XNOR U7453 ( .A(n7277), .B(n7278), .Z(n7279) );
  NANDN U7454 ( .A(n18113), .B(n7179), .Z(n7181) );
  XOR U7455 ( .A(b[13]), .B(a[51]), .Z(n7328) );
  NANDN U7456 ( .A(n18229), .B(n7328), .Z(n7180) );
  AND U7457 ( .A(n7181), .B(n7180), .Z(n7272) );
  NANDN U7458 ( .A(n17888), .B(n7182), .Z(n7184) );
  XOR U7459 ( .A(b[11]), .B(a[53]), .Z(n7331) );
  NANDN U7460 ( .A(n18025), .B(n7331), .Z(n7183) );
  NAND U7461 ( .A(n7184), .B(n7183), .Z(n7271) );
  XNOR U7462 ( .A(n7272), .B(n7271), .Z(n7273) );
  NANDN U7463 ( .A(n18487), .B(n7185), .Z(n7187) );
  XOR U7464 ( .A(b[15]), .B(a[49]), .Z(n7334) );
  NANDN U7465 ( .A(n18311), .B(n7334), .Z(n7186) );
  AND U7466 ( .A(n7187), .B(n7186), .Z(n7268) );
  NANDN U7467 ( .A(n18853), .B(n7188), .Z(n7190) );
  XOR U7468 ( .A(b[21]), .B(a[43]), .Z(n7337) );
  NANDN U7469 ( .A(n18926), .B(n7337), .Z(n7189) );
  AND U7470 ( .A(n7190), .B(n7189), .Z(n7266) );
  NANDN U7471 ( .A(n17613), .B(n7191), .Z(n7193) );
  XOR U7472 ( .A(b[9]), .B(a[55]), .Z(n7340) );
  NANDN U7473 ( .A(n17739), .B(n7340), .Z(n7192) );
  NAND U7474 ( .A(n7193), .B(n7192), .Z(n7265) );
  XNOR U7475 ( .A(n7266), .B(n7265), .Z(n7267) );
  XOR U7476 ( .A(n7268), .B(n7267), .Z(n7274) );
  XOR U7477 ( .A(n7273), .B(n7274), .Z(n7280) );
  XOR U7478 ( .A(n7279), .B(n7280), .Z(n7292) );
  XNOR U7479 ( .A(n7291), .B(n7292), .Z(n7223) );
  XNOR U7480 ( .A(n7224), .B(n7223), .Z(n7225) );
  XOR U7481 ( .A(n7226), .B(n7225), .Z(n7344) );
  XNOR U7482 ( .A(n7343), .B(n7344), .Z(n7345) );
  XNOR U7483 ( .A(n7346), .B(n7345), .Z(n7219) );
  XOR U7484 ( .A(n7220), .B(n7219), .Z(n7212) );
  NANDN U7485 ( .A(n7195), .B(n7194), .Z(n7199) );
  NANDN U7486 ( .A(n7197), .B(n7196), .Z(n7198) );
  AND U7487 ( .A(n7199), .B(n7198), .Z(n7211) );
  XOR U7488 ( .A(n7212), .B(n7211), .Z(n7214) );
  XNOR U7489 ( .A(n7213), .B(n7214), .Z(n7205) );
  XNOR U7490 ( .A(n7206), .B(n7205), .Z(n7207) );
  XNOR U7491 ( .A(n7208), .B(n7207), .Z(n7349) );
  XNOR U7492 ( .A(sreg[159]), .B(n7349), .Z(n7351) );
  NANDN U7493 ( .A(sreg[158]), .B(n7200), .Z(n7204) );
  NAND U7494 ( .A(n7202), .B(n7201), .Z(n7203) );
  NAND U7495 ( .A(n7204), .B(n7203), .Z(n7350) );
  XNOR U7496 ( .A(n7351), .B(n7350), .Z(c[159]) );
  NANDN U7497 ( .A(n7206), .B(n7205), .Z(n7210) );
  NANDN U7498 ( .A(n7208), .B(n7207), .Z(n7209) );
  AND U7499 ( .A(n7210), .B(n7209), .Z(n7357) );
  NANDN U7500 ( .A(n7212), .B(n7211), .Z(n7216) );
  NANDN U7501 ( .A(n7214), .B(n7213), .Z(n7215) );
  AND U7502 ( .A(n7216), .B(n7215), .Z(n7355) );
  NANDN U7503 ( .A(n7218), .B(n7217), .Z(n7222) );
  NAND U7504 ( .A(n7220), .B(n7219), .Z(n7221) );
  AND U7505 ( .A(n7222), .B(n7221), .Z(n7362) );
  NANDN U7506 ( .A(n7224), .B(n7223), .Z(n7228) );
  NANDN U7507 ( .A(n7226), .B(n7225), .Z(n7227) );
  AND U7508 ( .A(n7228), .B(n7227), .Z(n7367) );
  NANDN U7509 ( .A(n7230), .B(n7229), .Z(n7234) );
  NAND U7510 ( .A(n7232), .B(n7231), .Z(n7233) );
  AND U7511 ( .A(n7234), .B(n7233), .Z(n7366) );
  XNOR U7512 ( .A(n7367), .B(n7366), .Z(n7369) );
  NANDN U7513 ( .A(n7236), .B(n7235), .Z(n7240) );
  NANDN U7514 ( .A(n7238), .B(n7237), .Z(n7239) );
  AND U7515 ( .A(n7240), .B(n7239), .Z(n7446) );
  NANDN U7516 ( .A(n19237), .B(n7241), .Z(n7243) );
  XOR U7517 ( .A(b[27]), .B(a[38]), .Z(n7390) );
  NANDN U7518 ( .A(n19277), .B(n7390), .Z(n7242) );
  AND U7519 ( .A(n7243), .B(n7242), .Z(n7453) );
  NANDN U7520 ( .A(n17072), .B(n7244), .Z(n7246) );
  XOR U7521 ( .A(b[5]), .B(a[60]), .Z(n7393) );
  NANDN U7522 ( .A(n17223), .B(n7393), .Z(n7245) );
  AND U7523 ( .A(n7246), .B(n7245), .Z(n7451) );
  NANDN U7524 ( .A(n18673), .B(n7247), .Z(n7249) );
  XOR U7525 ( .A(b[19]), .B(a[46]), .Z(n7396) );
  NANDN U7526 ( .A(n18758), .B(n7396), .Z(n7248) );
  NAND U7527 ( .A(n7249), .B(n7248), .Z(n7450) );
  XNOR U7528 ( .A(n7451), .B(n7450), .Z(n7452) );
  XNOR U7529 ( .A(n7453), .B(n7452), .Z(n7444) );
  NANDN U7530 ( .A(n19425), .B(n7250), .Z(n7252) );
  XOR U7531 ( .A(b[31]), .B(a[34]), .Z(n7399) );
  NANDN U7532 ( .A(n19426), .B(n7399), .Z(n7251) );
  AND U7533 ( .A(n7252), .B(n7251), .Z(n7411) );
  NANDN U7534 ( .A(n17067), .B(n7253), .Z(n7255) );
  XOR U7535 ( .A(b[3]), .B(a[62]), .Z(n7402) );
  NANDN U7536 ( .A(n17068), .B(n7402), .Z(n7254) );
  AND U7537 ( .A(n7255), .B(n7254), .Z(n7409) );
  NANDN U7538 ( .A(n18514), .B(n7256), .Z(n7258) );
  XOR U7539 ( .A(b[17]), .B(a[48]), .Z(n7405) );
  NANDN U7540 ( .A(n18585), .B(n7405), .Z(n7257) );
  NAND U7541 ( .A(n7258), .B(n7257), .Z(n7408) );
  XNOR U7542 ( .A(n7409), .B(n7408), .Z(n7410) );
  XOR U7543 ( .A(n7411), .B(n7410), .Z(n7445) );
  XOR U7544 ( .A(n7444), .B(n7445), .Z(n7447) );
  XOR U7545 ( .A(n7446), .B(n7447), .Z(n7379) );
  NANDN U7546 ( .A(n7260), .B(n7259), .Z(n7264) );
  NANDN U7547 ( .A(n7262), .B(n7261), .Z(n7263) );
  AND U7548 ( .A(n7264), .B(n7263), .Z(n7432) );
  NANDN U7549 ( .A(n7266), .B(n7265), .Z(n7270) );
  NANDN U7550 ( .A(n7268), .B(n7267), .Z(n7269) );
  NAND U7551 ( .A(n7270), .B(n7269), .Z(n7433) );
  XNOR U7552 ( .A(n7432), .B(n7433), .Z(n7434) );
  NANDN U7553 ( .A(n7272), .B(n7271), .Z(n7276) );
  NANDN U7554 ( .A(n7274), .B(n7273), .Z(n7275) );
  NAND U7555 ( .A(n7276), .B(n7275), .Z(n7435) );
  XNOR U7556 ( .A(n7434), .B(n7435), .Z(n7378) );
  XNOR U7557 ( .A(n7379), .B(n7378), .Z(n7381) );
  NANDN U7558 ( .A(n7278), .B(n7277), .Z(n7282) );
  NANDN U7559 ( .A(n7280), .B(n7279), .Z(n7281) );
  AND U7560 ( .A(n7282), .B(n7281), .Z(n7380) );
  XOR U7561 ( .A(n7381), .B(n7380), .Z(n7495) );
  NANDN U7562 ( .A(n7284), .B(n7283), .Z(n7288) );
  NANDN U7563 ( .A(n7286), .B(n7285), .Z(n7287) );
  AND U7564 ( .A(n7288), .B(n7287), .Z(n7492) );
  NANDN U7565 ( .A(n7290), .B(n7289), .Z(n7294) );
  NANDN U7566 ( .A(n7292), .B(n7291), .Z(n7293) );
  AND U7567 ( .A(n7294), .B(n7293), .Z(n7375) );
  NANDN U7568 ( .A(n7296), .B(n7295), .Z(n7300) );
  OR U7569 ( .A(n7298), .B(n7297), .Z(n7299) );
  AND U7570 ( .A(n7300), .B(n7299), .Z(n7373) );
  NANDN U7571 ( .A(n7302), .B(n7301), .Z(n7306) );
  NANDN U7572 ( .A(n7304), .B(n7303), .Z(n7305) );
  AND U7573 ( .A(n7306), .B(n7305), .Z(n7439) );
  NANDN U7574 ( .A(n7308), .B(n7307), .Z(n7312) );
  NANDN U7575 ( .A(n7310), .B(n7309), .Z(n7311) );
  NAND U7576 ( .A(n7312), .B(n7311), .Z(n7438) );
  XNOR U7577 ( .A(n7439), .B(n7438), .Z(n7440) );
  NAND U7578 ( .A(b[0]), .B(a[64]), .Z(n7313) );
  XNOR U7579 ( .A(b[1]), .B(n7313), .Z(n7315) );
  NANDN U7580 ( .A(b[0]), .B(a[63]), .Z(n7314) );
  NAND U7581 ( .A(n7315), .B(n7314), .Z(n7387) );
  NANDN U7582 ( .A(n19394), .B(n7316), .Z(n7318) );
  XOR U7583 ( .A(b[29]), .B(a[36]), .Z(n7465) );
  NANDN U7584 ( .A(n19395), .B(n7465), .Z(n7317) );
  AND U7585 ( .A(n7318), .B(n7317), .Z(n7385) );
  AND U7586 ( .A(b[31]), .B(a[32]), .Z(n7384) );
  XNOR U7587 ( .A(n7385), .B(n7384), .Z(n7386) );
  XNOR U7588 ( .A(n7387), .B(n7386), .Z(n7426) );
  NANDN U7589 ( .A(n19005), .B(n7319), .Z(n7321) );
  XOR U7590 ( .A(b[23]), .B(a[42]), .Z(n7468) );
  NANDN U7591 ( .A(n19055), .B(n7468), .Z(n7320) );
  AND U7592 ( .A(n7321), .B(n7320), .Z(n7459) );
  NANDN U7593 ( .A(n17362), .B(n7322), .Z(n7324) );
  XOR U7594 ( .A(b[7]), .B(a[58]), .Z(n7471) );
  NANDN U7595 ( .A(n17522), .B(n7471), .Z(n7323) );
  AND U7596 ( .A(n7324), .B(n7323), .Z(n7457) );
  NANDN U7597 ( .A(n19116), .B(n7325), .Z(n7327) );
  XOR U7598 ( .A(b[25]), .B(a[40]), .Z(n7474) );
  NANDN U7599 ( .A(n19179), .B(n7474), .Z(n7326) );
  NAND U7600 ( .A(n7327), .B(n7326), .Z(n7456) );
  XNOR U7601 ( .A(n7457), .B(n7456), .Z(n7458) );
  XOR U7602 ( .A(n7459), .B(n7458), .Z(n7427) );
  XNOR U7603 ( .A(n7426), .B(n7427), .Z(n7428) );
  NANDN U7604 ( .A(n18113), .B(n7328), .Z(n7330) );
  XOR U7605 ( .A(b[13]), .B(a[52]), .Z(n7477) );
  NANDN U7606 ( .A(n18229), .B(n7477), .Z(n7329) );
  AND U7607 ( .A(n7330), .B(n7329), .Z(n7421) );
  NANDN U7608 ( .A(n17888), .B(n7331), .Z(n7333) );
  XOR U7609 ( .A(b[11]), .B(a[54]), .Z(n7480) );
  NANDN U7610 ( .A(n18025), .B(n7480), .Z(n7332) );
  NAND U7611 ( .A(n7333), .B(n7332), .Z(n7420) );
  XNOR U7612 ( .A(n7421), .B(n7420), .Z(n7422) );
  NANDN U7613 ( .A(n18487), .B(n7334), .Z(n7336) );
  XOR U7614 ( .A(b[15]), .B(a[50]), .Z(n7483) );
  NANDN U7615 ( .A(n18311), .B(n7483), .Z(n7335) );
  AND U7616 ( .A(n7336), .B(n7335), .Z(n7417) );
  NANDN U7617 ( .A(n18853), .B(n7337), .Z(n7339) );
  XOR U7618 ( .A(b[21]), .B(a[44]), .Z(n7486) );
  NANDN U7619 ( .A(n18926), .B(n7486), .Z(n7338) );
  AND U7620 ( .A(n7339), .B(n7338), .Z(n7415) );
  NANDN U7621 ( .A(n17613), .B(n7340), .Z(n7342) );
  XOR U7622 ( .A(b[9]), .B(a[56]), .Z(n7489) );
  NANDN U7623 ( .A(n17739), .B(n7489), .Z(n7341) );
  NAND U7624 ( .A(n7342), .B(n7341), .Z(n7414) );
  XNOR U7625 ( .A(n7415), .B(n7414), .Z(n7416) );
  XOR U7626 ( .A(n7417), .B(n7416), .Z(n7423) );
  XOR U7627 ( .A(n7422), .B(n7423), .Z(n7429) );
  XOR U7628 ( .A(n7428), .B(n7429), .Z(n7441) );
  XNOR U7629 ( .A(n7440), .B(n7441), .Z(n7372) );
  XNOR U7630 ( .A(n7373), .B(n7372), .Z(n7374) );
  XOR U7631 ( .A(n7375), .B(n7374), .Z(n7493) );
  XNOR U7632 ( .A(n7492), .B(n7493), .Z(n7494) );
  XNOR U7633 ( .A(n7495), .B(n7494), .Z(n7368) );
  XOR U7634 ( .A(n7369), .B(n7368), .Z(n7361) );
  NANDN U7635 ( .A(n7344), .B(n7343), .Z(n7348) );
  NANDN U7636 ( .A(n7346), .B(n7345), .Z(n7347) );
  AND U7637 ( .A(n7348), .B(n7347), .Z(n7360) );
  XOR U7638 ( .A(n7361), .B(n7360), .Z(n7363) );
  XNOR U7639 ( .A(n7362), .B(n7363), .Z(n7354) );
  XNOR U7640 ( .A(n7355), .B(n7354), .Z(n7356) );
  XNOR U7641 ( .A(n7357), .B(n7356), .Z(n7498) );
  XNOR U7642 ( .A(sreg[160]), .B(n7498), .Z(n7500) );
  NANDN U7643 ( .A(sreg[159]), .B(n7349), .Z(n7353) );
  NAND U7644 ( .A(n7351), .B(n7350), .Z(n7352) );
  NAND U7645 ( .A(n7353), .B(n7352), .Z(n7499) );
  XNOR U7646 ( .A(n7500), .B(n7499), .Z(c[160]) );
  NANDN U7647 ( .A(n7355), .B(n7354), .Z(n7359) );
  NANDN U7648 ( .A(n7357), .B(n7356), .Z(n7358) );
  AND U7649 ( .A(n7359), .B(n7358), .Z(n7506) );
  NANDN U7650 ( .A(n7361), .B(n7360), .Z(n7365) );
  NANDN U7651 ( .A(n7363), .B(n7362), .Z(n7364) );
  AND U7652 ( .A(n7365), .B(n7364), .Z(n7504) );
  NANDN U7653 ( .A(n7367), .B(n7366), .Z(n7371) );
  NAND U7654 ( .A(n7369), .B(n7368), .Z(n7370) );
  AND U7655 ( .A(n7371), .B(n7370), .Z(n7511) );
  NANDN U7656 ( .A(n7373), .B(n7372), .Z(n7377) );
  NANDN U7657 ( .A(n7375), .B(n7374), .Z(n7376) );
  AND U7658 ( .A(n7377), .B(n7376), .Z(n7516) );
  NANDN U7659 ( .A(n7379), .B(n7378), .Z(n7383) );
  NAND U7660 ( .A(n7381), .B(n7380), .Z(n7382) );
  AND U7661 ( .A(n7383), .B(n7382), .Z(n7515) );
  XNOR U7662 ( .A(n7516), .B(n7515), .Z(n7518) );
  NANDN U7663 ( .A(n7385), .B(n7384), .Z(n7389) );
  NANDN U7664 ( .A(n7387), .B(n7386), .Z(n7388) );
  AND U7665 ( .A(n7389), .B(n7388), .Z(n7595) );
  NANDN U7666 ( .A(n19237), .B(n7390), .Z(n7392) );
  XOR U7667 ( .A(b[27]), .B(a[39]), .Z(n7539) );
  NANDN U7668 ( .A(n19277), .B(n7539), .Z(n7391) );
  AND U7669 ( .A(n7392), .B(n7391), .Z(n7602) );
  NANDN U7670 ( .A(n17072), .B(n7393), .Z(n7395) );
  XOR U7671 ( .A(b[5]), .B(a[61]), .Z(n7542) );
  NANDN U7672 ( .A(n17223), .B(n7542), .Z(n7394) );
  AND U7673 ( .A(n7395), .B(n7394), .Z(n7600) );
  NANDN U7674 ( .A(n18673), .B(n7396), .Z(n7398) );
  XOR U7675 ( .A(b[19]), .B(a[47]), .Z(n7545) );
  NANDN U7676 ( .A(n18758), .B(n7545), .Z(n7397) );
  NAND U7677 ( .A(n7398), .B(n7397), .Z(n7599) );
  XNOR U7678 ( .A(n7600), .B(n7599), .Z(n7601) );
  XNOR U7679 ( .A(n7602), .B(n7601), .Z(n7593) );
  NANDN U7680 ( .A(n19425), .B(n7399), .Z(n7401) );
  XOR U7681 ( .A(b[31]), .B(a[35]), .Z(n7548) );
  NANDN U7682 ( .A(n19426), .B(n7548), .Z(n7400) );
  AND U7683 ( .A(n7401), .B(n7400), .Z(n7560) );
  NANDN U7684 ( .A(n17067), .B(n7402), .Z(n7404) );
  XOR U7685 ( .A(b[3]), .B(a[63]), .Z(n7551) );
  NANDN U7686 ( .A(n17068), .B(n7551), .Z(n7403) );
  AND U7687 ( .A(n7404), .B(n7403), .Z(n7558) );
  NANDN U7688 ( .A(n18514), .B(n7405), .Z(n7407) );
  XOR U7689 ( .A(b[17]), .B(a[49]), .Z(n7554) );
  NANDN U7690 ( .A(n18585), .B(n7554), .Z(n7406) );
  NAND U7691 ( .A(n7407), .B(n7406), .Z(n7557) );
  XNOR U7692 ( .A(n7558), .B(n7557), .Z(n7559) );
  XOR U7693 ( .A(n7560), .B(n7559), .Z(n7594) );
  XOR U7694 ( .A(n7593), .B(n7594), .Z(n7596) );
  XOR U7695 ( .A(n7595), .B(n7596), .Z(n7528) );
  NANDN U7696 ( .A(n7409), .B(n7408), .Z(n7413) );
  NANDN U7697 ( .A(n7411), .B(n7410), .Z(n7412) );
  AND U7698 ( .A(n7413), .B(n7412), .Z(n7581) );
  NANDN U7699 ( .A(n7415), .B(n7414), .Z(n7419) );
  NANDN U7700 ( .A(n7417), .B(n7416), .Z(n7418) );
  NAND U7701 ( .A(n7419), .B(n7418), .Z(n7582) );
  XNOR U7702 ( .A(n7581), .B(n7582), .Z(n7583) );
  NANDN U7703 ( .A(n7421), .B(n7420), .Z(n7425) );
  NANDN U7704 ( .A(n7423), .B(n7422), .Z(n7424) );
  NAND U7705 ( .A(n7425), .B(n7424), .Z(n7584) );
  XNOR U7706 ( .A(n7583), .B(n7584), .Z(n7527) );
  XNOR U7707 ( .A(n7528), .B(n7527), .Z(n7530) );
  NANDN U7708 ( .A(n7427), .B(n7426), .Z(n7431) );
  NANDN U7709 ( .A(n7429), .B(n7428), .Z(n7430) );
  AND U7710 ( .A(n7431), .B(n7430), .Z(n7529) );
  XOR U7711 ( .A(n7530), .B(n7529), .Z(n7644) );
  NANDN U7712 ( .A(n7433), .B(n7432), .Z(n7437) );
  NANDN U7713 ( .A(n7435), .B(n7434), .Z(n7436) );
  AND U7714 ( .A(n7437), .B(n7436), .Z(n7641) );
  NANDN U7715 ( .A(n7439), .B(n7438), .Z(n7443) );
  NANDN U7716 ( .A(n7441), .B(n7440), .Z(n7442) );
  AND U7717 ( .A(n7443), .B(n7442), .Z(n7524) );
  NANDN U7718 ( .A(n7445), .B(n7444), .Z(n7449) );
  OR U7719 ( .A(n7447), .B(n7446), .Z(n7448) );
  AND U7720 ( .A(n7449), .B(n7448), .Z(n7522) );
  NANDN U7721 ( .A(n7451), .B(n7450), .Z(n7455) );
  NANDN U7722 ( .A(n7453), .B(n7452), .Z(n7454) );
  AND U7723 ( .A(n7455), .B(n7454), .Z(n7588) );
  NANDN U7724 ( .A(n7457), .B(n7456), .Z(n7461) );
  NANDN U7725 ( .A(n7459), .B(n7458), .Z(n7460) );
  NAND U7726 ( .A(n7461), .B(n7460), .Z(n7587) );
  XNOR U7727 ( .A(n7588), .B(n7587), .Z(n7589) );
  NAND U7728 ( .A(b[0]), .B(a[65]), .Z(n7462) );
  XNOR U7729 ( .A(b[1]), .B(n7462), .Z(n7464) );
  NANDN U7730 ( .A(b[0]), .B(a[64]), .Z(n7463) );
  NAND U7731 ( .A(n7464), .B(n7463), .Z(n7536) );
  NANDN U7732 ( .A(n19394), .B(n7465), .Z(n7467) );
  XOR U7733 ( .A(b[29]), .B(a[37]), .Z(n7611) );
  NANDN U7734 ( .A(n19395), .B(n7611), .Z(n7466) );
  AND U7735 ( .A(n7467), .B(n7466), .Z(n7534) );
  AND U7736 ( .A(b[31]), .B(a[33]), .Z(n7533) );
  XNOR U7737 ( .A(n7534), .B(n7533), .Z(n7535) );
  XNOR U7738 ( .A(n7536), .B(n7535), .Z(n7575) );
  NANDN U7739 ( .A(n19005), .B(n7468), .Z(n7470) );
  XOR U7740 ( .A(b[23]), .B(a[43]), .Z(n7617) );
  NANDN U7741 ( .A(n19055), .B(n7617), .Z(n7469) );
  AND U7742 ( .A(n7470), .B(n7469), .Z(n7608) );
  NANDN U7743 ( .A(n17362), .B(n7471), .Z(n7473) );
  XOR U7744 ( .A(b[7]), .B(a[59]), .Z(n7620) );
  NANDN U7745 ( .A(n17522), .B(n7620), .Z(n7472) );
  AND U7746 ( .A(n7473), .B(n7472), .Z(n7606) );
  NANDN U7747 ( .A(n19116), .B(n7474), .Z(n7476) );
  XOR U7748 ( .A(b[25]), .B(a[41]), .Z(n7623) );
  NANDN U7749 ( .A(n19179), .B(n7623), .Z(n7475) );
  NAND U7750 ( .A(n7476), .B(n7475), .Z(n7605) );
  XNOR U7751 ( .A(n7606), .B(n7605), .Z(n7607) );
  XOR U7752 ( .A(n7608), .B(n7607), .Z(n7576) );
  XNOR U7753 ( .A(n7575), .B(n7576), .Z(n7577) );
  NANDN U7754 ( .A(n18113), .B(n7477), .Z(n7479) );
  XOR U7755 ( .A(b[13]), .B(a[53]), .Z(n7626) );
  NANDN U7756 ( .A(n18229), .B(n7626), .Z(n7478) );
  AND U7757 ( .A(n7479), .B(n7478), .Z(n7570) );
  NANDN U7758 ( .A(n17888), .B(n7480), .Z(n7482) );
  XOR U7759 ( .A(b[11]), .B(a[55]), .Z(n7629) );
  NANDN U7760 ( .A(n18025), .B(n7629), .Z(n7481) );
  NAND U7761 ( .A(n7482), .B(n7481), .Z(n7569) );
  XNOR U7762 ( .A(n7570), .B(n7569), .Z(n7571) );
  NANDN U7763 ( .A(n18487), .B(n7483), .Z(n7485) );
  XOR U7764 ( .A(b[15]), .B(a[51]), .Z(n7632) );
  NANDN U7765 ( .A(n18311), .B(n7632), .Z(n7484) );
  AND U7766 ( .A(n7485), .B(n7484), .Z(n7566) );
  NANDN U7767 ( .A(n18853), .B(n7486), .Z(n7488) );
  XOR U7768 ( .A(b[21]), .B(a[45]), .Z(n7635) );
  NANDN U7769 ( .A(n18926), .B(n7635), .Z(n7487) );
  AND U7770 ( .A(n7488), .B(n7487), .Z(n7564) );
  NANDN U7771 ( .A(n17613), .B(n7489), .Z(n7491) );
  XOR U7772 ( .A(b[9]), .B(a[57]), .Z(n7638) );
  NANDN U7773 ( .A(n17739), .B(n7638), .Z(n7490) );
  NAND U7774 ( .A(n7491), .B(n7490), .Z(n7563) );
  XNOR U7775 ( .A(n7564), .B(n7563), .Z(n7565) );
  XOR U7776 ( .A(n7566), .B(n7565), .Z(n7572) );
  XOR U7777 ( .A(n7571), .B(n7572), .Z(n7578) );
  XOR U7778 ( .A(n7577), .B(n7578), .Z(n7590) );
  XNOR U7779 ( .A(n7589), .B(n7590), .Z(n7521) );
  XNOR U7780 ( .A(n7522), .B(n7521), .Z(n7523) );
  XOR U7781 ( .A(n7524), .B(n7523), .Z(n7642) );
  XNOR U7782 ( .A(n7641), .B(n7642), .Z(n7643) );
  XNOR U7783 ( .A(n7644), .B(n7643), .Z(n7517) );
  XOR U7784 ( .A(n7518), .B(n7517), .Z(n7510) );
  NANDN U7785 ( .A(n7493), .B(n7492), .Z(n7497) );
  NANDN U7786 ( .A(n7495), .B(n7494), .Z(n7496) );
  AND U7787 ( .A(n7497), .B(n7496), .Z(n7509) );
  XOR U7788 ( .A(n7510), .B(n7509), .Z(n7512) );
  XNOR U7789 ( .A(n7511), .B(n7512), .Z(n7503) );
  XNOR U7790 ( .A(n7504), .B(n7503), .Z(n7505) );
  XNOR U7791 ( .A(n7506), .B(n7505), .Z(n7647) );
  XNOR U7792 ( .A(sreg[161]), .B(n7647), .Z(n7649) );
  NANDN U7793 ( .A(sreg[160]), .B(n7498), .Z(n7502) );
  NAND U7794 ( .A(n7500), .B(n7499), .Z(n7501) );
  NAND U7795 ( .A(n7502), .B(n7501), .Z(n7648) );
  XNOR U7796 ( .A(n7649), .B(n7648), .Z(c[161]) );
  NANDN U7797 ( .A(n7504), .B(n7503), .Z(n7508) );
  NANDN U7798 ( .A(n7506), .B(n7505), .Z(n7507) );
  AND U7799 ( .A(n7508), .B(n7507), .Z(n7655) );
  NANDN U7800 ( .A(n7510), .B(n7509), .Z(n7514) );
  NANDN U7801 ( .A(n7512), .B(n7511), .Z(n7513) );
  AND U7802 ( .A(n7514), .B(n7513), .Z(n7653) );
  NANDN U7803 ( .A(n7516), .B(n7515), .Z(n7520) );
  NAND U7804 ( .A(n7518), .B(n7517), .Z(n7519) );
  AND U7805 ( .A(n7520), .B(n7519), .Z(n7660) );
  NANDN U7806 ( .A(n7522), .B(n7521), .Z(n7526) );
  NANDN U7807 ( .A(n7524), .B(n7523), .Z(n7525) );
  AND U7808 ( .A(n7526), .B(n7525), .Z(n7665) );
  NANDN U7809 ( .A(n7528), .B(n7527), .Z(n7532) );
  NAND U7810 ( .A(n7530), .B(n7529), .Z(n7531) );
  AND U7811 ( .A(n7532), .B(n7531), .Z(n7664) );
  XNOR U7812 ( .A(n7665), .B(n7664), .Z(n7667) );
  NANDN U7813 ( .A(n7534), .B(n7533), .Z(n7538) );
  NANDN U7814 ( .A(n7536), .B(n7535), .Z(n7537) );
  AND U7815 ( .A(n7538), .B(n7537), .Z(n7744) );
  NANDN U7816 ( .A(n19237), .B(n7539), .Z(n7541) );
  XOR U7817 ( .A(b[27]), .B(a[40]), .Z(n7688) );
  NANDN U7818 ( .A(n19277), .B(n7688), .Z(n7540) );
  AND U7819 ( .A(n7541), .B(n7540), .Z(n7751) );
  NANDN U7820 ( .A(n17072), .B(n7542), .Z(n7544) );
  XOR U7821 ( .A(b[5]), .B(a[62]), .Z(n7691) );
  NANDN U7822 ( .A(n17223), .B(n7691), .Z(n7543) );
  AND U7823 ( .A(n7544), .B(n7543), .Z(n7749) );
  NANDN U7824 ( .A(n18673), .B(n7545), .Z(n7547) );
  XOR U7825 ( .A(b[19]), .B(a[48]), .Z(n7694) );
  NANDN U7826 ( .A(n18758), .B(n7694), .Z(n7546) );
  NAND U7827 ( .A(n7547), .B(n7546), .Z(n7748) );
  XNOR U7828 ( .A(n7749), .B(n7748), .Z(n7750) );
  XNOR U7829 ( .A(n7751), .B(n7750), .Z(n7742) );
  NANDN U7830 ( .A(n19425), .B(n7548), .Z(n7550) );
  XOR U7831 ( .A(b[31]), .B(a[36]), .Z(n7697) );
  NANDN U7832 ( .A(n19426), .B(n7697), .Z(n7549) );
  AND U7833 ( .A(n7550), .B(n7549), .Z(n7709) );
  NANDN U7834 ( .A(n17067), .B(n7551), .Z(n7553) );
  XOR U7835 ( .A(b[3]), .B(a[64]), .Z(n7700) );
  NANDN U7836 ( .A(n17068), .B(n7700), .Z(n7552) );
  AND U7837 ( .A(n7553), .B(n7552), .Z(n7707) );
  NANDN U7838 ( .A(n18514), .B(n7554), .Z(n7556) );
  XOR U7839 ( .A(b[17]), .B(a[50]), .Z(n7703) );
  NANDN U7840 ( .A(n18585), .B(n7703), .Z(n7555) );
  NAND U7841 ( .A(n7556), .B(n7555), .Z(n7706) );
  XNOR U7842 ( .A(n7707), .B(n7706), .Z(n7708) );
  XOR U7843 ( .A(n7709), .B(n7708), .Z(n7743) );
  XOR U7844 ( .A(n7742), .B(n7743), .Z(n7745) );
  XOR U7845 ( .A(n7744), .B(n7745), .Z(n7677) );
  NANDN U7846 ( .A(n7558), .B(n7557), .Z(n7562) );
  NANDN U7847 ( .A(n7560), .B(n7559), .Z(n7561) );
  AND U7848 ( .A(n7562), .B(n7561), .Z(n7730) );
  NANDN U7849 ( .A(n7564), .B(n7563), .Z(n7568) );
  NANDN U7850 ( .A(n7566), .B(n7565), .Z(n7567) );
  NAND U7851 ( .A(n7568), .B(n7567), .Z(n7731) );
  XNOR U7852 ( .A(n7730), .B(n7731), .Z(n7732) );
  NANDN U7853 ( .A(n7570), .B(n7569), .Z(n7574) );
  NANDN U7854 ( .A(n7572), .B(n7571), .Z(n7573) );
  NAND U7855 ( .A(n7574), .B(n7573), .Z(n7733) );
  XNOR U7856 ( .A(n7732), .B(n7733), .Z(n7676) );
  XNOR U7857 ( .A(n7677), .B(n7676), .Z(n7679) );
  NANDN U7858 ( .A(n7576), .B(n7575), .Z(n7580) );
  NANDN U7859 ( .A(n7578), .B(n7577), .Z(n7579) );
  AND U7860 ( .A(n7580), .B(n7579), .Z(n7678) );
  XOR U7861 ( .A(n7679), .B(n7678), .Z(n7793) );
  NANDN U7862 ( .A(n7582), .B(n7581), .Z(n7586) );
  NANDN U7863 ( .A(n7584), .B(n7583), .Z(n7585) );
  AND U7864 ( .A(n7586), .B(n7585), .Z(n7790) );
  NANDN U7865 ( .A(n7588), .B(n7587), .Z(n7592) );
  NANDN U7866 ( .A(n7590), .B(n7589), .Z(n7591) );
  AND U7867 ( .A(n7592), .B(n7591), .Z(n7673) );
  NANDN U7868 ( .A(n7594), .B(n7593), .Z(n7598) );
  OR U7869 ( .A(n7596), .B(n7595), .Z(n7597) );
  AND U7870 ( .A(n7598), .B(n7597), .Z(n7671) );
  NANDN U7871 ( .A(n7600), .B(n7599), .Z(n7604) );
  NANDN U7872 ( .A(n7602), .B(n7601), .Z(n7603) );
  AND U7873 ( .A(n7604), .B(n7603), .Z(n7737) );
  NANDN U7874 ( .A(n7606), .B(n7605), .Z(n7610) );
  NANDN U7875 ( .A(n7608), .B(n7607), .Z(n7609) );
  NAND U7876 ( .A(n7610), .B(n7609), .Z(n7736) );
  XNOR U7877 ( .A(n7737), .B(n7736), .Z(n7738) );
  NANDN U7878 ( .A(n19394), .B(n7611), .Z(n7613) );
  XOR U7879 ( .A(b[29]), .B(a[38]), .Z(n7763) );
  NANDN U7880 ( .A(n19395), .B(n7763), .Z(n7612) );
  AND U7881 ( .A(n7613), .B(n7612), .Z(n7683) );
  AND U7882 ( .A(b[31]), .B(a[34]), .Z(n7682) );
  XNOR U7883 ( .A(n7683), .B(n7682), .Z(n7684) );
  NAND U7884 ( .A(b[0]), .B(a[66]), .Z(n7614) );
  XNOR U7885 ( .A(b[1]), .B(n7614), .Z(n7616) );
  NANDN U7886 ( .A(b[0]), .B(a[65]), .Z(n7615) );
  NAND U7887 ( .A(n7616), .B(n7615), .Z(n7685) );
  XNOR U7888 ( .A(n7684), .B(n7685), .Z(n7724) );
  NANDN U7889 ( .A(n19005), .B(n7617), .Z(n7619) );
  XOR U7890 ( .A(b[23]), .B(a[44]), .Z(n7766) );
  NANDN U7891 ( .A(n19055), .B(n7766), .Z(n7618) );
  AND U7892 ( .A(n7619), .B(n7618), .Z(n7757) );
  NANDN U7893 ( .A(n17362), .B(n7620), .Z(n7622) );
  XOR U7894 ( .A(b[7]), .B(a[60]), .Z(n7769) );
  NANDN U7895 ( .A(n17522), .B(n7769), .Z(n7621) );
  AND U7896 ( .A(n7622), .B(n7621), .Z(n7755) );
  NANDN U7897 ( .A(n19116), .B(n7623), .Z(n7625) );
  XOR U7898 ( .A(b[25]), .B(a[42]), .Z(n7772) );
  NANDN U7899 ( .A(n19179), .B(n7772), .Z(n7624) );
  NAND U7900 ( .A(n7625), .B(n7624), .Z(n7754) );
  XNOR U7901 ( .A(n7755), .B(n7754), .Z(n7756) );
  XOR U7902 ( .A(n7757), .B(n7756), .Z(n7725) );
  XNOR U7903 ( .A(n7724), .B(n7725), .Z(n7726) );
  NANDN U7904 ( .A(n18113), .B(n7626), .Z(n7628) );
  XOR U7905 ( .A(b[13]), .B(a[54]), .Z(n7775) );
  NANDN U7906 ( .A(n18229), .B(n7775), .Z(n7627) );
  AND U7907 ( .A(n7628), .B(n7627), .Z(n7719) );
  NANDN U7908 ( .A(n17888), .B(n7629), .Z(n7631) );
  XOR U7909 ( .A(b[11]), .B(a[56]), .Z(n7778) );
  NANDN U7910 ( .A(n18025), .B(n7778), .Z(n7630) );
  NAND U7911 ( .A(n7631), .B(n7630), .Z(n7718) );
  XNOR U7912 ( .A(n7719), .B(n7718), .Z(n7720) );
  NANDN U7913 ( .A(n18487), .B(n7632), .Z(n7634) );
  XOR U7914 ( .A(b[15]), .B(a[52]), .Z(n7781) );
  NANDN U7915 ( .A(n18311), .B(n7781), .Z(n7633) );
  AND U7916 ( .A(n7634), .B(n7633), .Z(n7715) );
  NANDN U7917 ( .A(n18853), .B(n7635), .Z(n7637) );
  XOR U7918 ( .A(b[21]), .B(a[46]), .Z(n7784) );
  NANDN U7919 ( .A(n18926), .B(n7784), .Z(n7636) );
  AND U7920 ( .A(n7637), .B(n7636), .Z(n7713) );
  NANDN U7921 ( .A(n17613), .B(n7638), .Z(n7640) );
  XOR U7922 ( .A(b[9]), .B(a[58]), .Z(n7787) );
  NANDN U7923 ( .A(n17739), .B(n7787), .Z(n7639) );
  NAND U7924 ( .A(n7640), .B(n7639), .Z(n7712) );
  XNOR U7925 ( .A(n7713), .B(n7712), .Z(n7714) );
  XOR U7926 ( .A(n7715), .B(n7714), .Z(n7721) );
  XOR U7927 ( .A(n7720), .B(n7721), .Z(n7727) );
  XOR U7928 ( .A(n7726), .B(n7727), .Z(n7739) );
  XNOR U7929 ( .A(n7738), .B(n7739), .Z(n7670) );
  XNOR U7930 ( .A(n7671), .B(n7670), .Z(n7672) );
  XOR U7931 ( .A(n7673), .B(n7672), .Z(n7791) );
  XNOR U7932 ( .A(n7790), .B(n7791), .Z(n7792) );
  XNOR U7933 ( .A(n7793), .B(n7792), .Z(n7666) );
  XOR U7934 ( .A(n7667), .B(n7666), .Z(n7659) );
  NANDN U7935 ( .A(n7642), .B(n7641), .Z(n7646) );
  NANDN U7936 ( .A(n7644), .B(n7643), .Z(n7645) );
  AND U7937 ( .A(n7646), .B(n7645), .Z(n7658) );
  XOR U7938 ( .A(n7659), .B(n7658), .Z(n7661) );
  XNOR U7939 ( .A(n7660), .B(n7661), .Z(n7652) );
  XNOR U7940 ( .A(n7653), .B(n7652), .Z(n7654) );
  XNOR U7941 ( .A(n7655), .B(n7654), .Z(n7796) );
  XNOR U7942 ( .A(sreg[162]), .B(n7796), .Z(n7798) );
  NANDN U7943 ( .A(sreg[161]), .B(n7647), .Z(n7651) );
  NAND U7944 ( .A(n7649), .B(n7648), .Z(n7650) );
  NAND U7945 ( .A(n7651), .B(n7650), .Z(n7797) );
  XNOR U7946 ( .A(n7798), .B(n7797), .Z(c[162]) );
  NANDN U7947 ( .A(n7653), .B(n7652), .Z(n7657) );
  NANDN U7948 ( .A(n7655), .B(n7654), .Z(n7656) );
  AND U7949 ( .A(n7657), .B(n7656), .Z(n7804) );
  NANDN U7950 ( .A(n7659), .B(n7658), .Z(n7663) );
  NANDN U7951 ( .A(n7661), .B(n7660), .Z(n7662) );
  AND U7952 ( .A(n7663), .B(n7662), .Z(n7802) );
  NANDN U7953 ( .A(n7665), .B(n7664), .Z(n7669) );
  NAND U7954 ( .A(n7667), .B(n7666), .Z(n7668) );
  AND U7955 ( .A(n7669), .B(n7668), .Z(n7809) );
  NANDN U7956 ( .A(n7671), .B(n7670), .Z(n7675) );
  NANDN U7957 ( .A(n7673), .B(n7672), .Z(n7674) );
  AND U7958 ( .A(n7675), .B(n7674), .Z(n7938) );
  NANDN U7959 ( .A(n7677), .B(n7676), .Z(n7681) );
  NAND U7960 ( .A(n7679), .B(n7678), .Z(n7680) );
  AND U7961 ( .A(n7681), .B(n7680), .Z(n7937) );
  XNOR U7962 ( .A(n7938), .B(n7937), .Z(n7940) );
  NANDN U7963 ( .A(n7683), .B(n7682), .Z(n7687) );
  NANDN U7964 ( .A(n7685), .B(n7684), .Z(n7686) );
  AND U7965 ( .A(n7687), .B(n7686), .Z(n7885) );
  NANDN U7966 ( .A(n19237), .B(n7688), .Z(n7690) );
  XOR U7967 ( .A(b[27]), .B(a[41]), .Z(n7831) );
  NANDN U7968 ( .A(n19277), .B(n7831), .Z(n7689) );
  AND U7969 ( .A(n7690), .B(n7689), .Z(n7892) );
  NANDN U7970 ( .A(n17072), .B(n7691), .Z(n7693) );
  XOR U7971 ( .A(b[5]), .B(a[63]), .Z(n7834) );
  NANDN U7972 ( .A(n17223), .B(n7834), .Z(n7692) );
  AND U7973 ( .A(n7693), .B(n7692), .Z(n7890) );
  NANDN U7974 ( .A(n18673), .B(n7694), .Z(n7696) );
  XOR U7975 ( .A(b[19]), .B(a[49]), .Z(n7837) );
  NANDN U7976 ( .A(n18758), .B(n7837), .Z(n7695) );
  NAND U7977 ( .A(n7696), .B(n7695), .Z(n7889) );
  XNOR U7978 ( .A(n7890), .B(n7889), .Z(n7891) );
  XNOR U7979 ( .A(n7892), .B(n7891), .Z(n7883) );
  NANDN U7980 ( .A(n19425), .B(n7697), .Z(n7699) );
  XOR U7981 ( .A(b[31]), .B(a[37]), .Z(n7840) );
  NANDN U7982 ( .A(n19426), .B(n7840), .Z(n7698) );
  AND U7983 ( .A(n7699), .B(n7698), .Z(n7852) );
  NANDN U7984 ( .A(n17067), .B(n7700), .Z(n7702) );
  XOR U7985 ( .A(b[3]), .B(a[65]), .Z(n7843) );
  NANDN U7986 ( .A(n17068), .B(n7843), .Z(n7701) );
  AND U7987 ( .A(n7702), .B(n7701), .Z(n7850) );
  NANDN U7988 ( .A(n18514), .B(n7703), .Z(n7705) );
  XOR U7989 ( .A(b[17]), .B(a[51]), .Z(n7846) );
  NANDN U7990 ( .A(n18585), .B(n7846), .Z(n7704) );
  NAND U7991 ( .A(n7705), .B(n7704), .Z(n7849) );
  XNOR U7992 ( .A(n7850), .B(n7849), .Z(n7851) );
  XOR U7993 ( .A(n7852), .B(n7851), .Z(n7884) );
  XOR U7994 ( .A(n7883), .B(n7884), .Z(n7886) );
  XOR U7995 ( .A(n7885), .B(n7886), .Z(n7820) );
  NANDN U7996 ( .A(n7707), .B(n7706), .Z(n7711) );
  NANDN U7997 ( .A(n7709), .B(n7708), .Z(n7710) );
  AND U7998 ( .A(n7711), .B(n7710), .Z(n7873) );
  NANDN U7999 ( .A(n7713), .B(n7712), .Z(n7717) );
  NANDN U8000 ( .A(n7715), .B(n7714), .Z(n7716) );
  NAND U8001 ( .A(n7717), .B(n7716), .Z(n7874) );
  XNOR U8002 ( .A(n7873), .B(n7874), .Z(n7875) );
  NANDN U8003 ( .A(n7719), .B(n7718), .Z(n7723) );
  NANDN U8004 ( .A(n7721), .B(n7720), .Z(n7722) );
  NAND U8005 ( .A(n7723), .B(n7722), .Z(n7876) );
  XNOR U8006 ( .A(n7875), .B(n7876), .Z(n7819) );
  XNOR U8007 ( .A(n7820), .B(n7819), .Z(n7822) );
  NANDN U8008 ( .A(n7725), .B(n7724), .Z(n7729) );
  NANDN U8009 ( .A(n7727), .B(n7726), .Z(n7728) );
  AND U8010 ( .A(n7729), .B(n7728), .Z(n7821) );
  XOR U8011 ( .A(n7822), .B(n7821), .Z(n7934) );
  NANDN U8012 ( .A(n7731), .B(n7730), .Z(n7735) );
  NANDN U8013 ( .A(n7733), .B(n7732), .Z(n7734) );
  AND U8014 ( .A(n7735), .B(n7734), .Z(n7931) );
  NANDN U8015 ( .A(n7737), .B(n7736), .Z(n7741) );
  NANDN U8016 ( .A(n7739), .B(n7738), .Z(n7740) );
  AND U8017 ( .A(n7741), .B(n7740), .Z(n7816) );
  NANDN U8018 ( .A(n7743), .B(n7742), .Z(n7747) );
  OR U8019 ( .A(n7745), .B(n7744), .Z(n7746) );
  AND U8020 ( .A(n7747), .B(n7746), .Z(n7814) );
  NANDN U8021 ( .A(n7749), .B(n7748), .Z(n7753) );
  NANDN U8022 ( .A(n7751), .B(n7750), .Z(n7752) );
  AND U8023 ( .A(n7753), .B(n7752), .Z(n7880) );
  NANDN U8024 ( .A(n7755), .B(n7754), .Z(n7759) );
  NANDN U8025 ( .A(n7757), .B(n7756), .Z(n7758) );
  NAND U8026 ( .A(n7759), .B(n7758), .Z(n7879) );
  XNOR U8027 ( .A(n7880), .B(n7879), .Z(n7882) );
  NAND U8028 ( .A(b[0]), .B(a[67]), .Z(n7760) );
  XNOR U8029 ( .A(b[1]), .B(n7760), .Z(n7762) );
  NANDN U8030 ( .A(b[0]), .B(a[66]), .Z(n7761) );
  NAND U8031 ( .A(n7762), .B(n7761), .Z(n7828) );
  NANDN U8032 ( .A(n19394), .B(n7763), .Z(n7765) );
  XOR U8033 ( .A(b[29]), .B(a[39]), .Z(n7901) );
  NANDN U8034 ( .A(n19395), .B(n7901), .Z(n7764) );
  AND U8035 ( .A(n7765), .B(n7764), .Z(n7826) );
  AND U8036 ( .A(b[31]), .B(a[35]), .Z(n7825) );
  XNOR U8037 ( .A(n7826), .B(n7825), .Z(n7827) );
  XNOR U8038 ( .A(n7828), .B(n7827), .Z(n7868) );
  NANDN U8039 ( .A(n19005), .B(n7766), .Z(n7768) );
  XOR U8040 ( .A(b[23]), .B(a[45]), .Z(n7907) );
  NANDN U8041 ( .A(n19055), .B(n7907), .Z(n7767) );
  AND U8042 ( .A(n7768), .B(n7767), .Z(n7897) );
  NANDN U8043 ( .A(n17362), .B(n7769), .Z(n7771) );
  XOR U8044 ( .A(b[7]), .B(a[61]), .Z(n7910) );
  NANDN U8045 ( .A(n17522), .B(n7910), .Z(n7770) );
  AND U8046 ( .A(n7771), .B(n7770), .Z(n7896) );
  NANDN U8047 ( .A(n19116), .B(n7772), .Z(n7774) );
  XOR U8048 ( .A(b[25]), .B(a[43]), .Z(n7913) );
  NANDN U8049 ( .A(n19179), .B(n7913), .Z(n7773) );
  NAND U8050 ( .A(n7774), .B(n7773), .Z(n7895) );
  XOR U8051 ( .A(n7896), .B(n7895), .Z(n7898) );
  XOR U8052 ( .A(n7897), .B(n7898), .Z(n7867) );
  XOR U8053 ( .A(n7868), .B(n7867), .Z(n7870) );
  NANDN U8054 ( .A(n18113), .B(n7775), .Z(n7777) );
  XOR U8055 ( .A(b[13]), .B(a[55]), .Z(n7916) );
  NANDN U8056 ( .A(n18229), .B(n7916), .Z(n7776) );
  AND U8057 ( .A(n7777), .B(n7776), .Z(n7862) );
  NANDN U8058 ( .A(n17888), .B(n7778), .Z(n7780) );
  XOR U8059 ( .A(b[11]), .B(a[57]), .Z(n7919) );
  NANDN U8060 ( .A(n18025), .B(n7919), .Z(n7779) );
  NAND U8061 ( .A(n7780), .B(n7779), .Z(n7861) );
  XNOR U8062 ( .A(n7862), .B(n7861), .Z(n7864) );
  NANDN U8063 ( .A(n18487), .B(n7781), .Z(n7783) );
  XOR U8064 ( .A(b[15]), .B(a[53]), .Z(n7922) );
  NANDN U8065 ( .A(n18311), .B(n7922), .Z(n7782) );
  AND U8066 ( .A(n7783), .B(n7782), .Z(n7858) );
  NANDN U8067 ( .A(n18853), .B(n7784), .Z(n7786) );
  XOR U8068 ( .A(b[21]), .B(a[47]), .Z(n7925) );
  NANDN U8069 ( .A(n18926), .B(n7925), .Z(n7785) );
  AND U8070 ( .A(n7786), .B(n7785), .Z(n7856) );
  NANDN U8071 ( .A(n17613), .B(n7787), .Z(n7789) );
  XOR U8072 ( .A(b[9]), .B(a[59]), .Z(n7928) );
  NANDN U8073 ( .A(n17739), .B(n7928), .Z(n7788) );
  NAND U8074 ( .A(n7789), .B(n7788), .Z(n7855) );
  XNOR U8075 ( .A(n7856), .B(n7855), .Z(n7857) );
  XNOR U8076 ( .A(n7858), .B(n7857), .Z(n7863) );
  XOR U8077 ( .A(n7864), .B(n7863), .Z(n7869) );
  XOR U8078 ( .A(n7870), .B(n7869), .Z(n7881) );
  XOR U8079 ( .A(n7882), .B(n7881), .Z(n7813) );
  XNOR U8080 ( .A(n7814), .B(n7813), .Z(n7815) );
  XOR U8081 ( .A(n7816), .B(n7815), .Z(n7932) );
  XNOR U8082 ( .A(n7931), .B(n7932), .Z(n7933) );
  XNOR U8083 ( .A(n7934), .B(n7933), .Z(n7939) );
  XOR U8084 ( .A(n7940), .B(n7939), .Z(n7808) );
  NANDN U8085 ( .A(n7791), .B(n7790), .Z(n7795) );
  NANDN U8086 ( .A(n7793), .B(n7792), .Z(n7794) );
  AND U8087 ( .A(n7795), .B(n7794), .Z(n7807) );
  XOR U8088 ( .A(n7808), .B(n7807), .Z(n7810) );
  XNOR U8089 ( .A(n7809), .B(n7810), .Z(n7801) );
  XNOR U8090 ( .A(n7802), .B(n7801), .Z(n7803) );
  XNOR U8091 ( .A(n7804), .B(n7803), .Z(n7943) );
  XNOR U8092 ( .A(sreg[163]), .B(n7943), .Z(n7945) );
  NANDN U8093 ( .A(sreg[162]), .B(n7796), .Z(n7800) );
  NAND U8094 ( .A(n7798), .B(n7797), .Z(n7799) );
  NAND U8095 ( .A(n7800), .B(n7799), .Z(n7944) );
  XNOR U8096 ( .A(n7945), .B(n7944), .Z(c[163]) );
  NANDN U8097 ( .A(n7802), .B(n7801), .Z(n7806) );
  NANDN U8098 ( .A(n7804), .B(n7803), .Z(n7805) );
  AND U8099 ( .A(n7806), .B(n7805), .Z(n7951) );
  NANDN U8100 ( .A(n7808), .B(n7807), .Z(n7812) );
  NANDN U8101 ( .A(n7810), .B(n7809), .Z(n7811) );
  AND U8102 ( .A(n7812), .B(n7811), .Z(n7949) );
  NANDN U8103 ( .A(n7814), .B(n7813), .Z(n7818) );
  NANDN U8104 ( .A(n7816), .B(n7815), .Z(n7817) );
  AND U8105 ( .A(n7818), .B(n7817), .Z(n7961) );
  NANDN U8106 ( .A(n7820), .B(n7819), .Z(n7824) );
  NAND U8107 ( .A(n7822), .B(n7821), .Z(n7823) );
  AND U8108 ( .A(n7824), .B(n7823), .Z(n7960) );
  XNOR U8109 ( .A(n7961), .B(n7960), .Z(n7963) );
  NANDN U8110 ( .A(n7826), .B(n7825), .Z(n7830) );
  NANDN U8111 ( .A(n7828), .B(n7827), .Z(n7829) );
  AND U8112 ( .A(n7830), .B(n7829), .Z(n8028) );
  NANDN U8113 ( .A(n19237), .B(n7831), .Z(n7833) );
  XOR U8114 ( .A(b[27]), .B(a[42]), .Z(n7972) );
  NANDN U8115 ( .A(n19277), .B(n7972), .Z(n7832) );
  AND U8116 ( .A(n7833), .B(n7832), .Z(n8035) );
  NANDN U8117 ( .A(n17072), .B(n7834), .Z(n7836) );
  XOR U8118 ( .A(b[5]), .B(a[64]), .Z(n7975) );
  NANDN U8119 ( .A(n17223), .B(n7975), .Z(n7835) );
  AND U8120 ( .A(n7836), .B(n7835), .Z(n8033) );
  NANDN U8121 ( .A(n18673), .B(n7837), .Z(n7839) );
  XOR U8122 ( .A(b[19]), .B(a[50]), .Z(n7978) );
  NANDN U8123 ( .A(n18758), .B(n7978), .Z(n7838) );
  NAND U8124 ( .A(n7839), .B(n7838), .Z(n8032) );
  XNOR U8125 ( .A(n8033), .B(n8032), .Z(n8034) );
  XNOR U8126 ( .A(n8035), .B(n8034), .Z(n8026) );
  NANDN U8127 ( .A(n19425), .B(n7840), .Z(n7842) );
  XOR U8128 ( .A(b[31]), .B(a[38]), .Z(n7981) );
  NANDN U8129 ( .A(n19426), .B(n7981), .Z(n7841) );
  AND U8130 ( .A(n7842), .B(n7841), .Z(n7993) );
  NANDN U8131 ( .A(n17067), .B(n7843), .Z(n7845) );
  XOR U8132 ( .A(b[3]), .B(a[66]), .Z(n7984) );
  NANDN U8133 ( .A(n17068), .B(n7984), .Z(n7844) );
  AND U8134 ( .A(n7845), .B(n7844), .Z(n7991) );
  NANDN U8135 ( .A(n18514), .B(n7846), .Z(n7848) );
  XOR U8136 ( .A(b[17]), .B(a[52]), .Z(n7987) );
  NANDN U8137 ( .A(n18585), .B(n7987), .Z(n7847) );
  NAND U8138 ( .A(n7848), .B(n7847), .Z(n7990) );
  XNOR U8139 ( .A(n7991), .B(n7990), .Z(n7992) );
  XOR U8140 ( .A(n7993), .B(n7992), .Z(n8027) );
  XOR U8141 ( .A(n8026), .B(n8027), .Z(n8029) );
  XOR U8142 ( .A(n8028), .B(n8029), .Z(n8075) );
  NANDN U8143 ( .A(n7850), .B(n7849), .Z(n7854) );
  NANDN U8144 ( .A(n7852), .B(n7851), .Z(n7853) );
  AND U8145 ( .A(n7854), .B(n7853), .Z(n8014) );
  NANDN U8146 ( .A(n7856), .B(n7855), .Z(n7860) );
  NANDN U8147 ( .A(n7858), .B(n7857), .Z(n7859) );
  NAND U8148 ( .A(n7860), .B(n7859), .Z(n8015) );
  XNOR U8149 ( .A(n8014), .B(n8015), .Z(n8016) );
  NANDN U8150 ( .A(n7862), .B(n7861), .Z(n7866) );
  NAND U8151 ( .A(n7864), .B(n7863), .Z(n7865) );
  NAND U8152 ( .A(n7866), .B(n7865), .Z(n8017) );
  XNOR U8153 ( .A(n8016), .B(n8017), .Z(n8074) );
  XNOR U8154 ( .A(n8075), .B(n8074), .Z(n8077) );
  NAND U8155 ( .A(n7868), .B(n7867), .Z(n7872) );
  NAND U8156 ( .A(n7870), .B(n7869), .Z(n7871) );
  AND U8157 ( .A(n7872), .B(n7871), .Z(n8076) );
  XOR U8158 ( .A(n8077), .B(n8076), .Z(n8089) );
  NANDN U8159 ( .A(n7874), .B(n7873), .Z(n7878) );
  NANDN U8160 ( .A(n7876), .B(n7875), .Z(n7877) );
  AND U8161 ( .A(n7878), .B(n7877), .Z(n8086) );
  NANDN U8162 ( .A(n7884), .B(n7883), .Z(n7888) );
  OR U8163 ( .A(n7886), .B(n7885), .Z(n7887) );
  AND U8164 ( .A(n7888), .B(n7887), .Z(n8081) );
  NANDN U8165 ( .A(n7890), .B(n7889), .Z(n7894) );
  NANDN U8166 ( .A(n7892), .B(n7891), .Z(n7893) );
  AND U8167 ( .A(n7894), .B(n7893), .Z(n8021) );
  NANDN U8168 ( .A(n7896), .B(n7895), .Z(n7900) );
  OR U8169 ( .A(n7898), .B(n7897), .Z(n7899) );
  NAND U8170 ( .A(n7900), .B(n7899), .Z(n8020) );
  XNOR U8171 ( .A(n8021), .B(n8020), .Z(n8022) );
  NANDN U8172 ( .A(n19394), .B(n7901), .Z(n7903) );
  XOR U8173 ( .A(b[29]), .B(a[40]), .Z(n8047) );
  NANDN U8174 ( .A(n19395), .B(n8047), .Z(n7902) );
  AND U8175 ( .A(n7903), .B(n7902), .Z(n7967) );
  AND U8176 ( .A(b[31]), .B(a[36]), .Z(n7966) );
  XNOR U8177 ( .A(n7967), .B(n7966), .Z(n7968) );
  NAND U8178 ( .A(b[0]), .B(a[68]), .Z(n7904) );
  XNOR U8179 ( .A(b[1]), .B(n7904), .Z(n7906) );
  NANDN U8180 ( .A(b[0]), .B(a[67]), .Z(n7905) );
  NAND U8181 ( .A(n7906), .B(n7905), .Z(n7969) );
  XNOR U8182 ( .A(n7968), .B(n7969), .Z(n8008) );
  NANDN U8183 ( .A(n19005), .B(n7907), .Z(n7909) );
  XOR U8184 ( .A(b[23]), .B(a[46]), .Z(n8050) );
  NANDN U8185 ( .A(n19055), .B(n8050), .Z(n7908) );
  AND U8186 ( .A(n7909), .B(n7908), .Z(n8041) );
  NANDN U8187 ( .A(n17362), .B(n7910), .Z(n7912) );
  XOR U8188 ( .A(b[7]), .B(a[62]), .Z(n8053) );
  NANDN U8189 ( .A(n17522), .B(n8053), .Z(n7911) );
  AND U8190 ( .A(n7912), .B(n7911), .Z(n8039) );
  NANDN U8191 ( .A(n19116), .B(n7913), .Z(n7915) );
  XOR U8192 ( .A(b[25]), .B(a[44]), .Z(n8056) );
  NANDN U8193 ( .A(n19179), .B(n8056), .Z(n7914) );
  NAND U8194 ( .A(n7915), .B(n7914), .Z(n8038) );
  XNOR U8195 ( .A(n8039), .B(n8038), .Z(n8040) );
  XOR U8196 ( .A(n8041), .B(n8040), .Z(n8009) );
  XNOR U8197 ( .A(n8008), .B(n8009), .Z(n8010) );
  NANDN U8198 ( .A(n18113), .B(n7916), .Z(n7918) );
  XOR U8199 ( .A(b[13]), .B(a[56]), .Z(n8059) );
  NANDN U8200 ( .A(n18229), .B(n8059), .Z(n7917) );
  AND U8201 ( .A(n7918), .B(n7917), .Z(n8003) );
  NANDN U8202 ( .A(n17888), .B(n7919), .Z(n7921) );
  XOR U8203 ( .A(b[11]), .B(a[58]), .Z(n8062) );
  NANDN U8204 ( .A(n18025), .B(n8062), .Z(n7920) );
  NAND U8205 ( .A(n7921), .B(n7920), .Z(n8002) );
  XNOR U8206 ( .A(n8003), .B(n8002), .Z(n8004) );
  NANDN U8207 ( .A(n18487), .B(n7922), .Z(n7924) );
  XOR U8208 ( .A(b[15]), .B(a[54]), .Z(n8065) );
  NANDN U8209 ( .A(n18311), .B(n8065), .Z(n7923) );
  AND U8210 ( .A(n7924), .B(n7923), .Z(n7999) );
  NANDN U8211 ( .A(n18853), .B(n7925), .Z(n7927) );
  XOR U8212 ( .A(b[21]), .B(a[48]), .Z(n8068) );
  NANDN U8213 ( .A(n18926), .B(n8068), .Z(n7926) );
  AND U8214 ( .A(n7927), .B(n7926), .Z(n7997) );
  NANDN U8215 ( .A(n17613), .B(n7928), .Z(n7930) );
  XOR U8216 ( .A(b[9]), .B(a[60]), .Z(n8071) );
  NANDN U8217 ( .A(n17739), .B(n8071), .Z(n7929) );
  NAND U8218 ( .A(n7930), .B(n7929), .Z(n7996) );
  XNOR U8219 ( .A(n7997), .B(n7996), .Z(n7998) );
  XOR U8220 ( .A(n7999), .B(n7998), .Z(n8005) );
  XOR U8221 ( .A(n8004), .B(n8005), .Z(n8011) );
  XOR U8222 ( .A(n8010), .B(n8011), .Z(n8023) );
  XNOR U8223 ( .A(n8022), .B(n8023), .Z(n8080) );
  XNOR U8224 ( .A(n8081), .B(n8080), .Z(n8082) );
  XOR U8225 ( .A(n8083), .B(n8082), .Z(n8087) );
  XNOR U8226 ( .A(n8086), .B(n8087), .Z(n8088) );
  XNOR U8227 ( .A(n8089), .B(n8088), .Z(n7962) );
  XOR U8228 ( .A(n7963), .B(n7962), .Z(n7955) );
  NANDN U8229 ( .A(n7932), .B(n7931), .Z(n7936) );
  NANDN U8230 ( .A(n7934), .B(n7933), .Z(n7935) );
  AND U8231 ( .A(n7936), .B(n7935), .Z(n7954) );
  XNOR U8232 ( .A(n7955), .B(n7954), .Z(n7956) );
  NANDN U8233 ( .A(n7938), .B(n7937), .Z(n7942) );
  NAND U8234 ( .A(n7940), .B(n7939), .Z(n7941) );
  NAND U8235 ( .A(n7942), .B(n7941), .Z(n7957) );
  XNOR U8236 ( .A(n7956), .B(n7957), .Z(n7948) );
  XNOR U8237 ( .A(n7949), .B(n7948), .Z(n7950) );
  XNOR U8238 ( .A(n7951), .B(n7950), .Z(n8092) );
  XNOR U8239 ( .A(sreg[164]), .B(n8092), .Z(n8094) );
  NANDN U8240 ( .A(sreg[163]), .B(n7943), .Z(n7947) );
  NAND U8241 ( .A(n7945), .B(n7944), .Z(n7946) );
  NAND U8242 ( .A(n7947), .B(n7946), .Z(n8093) );
  XNOR U8243 ( .A(n8094), .B(n8093), .Z(c[164]) );
  NANDN U8244 ( .A(n7949), .B(n7948), .Z(n7953) );
  NANDN U8245 ( .A(n7951), .B(n7950), .Z(n7952) );
  AND U8246 ( .A(n7953), .B(n7952), .Z(n8100) );
  NANDN U8247 ( .A(n7955), .B(n7954), .Z(n7959) );
  NANDN U8248 ( .A(n7957), .B(n7956), .Z(n7958) );
  AND U8249 ( .A(n7959), .B(n7958), .Z(n8098) );
  NANDN U8250 ( .A(n7961), .B(n7960), .Z(n7965) );
  NAND U8251 ( .A(n7963), .B(n7962), .Z(n7964) );
  AND U8252 ( .A(n7965), .B(n7964), .Z(n8105) );
  NANDN U8253 ( .A(n7967), .B(n7966), .Z(n7971) );
  NANDN U8254 ( .A(n7969), .B(n7968), .Z(n7970) );
  AND U8255 ( .A(n7971), .B(n7970), .Z(n8189) );
  NANDN U8256 ( .A(n19237), .B(n7972), .Z(n7974) );
  XOR U8257 ( .A(b[27]), .B(a[43]), .Z(n8133) );
  NANDN U8258 ( .A(n19277), .B(n8133), .Z(n7973) );
  AND U8259 ( .A(n7974), .B(n7973), .Z(n8196) );
  NANDN U8260 ( .A(n17072), .B(n7975), .Z(n7977) );
  XOR U8261 ( .A(b[5]), .B(a[65]), .Z(n8136) );
  NANDN U8262 ( .A(n17223), .B(n8136), .Z(n7976) );
  AND U8263 ( .A(n7977), .B(n7976), .Z(n8194) );
  NANDN U8264 ( .A(n18673), .B(n7978), .Z(n7980) );
  XOR U8265 ( .A(b[19]), .B(a[51]), .Z(n8139) );
  NANDN U8266 ( .A(n18758), .B(n8139), .Z(n7979) );
  NAND U8267 ( .A(n7980), .B(n7979), .Z(n8193) );
  XNOR U8268 ( .A(n8194), .B(n8193), .Z(n8195) );
  XNOR U8269 ( .A(n8196), .B(n8195), .Z(n8187) );
  NANDN U8270 ( .A(n19425), .B(n7981), .Z(n7983) );
  XOR U8271 ( .A(b[31]), .B(a[39]), .Z(n8142) );
  NANDN U8272 ( .A(n19426), .B(n8142), .Z(n7982) );
  AND U8273 ( .A(n7983), .B(n7982), .Z(n8154) );
  NANDN U8274 ( .A(n17067), .B(n7984), .Z(n7986) );
  XOR U8275 ( .A(b[3]), .B(a[67]), .Z(n8145) );
  NANDN U8276 ( .A(n17068), .B(n8145), .Z(n7985) );
  AND U8277 ( .A(n7986), .B(n7985), .Z(n8152) );
  NANDN U8278 ( .A(n18514), .B(n7987), .Z(n7989) );
  XOR U8279 ( .A(b[17]), .B(a[53]), .Z(n8148) );
  NANDN U8280 ( .A(n18585), .B(n8148), .Z(n7988) );
  NAND U8281 ( .A(n7989), .B(n7988), .Z(n8151) );
  XNOR U8282 ( .A(n8152), .B(n8151), .Z(n8153) );
  XOR U8283 ( .A(n8154), .B(n8153), .Z(n8188) );
  XOR U8284 ( .A(n8187), .B(n8188), .Z(n8190) );
  XOR U8285 ( .A(n8189), .B(n8190), .Z(n8122) );
  NANDN U8286 ( .A(n7991), .B(n7990), .Z(n7995) );
  NANDN U8287 ( .A(n7993), .B(n7992), .Z(n7994) );
  AND U8288 ( .A(n7995), .B(n7994), .Z(n8175) );
  NANDN U8289 ( .A(n7997), .B(n7996), .Z(n8001) );
  NANDN U8290 ( .A(n7999), .B(n7998), .Z(n8000) );
  NAND U8291 ( .A(n8001), .B(n8000), .Z(n8176) );
  XNOR U8292 ( .A(n8175), .B(n8176), .Z(n8177) );
  NANDN U8293 ( .A(n8003), .B(n8002), .Z(n8007) );
  NANDN U8294 ( .A(n8005), .B(n8004), .Z(n8006) );
  NAND U8295 ( .A(n8007), .B(n8006), .Z(n8178) );
  XNOR U8296 ( .A(n8177), .B(n8178), .Z(n8121) );
  XNOR U8297 ( .A(n8122), .B(n8121), .Z(n8124) );
  NANDN U8298 ( .A(n8009), .B(n8008), .Z(n8013) );
  NANDN U8299 ( .A(n8011), .B(n8010), .Z(n8012) );
  AND U8300 ( .A(n8013), .B(n8012), .Z(n8123) );
  XOR U8301 ( .A(n8124), .B(n8123), .Z(n8237) );
  NANDN U8302 ( .A(n8015), .B(n8014), .Z(n8019) );
  NANDN U8303 ( .A(n8017), .B(n8016), .Z(n8018) );
  AND U8304 ( .A(n8019), .B(n8018), .Z(n8235) );
  NANDN U8305 ( .A(n8021), .B(n8020), .Z(n8025) );
  NANDN U8306 ( .A(n8023), .B(n8022), .Z(n8024) );
  AND U8307 ( .A(n8025), .B(n8024), .Z(n8118) );
  NANDN U8308 ( .A(n8027), .B(n8026), .Z(n8031) );
  OR U8309 ( .A(n8029), .B(n8028), .Z(n8030) );
  AND U8310 ( .A(n8031), .B(n8030), .Z(n8116) );
  NANDN U8311 ( .A(n8033), .B(n8032), .Z(n8037) );
  NANDN U8312 ( .A(n8035), .B(n8034), .Z(n8036) );
  AND U8313 ( .A(n8037), .B(n8036), .Z(n8182) );
  NANDN U8314 ( .A(n8039), .B(n8038), .Z(n8043) );
  NANDN U8315 ( .A(n8041), .B(n8040), .Z(n8042) );
  NAND U8316 ( .A(n8043), .B(n8042), .Z(n8181) );
  XNOR U8317 ( .A(n8182), .B(n8181), .Z(n8183) );
  NAND U8318 ( .A(b[0]), .B(a[69]), .Z(n8044) );
  XNOR U8319 ( .A(b[1]), .B(n8044), .Z(n8046) );
  NANDN U8320 ( .A(b[0]), .B(a[68]), .Z(n8045) );
  NAND U8321 ( .A(n8046), .B(n8045), .Z(n8130) );
  NANDN U8322 ( .A(n19394), .B(n8047), .Z(n8049) );
  XOR U8323 ( .A(b[29]), .B(a[41]), .Z(n8208) );
  NANDN U8324 ( .A(n19395), .B(n8208), .Z(n8048) );
  AND U8325 ( .A(n8049), .B(n8048), .Z(n8128) );
  AND U8326 ( .A(b[31]), .B(a[37]), .Z(n8127) );
  XNOR U8327 ( .A(n8128), .B(n8127), .Z(n8129) );
  XNOR U8328 ( .A(n8130), .B(n8129), .Z(n8169) );
  NANDN U8329 ( .A(n19005), .B(n8050), .Z(n8052) );
  XOR U8330 ( .A(b[23]), .B(a[47]), .Z(n8211) );
  NANDN U8331 ( .A(n19055), .B(n8211), .Z(n8051) );
  AND U8332 ( .A(n8052), .B(n8051), .Z(n8202) );
  NANDN U8333 ( .A(n17362), .B(n8053), .Z(n8055) );
  XOR U8334 ( .A(b[7]), .B(a[63]), .Z(n8214) );
  NANDN U8335 ( .A(n17522), .B(n8214), .Z(n8054) );
  AND U8336 ( .A(n8055), .B(n8054), .Z(n8200) );
  NANDN U8337 ( .A(n19116), .B(n8056), .Z(n8058) );
  XOR U8338 ( .A(b[25]), .B(a[45]), .Z(n8217) );
  NANDN U8339 ( .A(n19179), .B(n8217), .Z(n8057) );
  NAND U8340 ( .A(n8058), .B(n8057), .Z(n8199) );
  XNOR U8341 ( .A(n8200), .B(n8199), .Z(n8201) );
  XOR U8342 ( .A(n8202), .B(n8201), .Z(n8170) );
  XNOR U8343 ( .A(n8169), .B(n8170), .Z(n8171) );
  NANDN U8344 ( .A(n18113), .B(n8059), .Z(n8061) );
  XOR U8345 ( .A(b[13]), .B(a[57]), .Z(n8220) );
  NANDN U8346 ( .A(n18229), .B(n8220), .Z(n8060) );
  AND U8347 ( .A(n8061), .B(n8060), .Z(n8164) );
  NANDN U8348 ( .A(n17888), .B(n8062), .Z(n8064) );
  XOR U8349 ( .A(b[11]), .B(a[59]), .Z(n8223) );
  NANDN U8350 ( .A(n18025), .B(n8223), .Z(n8063) );
  NAND U8351 ( .A(n8064), .B(n8063), .Z(n8163) );
  XNOR U8352 ( .A(n8164), .B(n8163), .Z(n8165) );
  NANDN U8353 ( .A(n18487), .B(n8065), .Z(n8067) );
  XOR U8354 ( .A(b[15]), .B(a[55]), .Z(n8226) );
  NANDN U8355 ( .A(n18311), .B(n8226), .Z(n8066) );
  AND U8356 ( .A(n8067), .B(n8066), .Z(n8160) );
  NANDN U8357 ( .A(n18853), .B(n8068), .Z(n8070) );
  XOR U8358 ( .A(b[21]), .B(a[49]), .Z(n8229) );
  NANDN U8359 ( .A(n18926), .B(n8229), .Z(n8069) );
  AND U8360 ( .A(n8070), .B(n8069), .Z(n8158) );
  NANDN U8361 ( .A(n17613), .B(n8071), .Z(n8073) );
  XOR U8362 ( .A(b[9]), .B(a[61]), .Z(n8232) );
  NANDN U8363 ( .A(n17739), .B(n8232), .Z(n8072) );
  NAND U8364 ( .A(n8073), .B(n8072), .Z(n8157) );
  XNOR U8365 ( .A(n8158), .B(n8157), .Z(n8159) );
  XOR U8366 ( .A(n8160), .B(n8159), .Z(n8166) );
  XOR U8367 ( .A(n8165), .B(n8166), .Z(n8172) );
  XOR U8368 ( .A(n8171), .B(n8172), .Z(n8184) );
  XNOR U8369 ( .A(n8183), .B(n8184), .Z(n8115) );
  XNOR U8370 ( .A(n8116), .B(n8115), .Z(n8117) );
  XOR U8371 ( .A(n8118), .B(n8117), .Z(n8236) );
  XOR U8372 ( .A(n8235), .B(n8236), .Z(n8238) );
  XOR U8373 ( .A(n8237), .B(n8238), .Z(n8112) );
  NANDN U8374 ( .A(n8075), .B(n8074), .Z(n8079) );
  NAND U8375 ( .A(n8077), .B(n8076), .Z(n8078) );
  AND U8376 ( .A(n8079), .B(n8078), .Z(n8110) );
  NANDN U8377 ( .A(n8081), .B(n8080), .Z(n8085) );
  NANDN U8378 ( .A(n8083), .B(n8082), .Z(n8084) );
  AND U8379 ( .A(n8085), .B(n8084), .Z(n8109) );
  XNOR U8380 ( .A(n8110), .B(n8109), .Z(n8111) );
  XNOR U8381 ( .A(n8112), .B(n8111), .Z(n8103) );
  NANDN U8382 ( .A(n8087), .B(n8086), .Z(n8091) );
  NANDN U8383 ( .A(n8089), .B(n8088), .Z(n8090) );
  NAND U8384 ( .A(n8091), .B(n8090), .Z(n8104) );
  XOR U8385 ( .A(n8103), .B(n8104), .Z(n8106) );
  XNOR U8386 ( .A(n8105), .B(n8106), .Z(n8097) );
  XNOR U8387 ( .A(n8098), .B(n8097), .Z(n8099) );
  XNOR U8388 ( .A(n8100), .B(n8099), .Z(n8241) );
  XNOR U8389 ( .A(sreg[165]), .B(n8241), .Z(n8243) );
  NANDN U8390 ( .A(sreg[164]), .B(n8092), .Z(n8096) );
  NAND U8391 ( .A(n8094), .B(n8093), .Z(n8095) );
  NAND U8392 ( .A(n8096), .B(n8095), .Z(n8242) );
  XNOR U8393 ( .A(n8243), .B(n8242), .Z(c[165]) );
  NANDN U8394 ( .A(n8098), .B(n8097), .Z(n8102) );
  NANDN U8395 ( .A(n8100), .B(n8099), .Z(n8101) );
  AND U8396 ( .A(n8102), .B(n8101), .Z(n8249) );
  NANDN U8397 ( .A(n8104), .B(n8103), .Z(n8108) );
  NANDN U8398 ( .A(n8106), .B(n8105), .Z(n8107) );
  AND U8399 ( .A(n8108), .B(n8107), .Z(n8247) );
  NANDN U8400 ( .A(n8110), .B(n8109), .Z(n8114) );
  NANDN U8401 ( .A(n8112), .B(n8111), .Z(n8113) );
  AND U8402 ( .A(n8114), .B(n8113), .Z(n8255) );
  NANDN U8403 ( .A(n8116), .B(n8115), .Z(n8120) );
  NANDN U8404 ( .A(n8118), .B(n8117), .Z(n8119) );
  AND U8405 ( .A(n8120), .B(n8119), .Z(n8259) );
  NANDN U8406 ( .A(n8122), .B(n8121), .Z(n8126) );
  NAND U8407 ( .A(n8124), .B(n8123), .Z(n8125) );
  AND U8408 ( .A(n8126), .B(n8125), .Z(n8258) );
  XNOR U8409 ( .A(n8259), .B(n8258), .Z(n8261) );
  NANDN U8410 ( .A(n8128), .B(n8127), .Z(n8132) );
  NANDN U8411 ( .A(n8130), .B(n8129), .Z(n8131) );
  AND U8412 ( .A(n8132), .B(n8131), .Z(n8338) );
  NANDN U8413 ( .A(n19237), .B(n8133), .Z(n8135) );
  XOR U8414 ( .A(b[27]), .B(a[44]), .Z(n8282) );
  NANDN U8415 ( .A(n19277), .B(n8282), .Z(n8134) );
  AND U8416 ( .A(n8135), .B(n8134), .Z(n8345) );
  NANDN U8417 ( .A(n17072), .B(n8136), .Z(n8138) );
  XOR U8418 ( .A(b[5]), .B(a[66]), .Z(n8285) );
  NANDN U8419 ( .A(n17223), .B(n8285), .Z(n8137) );
  AND U8420 ( .A(n8138), .B(n8137), .Z(n8343) );
  NANDN U8421 ( .A(n18673), .B(n8139), .Z(n8141) );
  XOR U8422 ( .A(b[19]), .B(a[52]), .Z(n8288) );
  NANDN U8423 ( .A(n18758), .B(n8288), .Z(n8140) );
  NAND U8424 ( .A(n8141), .B(n8140), .Z(n8342) );
  XNOR U8425 ( .A(n8343), .B(n8342), .Z(n8344) );
  XNOR U8426 ( .A(n8345), .B(n8344), .Z(n8336) );
  NANDN U8427 ( .A(n19425), .B(n8142), .Z(n8144) );
  XOR U8428 ( .A(b[31]), .B(a[40]), .Z(n8291) );
  NANDN U8429 ( .A(n19426), .B(n8291), .Z(n8143) );
  AND U8430 ( .A(n8144), .B(n8143), .Z(n8303) );
  NANDN U8431 ( .A(n17067), .B(n8145), .Z(n8147) );
  XOR U8432 ( .A(b[3]), .B(a[68]), .Z(n8294) );
  NANDN U8433 ( .A(n17068), .B(n8294), .Z(n8146) );
  AND U8434 ( .A(n8147), .B(n8146), .Z(n8301) );
  NANDN U8435 ( .A(n18514), .B(n8148), .Z(n8150) );
  XOR U8436 ( .A(b[17]), .B(a[54]), .Z(n8297) );
  NANDN U8437 ( .A(n18585), .B(n8297), .Z(n8149) );
  NAND U8438 ( .A(n8150), .B(n8149), .Z(n8300) );
  XNOR U8439 ( .A(n8301), .B(n8300), .Z(n8302) );
  XOR U8440 ( .A(n8303), .B(n8302), .Z(n8337) );
  XOR U8441 ( .A(n8336), .B(n8337), .Z(n8339) );
  XOR U8442 ( .A(n8338), .B(n8339), .Z(n8271) );
  NANDN U8443 ( .A(n8152), .B(n8151), .Z(n8156) );
  NANDN U8444 ( .A(n8154), .B(n8153), .Z(n8155) );
  AND U8445 ( .A(n8156), .B(n8155), .Z(n8324) );
  NANDN U8446 ( .A(n8158), .B(n8157), .Z(n8162) );
  NANDN U8447 ( .A(n8160), .B(n8159), .Z(n8161) );
  NAND U8448 ( .A(n8162), .B(n8161), .Z(n8325) );
  XNOR U8449 ( .A(n8324), .B(n8325), .Z(n8326) );
  NANDN U8450 ( .A(n8164), .B(n8163), .Z(n8168) );
  NANDN U8451 ( .A(n8166), .B(n8165), .Z(n8167) );
  NAND U8452 ( .A(n8168), .B(n8167), .Z(n8327) );
  XNOR U8453 ( .A(n8326), .B(n8327), .Z(n8270) );
  XNOR U8454 ( .A(n8271), .B(n8270), .Z(n8273) );
  NANDN U8455 ( .A(n8170), .B(n8169), .Z(n8174) );
  NANDN U8456 ( .A(n8172), .B(n8171), .Z(n8173) );
  AND U8457 ( .A(n8174), .B(n8173), .Z(n8272) );
  XOR U8458 ( .A(n8273), .B(n8272), .Z(n8387) );
  NANDN U8459 ( .A(n8176), .B(n8175), .Z(n8180) );
  NANDN U8460 ( .A(n8178), .B(n8177), .Z(n8179) );
  AND U8461 ( .A(n8180), .B(n8179), .Z(n8384) );
  NANDN U8462 ( .A(n8182), .B(n8181), .Z(n8186) );
  NANDN U8463 ( .A(n8184), .B(n8183), .Z(n8185) );
  AND U8464 ( .A(n8186), .B(n8185), .Z(n8267) );
  NANDN U8465 ( .A(n8188), .B(n8187), .Z(n8192) );
  OR U8466 ( .A(n8190), .B(n8189), .Z(n8191) );
  AND U8467 ( .A(n8192), .B(n8191), .Z(n8265) );
  NANDN U8468 ( .A(n8194), .B(n8193), .Z(n8198) );
  NANDN U8469 ( .A(n8196), .B(n8195), .Z(n8197) );
  AND U8470 ( .A(n8198), .B(n8197), .Z(n8331) );
  NANDN U8471 ( .A(n8200), .B(n8199), .Z(n8204) );
  NANDN U8472 ( .A(n8202), .B(n8201), .Z(n8203) );
  NAND U8473 ( .A(n8204), .B(n8203), .Z(n8330) );
  XNOR U8474 ( .A(n8331), .B(n8330), .Z(n8332) );
  NAND U8475 ( .A(b[0]), .B(a[70]), .Z(n8205) );
  XNOR U8476 ( .A(b[1]), .B(n8205), .Z(n8207) );
  NANDN U8477 ( .A(b[0]), .B(a[69]), .Z(n8206) );
  NAND U8478 ( .A(n8207), .B(n8206), .Z(n8279) );
  NANDN U8479 ( .A(n19394), .B(n8208), .Z(n8210) );
  XOR U8480 ( .A(b[29]), .B(a[42]), .Z(n8357) );
  NANDN U8481 ( .A(n19395), .B(n8357), .Z(n8209) );
  AND U8482 ( .A(n8210), .B(n8209), .Z(n8277) );
  AND U8483 ( .A(b[31]), .B(a[38]), .Z(n8276) );
  XNOR U8484 ( .A(n8277), .B(n8276), .Z(n8278) );
  XNOR U8485 ( .A(n8279), .B(n8278), .Z(n8318) );
  NANDN U8486 ( .A(n19005), .B(n8211), .Z(n8213) );
  XOR U8487 ( .A(b[23]), .B(a[48]), .Z(n8360) );
  NANDN U8488 ( .A(n19055), .B(n8360), .Z(n8212) );
  AND U8489 ( .A(n8213), .B(n8212), .Z(n8351) );
  NANDN U8490 ( .A(n17362), .B(n8214), .Z(n8216) );
  XOR U8491 ( .A(b[7]), .B(a[64]), .Z(n8363) );
  NANDN U8492 ( .A(n17522), .B(n8363), .Z(n8215) );
  AND U8493 ( .A(n8216), .B(n8215), .Z(n8349) );
  NANDN U8494 ( .A(n19116), .B(n8217), .Z(n8219) );
  XOR U8495 ( .A(b[25]), .B(a[46]), .Z(n8366) );
  NANDN U8496 ( .A(n19179), .B(n8366), .Z(n8218) );
  NAND U8497 ( .A(n8219), .B(n8218), .Z(n8348) );
  XNOR U8498 ( .A(n8349), .B(n8348), .Z(n8350) );
  XOR U8499 ( .A(n8351), .B(n8350), .Z(n8319) );
  XNOR U8500 ( .A(n8318), .B(n8319), .Z(n8320) );
  NANDN U8501 ( .A(n18113), .B(n8220), .Z(n8222) );
  XOR U8502 ( .A(b[13]), .B(a[58]), .Z(n8369) );
  NANDN U8503 ( .A(n18229), .B(n8369), .Z(n8221) );
  AND U8504 ( .A(n8222), .B(n8221), .Z(n8313) );
  NANDN U8505 ( .A(n17888), .B(n8223), .Z(n8225) );
  XOR U8506 ( .A(b[11]), .B(a[60]), .Z(n8372) );
  NANDN U8507 ( .A(n18025), .B(n8372), .Z(n8224) );
  NAND U8508 ( .A(n8225), .B(n8224), .Z(n8312) );
  XNOR U8509 ( .A(n8313), .B(n8312), .Z(n8314) );
  NANDN U8510 ( .A(n18487), .B(n8226), .Z(n8228) );
  XOR U8511 ( .A(b[15]), .B(a[56]), .Z(n8375) );
  NANDN U8512 ( .A(n18311), .B(n8375), .Z(n8227) );
  AND U8513 ( .A(n8228), .B(n8227), .Z(n8309) );
  NANDN U8514 ( .A(n18853), .B(n8229), .Z(n8231) );
  XOR U8515 ( .A(b[21]), .B(a[50]), .Z(n8378) );
  NANDN U8516 ( .A(n18926), .B(n8378), .Z(n8230) );
  AND U8517 ( .A(n8231), .B(n8230), .Z(n8307) );
  NANDN U8518 ( .A(n17613), .B(n8232), .Z(n8234) );
  XOR U8519 ( .A(b[9]), .B(a[62]), .Z(n8381) );
  NANDN U8520 ( .A(n17739), .B(n8381), .Z(n8233) );
  NAND U8521 ( .A(n8234), .B(n8233), .Z(n8306) );
  XNOR U8522 ( .A(n8307), .B(n8306), .Z(n8308) );
  XOR U8523 ( .A(n8309), .B(n8308), .Z(n8315) );
  XOR U8524 ( .A(n8314), .B(n8315), .Z(n8321) );
  XOR U8525 ( .A(n8320), .B(n8321), .Z(n8333) );
  XNOR U8526 ( .A(n8332), .B(n8333), .Z(n8264) );
  XNOR U8527 ( .A(n8265), .B(n8264), .Z(n8266) );
  XOR U8528 ( .A(n8267), .B(n8266), .Z(n8385) );
  XNOR U8529 ( .A(n8384), .B(n8385), .Z(n8386) );
  XNOR U8530 ( .A(n8387), .B(n8386), .Z(n8260) );
  XOR U8531 ( .A(n8261), .B(n8260), .Z(n8253) );
  NANDN U8532 ( .A(n8236), .B(n8235), .Z(n8240) );
  OR U8533 ( .A(n8238), .B(n8237), .Z(n8239) );
  AND U8534 ( .A(n8240), .B(n8239), .Z(n8252) );
  XNOR U8535 ( .A(n8253), .B(n8252), .Z(n8254) );
  XNOR U8536 ( .A(n8255), .B(n8254), .Z(n8246) );
  XNOR U8537 ( .A(n8247), .B(n8246), .Z(n8248) );
  XNOR U8538 ( .A(n8249), .B(n8248), .Z(n8390) );
  XNOR U8539 ( .A(sreg[166]), .B(n8390), .Z(n8392) );
  NANDN U8540 ( .A(sreg[165]), .B(n8241), .Z(n8245) );
  NAND U8541 ( .A(n8243), .B(n8242), .Z(n8244) );
  NAND U8542 ( .A(n8245), .B(n8244), .Z(n8391) );
  XNOR U8543 ( .A(n8392), .B(n8391), .Z(c[166]) );
  NANDN U8544 ( .A(n8247), .B(n8246), .Z(n8251) );
  NANDN U8545 ( .A(n8249), .B(n8248), .Z(n8250) );
  AND U8546 ( .A(n8251), .B(n8250), .Z(n8398) );
  NANDN U8547 ( .A(n8253), .B(n8252), .Z(n8257) );
  NANDN U8548 ( .A(n8255), .B(n8254), .Z(n8256) );
  AND U8549 ( .A(n8257), .B(n8256), .Z(n8396) );
  NANDN U8550 ( .A(n8259), .B(n8258), .Z(n8263) );
  NAND U8551 ( .A(n8261), .B(n8260), .Z(n8262) );
  AND U8552 ( .A(n8263), .B(n8262), .Z(n8403) );
  NANDN U8553 ( .A(n8265), .B(n8264), .Z(n8269) );
  NANDN U8554 ( .A(n8267), .B(n8266), .Z(n8268) );
  AND U8555 ( .A(n8269), .B(n8268), .Z(n8408) );
  NANDN U8556 ( .A(n8271), .B(n8270), .Z(n8275) );
  NAND U8557 ( .A(n8273), .B(n8272), .Z(n8274) );
  AND U8558 ( .A(n8275), .B(n8274), .Z(n8407) );
  XNOR U8559 ( .A(n8408), .B(n8407), .Z(n8410) );
  NANDN U8560 ( .A(n8277), .B(n8276), .Z(n8281) );
  NANDN U8561 ( .A(n8279), .B(n8278), .Z(n8280) );
  AND U8562 ( .A(n8281), .B(n8280), .Z(n8487) );
  NANDN U8563 ( .A(n19237), .B(n8282), .Z(n8284) );
  XOR U8564 ( .A(b[27]), .B(a[45]), .Z(n8431) );
  NANDN U8565 ( .A(n19277), .B(n8431), .Z(n8283) );
  AND U8566 ( .A(n8284), .B(n8283), .Z(n8494) );
  NANDN U8567 ( .A(n17072), .B(n8285), .Z(n8287) );
  XOR U8568 ( .A(b[5]), .B(a[67]), .Z(n8434) );
  NANDN U8569 ( .A(n17223), .B(n8434), .Z(n8286) );
  AND U8570 ( .A(n8287), .B(n8286), .Z(n8492) );
  NANDN U8571 ( .A(n18673), .B(n8288), .Z(n8290) );
  XOR U8572 ( .A(b[19]), .B(a[53]), .Z(n8437) );
  NANDN U8573 ( .A(n18758), .B(n8437), .Z(n8289) );
  NAND U8574 ( .A(n8290), .B(n8289), .Z(n8491) );
  XNOR U8575 ( .A(n8492), .B(n8491), .Z(n8493) );
  XNOR U8576 ( .A(n8494), .B(n8493), .Z(n8485) );
  NANDN U8577 ( .A(n19425), .B(n8291), .Z(n8293) );
  XOR U8578 ( .A(b[31]), .B(a[41]), .Z(n8440) );
  NANDN U8579 ( .A(n19426), .B(n8440), .Z(n8292) );
  AND U8580 ( .A(n8293), .B(n8292), .Z(n8452) );
  NANDN U8581 ( .A(n17067), .B(n8294), .Z(n8296) );
  XOR U8582 ( .A(b[3]), .B(a[69]), .Z(n8443) );
  NANDN U8583 ( .A(n17068), .B(n8443), .Z(n8295) );
  AND U8584 ( .A(n8296), .B(n8295), .Z(n8450) );
  NANDN U8585 ( .A(n18514), .B(n8297), .Z(n8299) );
  XOR U8586 ( .A(b[17]), .B(a[55]), .Z(n8446) );
  NANDN U8587 ( .A(n18585), .B(n8446), .Z(n8298) );
  NAND U8588 ( .A(n8299), .B(n8298), .Z(n8449) );
  XNOR U8589 ( .A(n8450), .B(n8449), .Z(n8451) );
  XOR U8590 ( .A(n8452), .B(n8451), .Z(n8486) );
  XOR U8591 ( .A(n8485), .B(n8486), .Z(n8488) );
  XOR U8592 ( .A(n8487), .B(n8488), .Z(n8420) );
  NANDN U8593 ( .A(n8301), .B(n8300), .Z(n8305) );
  NANDN U8594 ( .A(n8303), .B(n8302), .Z(n8304) );
  AND U8595 ( .A(n8305), .B(n8304), .Z(n8473) );
  NANDN U8596 ( .A(n8307), .B(n8306), .Z(n8311) );
  NANDN U8597 ( .A(n8309), .B(n8308), .Z(n8310) );
  NAND U8598 ( .A(n8311), .B(n8310), .Z(n8474) );
  XNOR U8599 ( .A(n8473), .B(n8474), .Z(n8475) );
  NANDN U8600 ( .A(n8313), .B(n8312), .Z(n8317) );
  NANDN U8601 ( .A(n8315), .B(n8314), .Z(n8316) );
  NAND U8602 ( .A(n8317), .B(n8316), .Z(n8476) );
  XNOR U8603 ( .A(n8475), .B(n8476), .Z(n8419) );
  XNOR U8604 ( .A(n8420), .B(n8419), .Z(n8422) );
  NANDN U8605 ( .A(n8319), .B(n8318), .Z(n8323) );
  NANDN U8606 ( .A(n8321), .B(n8320), .Z(n8322) );
  AND U8607 ( .A(n8323), .B(n8322), .Z(n8421) );
  XOR U8608 ( .A(n8422), .B(n8421), .Z(n8536) );
  NANDN U8609 ( .A(n8325), .B(n8324), .Z(n8329) );
  NANDN U8610 ( .A(n8327), .B(n8326), .Z(n8328) );
  AND U8611 ( .A(n8329), .B(n8328), .Z(n8533) );
  NANDN U8612 ( .A(n8331), .B(n8330), .Z(n8335) );
  NANDN U8613 ( .A(n8333), .B(n8332), .Z(n8334) );
  AND U8614 ( .A(n8335), .B(n8334), .Z(n8416) );
  NANDN U8615 ( .A(n8337), .B(n8336), .Z(n8341) );
  OR U8616 ( .A(n8339), .B(n8338), .Z(n8340) );
  AND U8617 ( .A(n8341), .B(n8340), .Z(n8414) );
  NANDN U8618 ( .A(n8343), .B(n8342), .Z(n8347) );
  NANDN U8619 ( .A(n8345), .B(n8344), .Z(n8346) );
  AND U8620 ( .A(n8347), .B(n8346), .Z(n8480) );
  NANDN U8621 ( .A(n8349), .B(n8348), .Z(n8353) );
  NANDN U8622 ( .A(n8351), .B(n8350), .Z(n8352) );
  NAND U8623 ( .A(n8353), .B(n8352), .Z(n8479) );
  XNOR U8624 ( .A(n8480), .B(n8479), .Z(n8481) );
  NAND U8625 ( .A(b[0]), .B(a[71]), .Z(n8354) );
  XNOR U8626 ( .A(b[1]), .B(n8354), .Z(n8356) );
  NANDN U8627 ( .A(b[0]), .B(a[70]), .Z(n8355) );
  NAND U8628 ( .A(n8356), .B(n8355), .Z(n8428) );
  NANDN U8629 ( .A(n19394), .B(n8357), .Z(n8359) );
  XOR U8630 ( .A(b[29]), .B(a[43]), .Z(n8506) );
  NANDN U8631 ( .A(n19395), .B(n8506), .Z(n8358) );
  AND U8632 ( .A(n8359), .B(n8358), .Z(n8426) );
  AND U8633 ( .A(b[31]), .B(a[39]), .Z(n8425) );
  XNOR U8634 ( .A(n8426), .B(n8425), .Z(n8427) );
  XNOR U8635 ( .A(n8428), .B(n8427), .Z(n8467) );
  NANDN U8636 ( .A(n19005), .B(n8360), .Z(n8362) );
  XOR U8637 ( .A(b[23]), .B(a[49]), .Z(n8509) );
  NANDN U8638 ( .A(n19055), .B(n8509), .Z(n8361) );
  AND U8639 ( .A(n8362), .B(n8361), .Z(n8500) );
  NANDN U8640 ( .A(n17362), .B(n8363), .Z(n8365) );
  XOR U8641 ( .A(b[7]), .B(a[65]), .Z(n8512) );
  NANDN U8642 ( .A(n17522), .B(n8512), .Z(n8364) );
  AND U8643 ( .A(n8365), .B(n8364), .Z(n8498) );
  NANDN U8644 ( .A(n19116), .B(n8366), .Z(n8368) );
  XOR U8645 ( .A(b[25]), .B(a[47]), .Z(n8515) );
  NANDN U8646 ( .A(n19179), .B(n8515), .Z(n8367) );
  NAND U8647 ( .A(n8368), .B(n8367), .Z(n8497) );
  XNOR U8648 ( .A(n8498), .B(n8497), .Z(n8499) );
  XOR U8649 ( .A(n8500), .B(n8499), .Z(n8468) );
  XNOR U8650 ( .A(n8467), .B(n8468), .Z(n8469) );
  NANDN U8651 ( .A(n18113), .B(n8369), .Z(n8371) );
  XOR U8652 ( .A(b[13]), .B(a[59]), .Z(n8518) );
  NANDN U8653 ( .A(n18229), .B(n8518), .Z(n8370) );
  AND U8654 ( .A(n8371), .B(n8370), .Z(n8462) );
  NANDN U8655 ( .A(n17888), .B(n8372), .Z(n8374) );
  XOR U8656 ( .A(b[11]), .B(a[61]), .Z(n8521) );
  NANDN U8657 ( .A(n18025), .B(n8521), .Z(n8373) );
  NAND U8658 ( .A(n8374), .B(n8373), .Z(n8461) );
  XNOR U8659 ( .A(n8462), .B(n8461), .Z(n8463) );
  NANDN U8660 ( .A(n18487), .B(n8375), .Z(n8377) );
  XOR U8661 ( .A(b[15]), .B(a[57]), .Z(n8524) );
  NANDN U8662 ( .A(n18311), .B(n8524), .Z(n8376) );
  AND U8663 ( .A(n8377), .B(n8376), .Z(n8458) );
  NANDN U8664 ( .A(n18853), .B(n8378), .Z(n8380) );
  XOR U8665 ( .A(b[21]), .B(a[51]), .Z(n8527) );
  NANDN U8666 ( .A(n18926), .B(n8527), .Z(n8379) );
  AND U8667 ( .A(n8380), .B(n8379), .Z(n8456) );
  NANDN U8668 ( .A(n17613), .B(n8381), .Z(n8383) );
  XOR U8669 ( .A(b[9]), .B(a[63]), .Z(n8530) );
  NANDN U8670 ( .A(n17739), .B(n8530), .Z(n8382) );
  NAND U8671 ( .A(n8383), .B(n8382), .Z(n8455) );
  XNOR U8672 ( .A(n8456), .B(n8455), .Z(n8457) );
  XOR U8673 ( .A(n8458), .B(n8457), .Z(n8464) );
  XOR U8674 ( .A(n8463), .B(n8464), .Z(n8470) );
  XOR U8675 ( .A(n8469), .B(n8470), .Z(n8482) );
  XNOR U8676 ( .A(n8481), .B(n8482), .Z(n8413) );
  XNOR U8677 ( .A(n8414), .B(n8413), .Z(n8415) );
  XOR U8678 ( .A(n8416), .B(n8415), .Z(n8534) );
  XNOR U8679 ( .A(n8533), .B(n8534), .Z(n8535) );
  XNOR U8680 ( .A(n8536), .B(n8535), .Z(n8409) );
  XOR U8681 ( .A(n8410), .B(n8409), .Z(n8402) );
  NANDN U8682 ( .A(n8385), .B(n8384), .Z(n8389) );
  NANDN U8683 ( .A(n8387), .B(n8386), .Z(n8388) );
  AND U8684 ( .A(n8389), .B(n8388), .Z(n8401) );
  XOR U8685 ( .A(n8402), .B(n8401), .Z(n8404) );
  XNOR U8686 ( .A(n8403), .B(n8404), .Z(n8395) );
  XNOR U8687 ( .A(n8396), .B(n8395), .Z(n8397) );
  XNOR U8688 ( .A(n8398), .B(n8397), .Z(n8539) );
  XNOR U8689 ( .A(sreg[167]), .B(n8539), .Z(n8541) );
  NANDN U8690 ( .A(sreg[166]), .B(n8390), .Z(n8394) );
  NAND U8691 ( .A(n8392), .B(n8391), .Z(n8393) );
  NAND U8692 ( .A(n8394), .B(n8393), .Z(n8540) );
  XNOR U8693 ( .A(n8541), .B(n8540), .Z(c[167]) );
  NANDN U8694 ( .A(n8396), .B(n8395), .Z(n8400) );
  NANDN U8695 ( .A(n8398), .B(n8397), .Z(n8399) );
  AND U8696 ( .A(n8400), .B(n8399), .Z(n8547) );
  NANDN U8697 ( .A(n8402), .B(n8401), .Z(n8406) );
  NANDN U8698 ( .A(n8404), .B(n8403), .Z(n8405) );
  AND U8699 ( .A(n8406), .B(n8405), .Z(n8545) );
  NANDN U8700 ( .A(n8408), .B(n8407), .Z(n8412) );
  NAND U8701 ( .A(n8410), .B(n8409), .Z(n8411) );
  AND U8702 ( .A(n8412), .B(n8411), .Z(n8552) );
  NANDN U8703 ( .A(n8414), .B(n8413), .Z(n8418) );
  NANDN U8704 ( .A(n8416), .B(n8415), .Z(n8417) );
  AND U8705 ( .A(n8418), .B(n8417), .Z(n8557) );
  NANDN U8706 ( .A(n8420), .B(n8419), .Z(n8424) );
  NAND U8707 ( .A(n8422), .B(n8421), .Z(n8423) );
  AND U8708 ( .A(n8424), .B(n8423), .Z(n8556) );
  XNOR U8709 ( .A(n8557), .B(n8556), .Z(n8559) );
  NANDN U8710 ( .A(n8426), .B(n8425), .Z(n8430) );
  NANDN U8711 ( .A(n8428), .B(n8427), .Z(n8429) );
  AND U8712 ( .A(n8430), .B(n8429), .Z(n8636) );
  NANDN U8713 ( .A(n19237), .B(n8431), .Z(n8433) );
  XOR U8714 ( .A(b[27]), .B(a[46]), .Z(n8580) );
  NANDN U8715 ( .A(n19277), .B(n8580), .Z(n8432) );
  AND U8716 ( .A(n8433), .B(n8432), .Z(n8643) );
  NANDN U8717 ( .A(n17072), .B(n8434), .Z(n8436) );
  XOR U8718 ( .A(b[5]), .B(a[68]), .Z(n8583) );
  NANDN U8719 ( .A(n17223), .B(n8583), .Z(n8435) );
  AND U8720 ( .A(n8436), .B(n8435), .Z(n8641) );
  NANDN U8721 ( .A(n18673), .B(n8437), .Z(n8439) );
  XOR U8722 ( .A(b[19]), .B(a[54]), .Z(n8586) );
  NANDN U8723 ( .A(n18758), .B(n8586), .Z(n8438) );
  NAND U8724 ( .A(n8439), .B(n8438), .Z(n8640) );
  XNOR U8725 ( .A(n8641), .B(n8640), .Z(n8642) );
  XNOR U8726 ( .A(n8643), .B(n8642), .Z(n8634) );
  NANDN U8727 ( .A(n19425), .B(n8440), .Z(n8442) );
  XOR U8728 ( .A(b[31]), .B(a[42]), .Z(n8589) );
  NANDN U8729 ( .A(n19426), .B(n8589), .Z(n8441) );
  AND U8730 ( .A(n8442), .B(n8441), .Z(n8601) );
  NANDN U8731 ( .A(n17067), .B(n8443), .Z(n8445) );
  XOR U8732 ( .A(b[3]), .B(a[70]), .Z(n8592) );
  NANDN U8733 ( .A(n17068), .B(n8592), .Z(n8444) );
  AND U8734 ( .A(n8445), .B(n8444), .Z(n8599) );
  NANDN U8735 ( .A(n18514), .B(n8446), .Z(n8448) );
  XOR U8736 ( .A(b[17]), .B(a[56]), .Z(n8595) );
  NANDN U8737 ( .A(n18585), .B(n8595), .Z(n8447) );
  NAND U8738 ( .A(n8448), .B(n8447), .Z(n8598) );
  XNOR U8739 ( .A(n8599), .B(n8598), .Z(n8600) );
  XOR U8740 ( .A(n8601), .B(n8600), .Z(n8635) );
  XOR U8741 ( .A(n8634), .B(n8635), .Z(n8637) );
  XOR U8742 ( .A(n8636), .B(n8637), .Z(n8569) );
  NANDN U8743 ( .A(n8450), .B(n8449), .Z(n8454) );
  NANDN U8744 ( .A(n8452), .B(n8451), .Z(n8453) );
  AND U8745 ( .A(n8454), .B(n8453), .Z(n8622) );
  NANDN U8746 ( .A(n8456), .B(n8455), .Z(n8460) );
  NANDN U8747 ( .A(n8458), .B(n8457), .Z(n8459) );
  NAND U8748 ( .A(n8460), .B(n8459), .Z(n8623) );
  XNOR U8749 ( .A(n8622), .B(n8623), .Z(n8624) );
  NANDN U8750 ( .A(n8462), .B(n8461), .Z(n8466) );
  NANDN U8751 ( .A(n8464), .B(n8463), .Z(n8465) );
  NAND U8752 ( .A(n8466), .B(n8465), .Z(n8625) );
  XNOR U8753 ( .A(n8624), .B(n8625), .Z(n8568) );
  XNOR U8754 ( .A(n8569), .B(n8568), .Z(n8571) );
  NANDN U8755 ( .A(n8468), .B(n8467), .Z(n8472) );
  NANDN U8756 ( .A(n8470), .B(n8469), .Z(n8471) );
  AND U8757 ( .A(n8472), .B(n8471), .Z(n8570) );
  XOR U8758 ( .A(n8571), .B(n8570), .Z(n8685) );
  NANDN U8759 ( .A(n8474), .B(n8473), .Z(n8478) );
  NANDN U8760 ( .A(n8476), .B(n8475), .Z(n8477) );
  AND U8761 ( .A(n8478), .B(n8477), .Z(n8682) );
  NANDN U8762 ( .A(n8480), .B(n8479), .Z(n8484) );
  NANDN U8763 ( .A(n8482), .B(n8481), .Z(n8483) );
  AND U8764 ( .A(n8484), .B(n8483), .Z(n8565) );
  NANDN U8765 ( .A(n8486), .B(n8485), .Z(n8490) );
  OR U8766 ( .A(n8488), .B(n8487), .Z(n8489) );
  AND U8767 ( .A(n8490), .B(n8489), .Z(n8563) );
  NANDN U8768 ( .A(n8492), .B(n8491), .Z(n8496) );
  NANDN U8769 ( .A(n8494), .B(n8493), .Z(n8495) );
  AND U8770 ( .A(n8496), .B(n8495), .Z(n8629) );
  NANDN U8771 ( .A(n8498), .B(n8497), .Z(n8502) );
  NANDN U8772 ( .A(n8500), .B(n8499), .Z(n8501) );
  NAND U8773 ( .A(n8502), .B(n8501), .Z(n8628) );
  XNOR U8774 ( .A(n8629), .B(n8628), .Z(n8630) );
  NAND U8775 ( .A(b[0]), .B(a[72]), .Z(n8503) );
  XNOR U8776 ( .A(b[1]), .B(n8503), .Z(n8505) );
  NANDN U8777 ( .A(b[0]), .B(a[71]), .Z(n8504) );
  NAND U8778 ( .A(n8505), .B(n8504), .Z(n8577) );
  NANDN U8779 ( .A(n19394), .B(n8506), .Z(n8508) );
  XOR U8780 ( .A(b[29]), .B(a[44]), .Z(n8655) );
  NANDN U8781 ( .A(n19395), .B(n8655), .Z(n8507) );
  AND U8782 ( .A(n8508), .B(n8507), .Z(n8575) );
  AND U8783 ( .A(b[31]), .B(a[40]), .Z(n8574) );
  XNOR U8784 ( .A(n8575), .B(n8574), .Z(n8576) );
  XNOR U8785 ( .A(n8577), .B(n8576), .Z(n8616) );
  NANDN U8786 ( .A(n19005), .B(n8509), .Z(n8511) );
  XOR U8787 ( .A(b[23]), .B(a[50]), .Z(n8658) );
  NANDN U8788 ( .A(n19055), .B(n8658), .Z(n8510) );
  AND U8789 ( .A(n8511), .B(n8510), .Z(n8649) );
  NANDN U8790 ( .A(n17362), .B(n8512), .Z(n8514) );
  XOR U8791 ( .A(b[7]), .B(a[66]), .Z(n8661) );
  NANDN U8792 ( .A(n17522), .B(n8661), .Z(n8513) );
  AND U8793 ( .A(n8514), .B(n8513), .Z(n8647) );
  NANDN U8794 ( .A(n19116), .B(n8515), .Z(n8517) );
  XOR U8795 ( .A(b[25]), .B(a[48]), .Z(n8664) );
  NANDN U8796 ( .A(n19179), .B(n8664), .Z(n8516) );
  NAND U8797 ( .A(n8517), .B(n8516), .Z(n8646) );
  XNOR U8798 ( .A(n8647), .B(n8646), .Z(n8648) );
  XOR U8799 ( .A(n8649), .B(n8648), .Z(n8617) );
  XNOR U8800 ( .A(n8616), .B(n8617), .Z(n8618) );
  NANDN U8801 ( .A(n18113), .B(n8518), .Z(n8520) );
  XOR U8802 ( .A(b[13]), .B(a[60]), .Z(n8667) );
  NANDN U8803 ( .A(n18229), .B(n8667), .Z(n8519) );
  AND U8804 ( .A(n8520), .B(n8519), .Z(n8611) );
  NANDN U8805 ( .A(n17888), .B(n8521), .Z(n8523) );
  XOR U8806 ( .A(b[11]), .B(a[62]), .Z(n8670) );
  NANDN U8807 ( .A(n18025), .B(n8670), .Z(n8522) );
  NAND U8808 ( .A(n8523), .B(n8522), .Z(n8610) );
  XNOR U8809 ( .A(n8611), .B(n8610), .Z(n8612) );
  NANDN U8810 ( .A(n18487), .B(n8524), .Z(n8526) );
  XOR U8811 ( .A(b[15]), .B(a[58]), .Z(n8673) );
  NANDN U8812 ( .A(n18311), .B(n8673), .Z(n8525) );
  AND U8813 ( .A(n8526), .B(n8525), .Z(n8607) );
  NANDN U8814 ( .A(n18853), .B(n8527), .Z(n8529) );
  XOR U8815 ( .A(b[21]), .B(a[52]), .Z(n8676) );
  NANDN U8816 ( .A(n18926), .B(n8676), .Z(n8528) );
  AND U8817 ( .A(n8529), .B(n8528), .Z(n8605) );
  NANDN U8818 ( .A(n17613), .B(n8530), .Z(n8532) );
  XOR U8819 ( .A(b[9]), .B(a[64]), .Z(n8679) );
  NANDN U8820 ( .A(n17739), .B(n8679), .Z(n8531) );
  NAND U8821 ( .A(n8532), .B(n8531), .Z(n8604) );
  XNOR U8822 ( .A(n8605), .B(n8604), .Z(n8606) );
  XOR U8823 ( .A(n8607), .B(n8606), .Z(n8613) );
  XOR U8824 ( .A(n8612), .B(n8613), .Z(n8619) );
  XOR U8825 ( .A(n8618), .B(n8619), .Z(n8631) );
  XNOR U8826 ( .A(n8630), .B(n8631), .Z(n8562) );
  XNOR U8827 ( .A(n8563), .B(n8562), .Z(n8564) );
  XOR U8828 ( .A(n8565), .B(n8564), .Z(n8683) );
  XNOR U8829 ( .A(n8682), .B(n8683), .Z(n8684) );
  XNOR U8830 ( .A(n8685), .B(n8684), .Z(n8558) );
  XOR U8831 ( .A(n8559), .B(n8558), .Z(n8551) );
  NANDN U8832 ( .A(n8534), .B(n8533), .Z(n8538) );
  NANDN U8833 ( .A(n8536), .B(n8535), .Z(n8537) );
  AND U8834 ( .A(n8538), .B(n8537), .Z(n8550) );
  XOR U8835 ( .A(n8551), .B(n8550), .Z(n8553) );
  XNOR U8836 ( .A(n8552), .B(n8553), .Z(n8544) );
  XNOR U8837 ( .A(n8545), .B(n8544), .Z(n8546) );
  XNOR U8838 ( .A(n8547), .B(n8546), .Z(n8688) );
  XNOR U8839 ( .A(sreg[168]), .B(n8688), .Z(n8690) );
  NANDN U8840 ( .A(sreg[167]), .B(n8539), .Z(n8543) );
  NAND U8841 ( .A(n8541), .B(n8540), .Z(n8542) );
  NAND U8842 ( .A(n8543), .B(n8542), .Z(n8689) );
  XNOR U8843 ( .A(n8690), .B(n8689), .Z(c[168]) );
  NANDN U8844 ( .A(n8545), .B(n8544), .Z(n8549) );
  NANDN U8845 ( .A(n8547), .B(n8546), .Z(n8548) );
  AND U8846 ( .A(n8549), .B(n8548), .Z(n8696) );
  NANDN U8847 ( .A(n8551), .B(n8550), .Z(n8555) );
  NANDN U8848 ( .A(n8553), .B(n8552), .Z(n8554) );
  AND U8849 ( .A(n8555), .B(n8554), .Z(n8694) );
  NANDN U8850 ( .A(n8557), .B(n8556), .Z(n8561) );
  NAND U8851 ( .A(n8559), .B(n8558), .Z(n8560) );
  AND U8852 ( .A(n8561), .B(n8560), .Z(n8701) );
  NANDN U8853 ( .A(n8563), .B(n8562), .Z(n8567) );
  NANDN U8854 ( .A(n8565), .B(n8564), .Z(n8566) );
  AND U8855 ( .A(n8567), .B(n8566), .Z(n8706) );
  NANDN U8856 ( .A(n8569), .B(n8568), .Z(n8573) );
  NAND U8857 ( .A(n8571), .B(n8570), .Z(n8572) );
  AND U8858 ( .A(n8573), .B(n8572), .Z(n8705) );
  XNOR U8859 ( .A(n8706), .B(n8705), .Z(n8708) );
  NANDN U8860 ( .A(n8575), .B(n8574), .Z(n8579) );
  NANDN U8861 ( .A(n8577), .B(n8576), .Z(n8578) );
  AND U8862 ( .A(n8579), .B(n8578), .Z(n8785) );
  NANDN U8863 ( .A(n19237), .B(n8580), .Z(n8582) );
  XOR U8864 ( .A(b[27]), .B(a[47]), .Z(n8729) );
  NANDN U8865 ( .A(n19277), .B(n8729), .Z(n8581) );
  AND U8866 ( .A(n8582), .B(n8581), .Z(n8792) );
  NANDN U8867 ( .A(n17072), .B(n8583), .Z(n8585) );
  XOR U8868 ( .A(b[5]), .B(a[69]), .Z(n8732) );
  NANDN U8869 ( .A(n17223), .B(n8732), .Z(n8584) );
  AND U8870 ( .A(n8585), .B(n8584), .Z(n8790) );
  NANDN U8871 ( .A(n18673), .B(n8586), .Z(n8588) );
  XOR U8872 ( .A(b[19]), .B(a[55]), .Z(n8735) );
  NANDN U8873 ( .A(n18758), .B(n8735), .Z(n8587) );
  NAND U8874 ( .A(n8588), .B(n8587), .Z(n8789) );
  XNOR U8875 ( .A(n8790), .B(n8789), .Z(n8791) );
  XNOR U8876 ( .A(n8792), .B(n8791), .Z(n8783) );
  NANDN U8877 ( .A(n19425), .B(n8589), .Z(n8591) );
  XOR U8878 ( .A(b[31]), .B(a[43]), .Z(n8738) );
  NANDN U8879 ( .A(n19426), .B(n8738), .Z(n8590) );
  AND U8880 ( .A(n8591), .B(n8590), .Z(n8750) );
  NANDN U8881 ( .A(n17067), .B(n8592), .Z(n8594) );
  XOR U8882 ( .A(b[3]), .B(a[71]), .Z(n8741) );
  NANDN U8883 ( .A(n17068), .B(n8741), .Z(n8593) );
  AND U8884 ( .A(n8594), .B(n8593), .Z(n8748) );
  NANDN U8885 ( .A(n18514), .B(n8595), .Z(n8597) );
  XOR U8886 ( .A(b[17]), .B(a[57]), .Z(n8744) );
  NANDN U8887 ( .A(n18585), .B(n8744), .Z(n8596) );
  NAND U8888 ( .A(n8597), .B(n8596), .Z(n8747) );
  XNOR U8889 ( .A(n8748), .B(n8747), .Z(n8749) );
  XOR U8890 ( .A(n8750), .B(n8749), .Z(n8784) );
  XOR U8891 ( .A(n8783), .B(n8784), .Z(n8786) );
  XOR U8892 ( .A(n8785), .B(n8786), .Z(n8718) );
  NANDN U8893 ( .A(n8599), .B(n8598), .Z(n8603) );
  NANDN U8894 ( .A(n8601), .B(n8600), .Z(n8602) );
  AND U8895 ( .A(n8603), .B(n8602), .Z(n8771) );
  NANDN U8896 ( .A(n8605), .B(n8604), .Z(n8609) );
  NANDN U8897 ( .A(n8607), .B(n8606), .Z(n8608) );
  NAND U8898 ( .A(n8609), .B(n8608), .Z(n8772) );
  XNOR U8899 ( .A(n8771), .B(n8772), .Z(n8773) );
  NANDN U8900 ( .A(n8611), .B(n8610), .Z(n8615) );
  NANDN U8901 ( .A(n8613), .B(n8612), .Z(n8614) );
  NAND U8902 ( .A(n8615), .B(n8614), .Z(n8774) );
  XNOR U8903 ( .A(n8773), .B(n8774), .Z(n8717) );
  XNOR U8904 ( .A(n8718), .B(n8717), .Z(n8720) );
  NANDN U8905 ( .A(n8617), .B(n8616), .Z(n8621) );
  NANDN U8906 ( .A(n8619), .B(n8618), .Z(n8620) );
  AND U8907 ( .A(n8621), .B(n8620), .Z(n8719) );
  XOR U8908 ( .A(n8720), .B(n8719), .Z(n8834) );
  NANDN U8909 ( .A(n8623), .B(n8622), .Z(n8627) );
  NANDN U8910 ( .A(n8625), .B(n8624), .Z(n8626) );
  AND U8911 ( .A(n8627), .B(n8626), .Z(n8831) );
  NANDN U8912 ( .A(n8629), .B(n8628), .Z(n8633) );
  NANDN U8913 ( .A(n8631), .B(n8630), .Z(n8632) );
  AND U8914 ( .A(n8633), .B(n8632), .Z(n8714) );
  NANDN U8915 ( .A(n8635), .B(n8634), .Z(n8639) );
  OR U8916 ( .A(n8637), .B(n8636), .Z(n8638) );
  AND U8917 ( .A(n8639), .B(n8638), .Z(n8712) );
  NANDN U8918 ( .A(n8641), .B(n8640), .Z(n8645) );
  NANDN U8919 ( .A(n8643), .B(n8642), .Z(n8644) );
  AND U8920 ( .A(n8645), .B(n8644), .Z(n8778) );
  NANDN U8921 ( .A(n8647), .B(n8646), .Z(n8651) );
  NANDN U8922 ( .A(n8649), .B(n8648), .Z(n8650) );
  NAND U8923 ( .A(n8651), .B(n8650), .Z(n8777) );
  XNOR U8924 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U8925 ( .A(b[0]), .B(a[73]), .Z(n8652) );
  XNOR U8926 ( .A(b[1]), .B(n8652), .Z(n8654) );
  NANDN U8927 ( .A(b[0]), .B(a[72]), .Z(n8653) );
  NAND U8928 ( .A(n8654), .B(n8653), .Z(n8726) );
  NANDN U8929 ( .A(n19394), .B(n8655), .Z(n8657) );
  XOR U8930 ( .A(b[29]), .B(a[45]), .Z(n8801) );
  NANDN U8931 ( .A(n19395), .B(n8801), .Z(n8656) );
  AND U8932 ( .A(n8657), .B(n8656), .Z(n8724) );
  AND U8933 ( .A(b[31]), .B(a[41]), .Z(n8723) );
  XNOR U8934 ( .A(n8724), .B(n8723), .Z(n8725) );
  XNOR U8935 ( .A(n8726), .B(n8725), .Z(n8765) );
  NANDN U8936 ( .A(n19005), .B(n8658), .Z(n8660) );
  XOR U8937 ( .A(b[23]), .B(a[51]), .Z(n8807) );
  NANDN U8938 ( .A(n19055), .B(n8807), .Z(n8659) );
  AND U8939 ( .A(n8660), .B(n8659), .Z(n8798) );
  NANDN U8940 ( .A(n17362), .B(n8661), .Z(n8663) );
  XOR U8941 ( .A(b[7]), .B(a[67]), .Z(n8810) );
  NANDN U8942 ( .A(n17522), .B(n8810), .Z(n8662) );
  AND U8943 ( .A(n8663), .B(n8662), .Z(n8796) );
  NANDN U8944 ( .A(n19116), .B(n8664), .Z(n8666) );
  XOR U8945 ( .A(b[25]), .B(a[49]), .Z(n8813) );
  NANDN U8946 ( .A(n19179), .B(n8813), .Z(n8665) );
  NAND U8947 ( .A(n8666), .B(n8665), .Z(n8795) );
  XNOR U8948 ( .A(n8796), .B(n8795), .Z(n8797) );
  XOR U8949 ( .A(n8798), .B(n8797), .Z(n8766) );
  XNOR U8950 ( .A(n8765), .B(n8766), .Z(n8767) );
  NANDN U8951 ( .A(n18113), .B(n8667), .Z(n8669) );
  XOR U8952 ( .A(b[13]), .B(a[61]), .Z(n8816) );
  NANDN U8953 ( .A(n18229), .B(n8816), .Z(n8668) );
  AND U8954 ( .A(n8669), .B(n8668), .Z(n8760) );
  NANDN U8955 ( .A(n17888), .B(n8670), .Z(n8672) );
  XOR U8956 ( .A(b[11]), .B(a[63]), .Z(n8819) );
  NANDN U8957 ( .A(n18025), .B(n8819), .Z(n8671) );
  NAND U8958 ( .A(n8672), .B(n8671), .Z(n8759) );
  XNOR U8959 ( .A(n8760), .B(n8759), .Z(n8761) );
  NANDN U8960 ( .A(n18487), .B(n8673), .Z(n8675) );
  XOR U8961 ( .A(b[15]), .B(a[59]), .Z(n8822) );
  NANDN U8962 ( .A(n18311), .B(n8822), .Z(n8674) );
  AND U8963 ( .A(n8675), .B(n8674), .Z(n8756) );
  NANDN U8964 ( .A(n18853), .B(n8676), .Z(n8678) );
  XOR U8965 ( .A(b[21]), .B(a[53]), .Z(n8825) );
  NANDN U8966 ( .A(n18926), .B(n8825), .Z(n8677) );
  AND U8967 ( .A(n8678), .B(n8677), .Z(n8754) );
  NANDN U8968 ( .A(n17613), .B(n8679), .Z(n8681) );
  XOR U8969 ( .A(b[9]), .B(a[65]), .Z(n8828) );
  NANDN U8970 ( .A(n17739), .B(n8828), .Z(n8680) );
  NAND U8971 ( .A(n8681), .B(n8680), .Z(n8753) );
  XNOR U8972 ( .A(n8754), .B(n8753), .Z(n8755) );
  XOR U8973 ( .A(n8756), .B(n8755), .Z(n8762) );
  XOR U8974 ( .A(n8761), .B(n8762), .Z(n8768) );
  XOR U8975 ( .A(n8767), .B(n8768), .Z(n8780) );
  XNOR U8976 ( .A(n8779), .B(n8780), .Z(n8711) );
  XNOR U8977 ( .A(n8712), .B(n8711), .Z(n8713) );
  XOR U8978 ( .A(n8714), .B(n8713), .Z(n8832) );
  XNOR U8979 ( .A(n8831), .B(n8832), .Z(n8833) );
  XNOR U8980 ( .A(n8834), .B(n8833), .Z(n8707) );
  XOR U8981 ( .A(n8708), .B(n8707), .Z(n8700) );
  NANDN U8982 ( .A(n8683), .B(n8682), .Z(n8687) );
  NANDN U8983 ( .A(n8685), .B(n8684), .Z(n8686) );
  AND U8984 ( .A(n8687), .B(n8686), .Z(n8699) );
  XOR U8985 ( .A(n8700), .B(n8699), .Z(n8702) );
  XNOR U8986 ( .A(n8701), .B(n8702), .Z(n8693) );
  XNOR U8987 ( .A(n8694), .B(n8693), .Z(n8695) );
  XNOR U8988 ( .A(n8696), .B(n8695), .Z(n8837) );
  XNOR U8989 ( .A(sreg[169]), .B(n8837), .Z(n8839) );
  NANDN U8990 ( .A(sreg[168]), .B(n8688), .Z(n8692) );
  NAND U8991 ( .A(n8690), .B(n8689), .Z(n8691) );
  NAND U8992 ( .A(n8692), .B(n8691), .Z(n8838) );
  XNOR U8993 ( .A(n8839), .B(n8838), .Z(c[169]) );
  NANDN U8994 ( .A(n8694), .B(n8693), .Z(n8698) );
  NANDN U8995 ( .A(n8696), .B(n8695), .Z(n8697) );
  AND U8996 ( .A(n8698), .B(n8697), .Z(n8845) );
  NANDN U8997 ( .A(n8700), .B(n8699), .Z(n8704) );
  NANDN U8998 ( .A(n8702), .B(n8701), .Z(n8703) );
  AND U8999 ( .A(n8704), .B(n8703), .Z(n8843) );
  NANDN U9000 ( .A(n8706), .B(n8705), .Z(n8710) );
  NAND U9001 ( .A(n8708), .B(n8707), .Z(n8709) );
  AND U9002 ( .A(n8710), .B(n8709), .Z(n8850) );
  NANDN U9003 ( .A(n8712), .B(n8711), .Z(n8716) );
  NANDN U9004 ( .A(n8714), .B(n8713), .Z(n8715) );
  AND U9005 ( .A(n8716), .B(n8715), .Z(n8855) );
  NANDN U9006 ( .A(n8718), .B(n8717), .Z(n8722) );
  NAND U9007 ( .A(n8720), .B(n8719), .Z(n8721) );
  AND U9008 ( .A(n8722), .B(n8721), .Z(n8854) );
  XNOR U9009 ( .A(n8855), .B(n8854), .Z(n8857) );
  NANDN U9010 ( .A(n8724), .B(n8723), .Z(n8728) );
  NANDN U9011 ( .A(n8726), .B(n8725), .Z(n8727) );
  AND U9012 ( .A(n8728), .B(n8727), .Z(n8934) );
  NANDN U9013 ( .A(n19237), .B(n8729), .Z(n8731) );
  XOR U9014 ( .A(b[27]), .B(a[48]), .Z(n8878) );
  NANDN U9015 ( .A(n19277), .B(n8878), .Z(n8730) );
  AND U9016 ( .A(n8731), .B(n8730), .Z(n8941) );
  NANDN U9017 ( .A(n17072), .B(n8732), .Z(n8734) );
  XOR U9018 ( .A(b[5]), .B(a[70]), .Z(n8881) );
  NANDN U9019 ( .A(n17223), .B(n8881), .Z(n8733) );
  AND U9020 ( .A(n8734), .B(n8733), .Z(n8939) );
  NANDN U9021 ( .A(n18673), .B(n8735), .Z(n8737) );
  XOR U9022 ( .A(b[19]), .B(a[56]), .Z(n8884) );
  NANDN U9023 ( .A(n18758), .B(n8884), .Z(n8736) );
  NAND U9024 ( .A(n8737), .B(n8736), .Z(n8938) );
  XNOR U9025 ( .A(n8939), .B(n8938), .Z(n8940) );
  XNOR U9026 ( .A(n8941), .B(n8940), .Z(n8932) );
  NANDN U9027 ( .A(n19425), .B(n8738), .Z(n8740) );
  XOR U9028 ( .A(b[31]), .B(a[44]), .Z(n8887) );
  NANDN U9029 ( .A(n19426), .B(n8887), .Z(n8739) );
  AND U9030 ( .A(n8740), .B(n8739), .Z(n8899) );
  NANDN U9031 ( .A(n17067), .B(n8741), .Z(n8743) );
  XOR U9032 ( .A(b[3]), .B(a[72]), .Z(n8890) );
  NANDN U9033 ( .A(n17068), .B(n8890), .Z(n8742) );
  AND U9034 ( .A(n8743), .B(n8742), .Z(n8897) );
  NANDN U9035 ( .A(n18514), .B(n8744), .Z(n8746) );
  XOR U9036 ( .A(b[17]), .B(a[58]), .Z(n8893) );
  NANDN U9037 ( .A(n18585), .B(n8893), .Z(n8745) );
  NAND U9038 ( .A(n8746), .B(n8745), .Z(n8896) );
  XNOR U9039 ( .A(n8897), .B(n8896), .Z(n8898) );
  XOR U9040 ( .A(n8899), .B(n8898), .Z(n8933) );
  XOR U9041 ( .A(n8932), .B(n8933), .Z(n8935) );
  XOR U9042 ( .A(n8934), .B(n8935), .Z(n8867) );
  NANDN U9043 ( .A(n8748), .B(n8747), .Z(n8752) );
  NANDN U9044 ( .A(n8750), .B(n8749), .Z(n8751) );
  AND U9045 ( .A(n8752), .B(n8751), .Z(n8920) );
  NANDN U9046 ( .A(n8754), .B(n8753), .Z(n8758) );
  NANDN U9047 ( .A(n8756), .B(n8755), .Z(n8757) );
  NAND U9048 ( .A(n8758), .B(n8757), .Z(n8921) );
  XNOR U9049 ( .A(n8920), .B(n8921), .Z(n8922) );
  NANDN U9050 ( .A(n8760), .B(n8759), .Z(n8764) );
  NANDN U9051 ( .A(n8762), .B(n8761), .Z(n8763) );
  NAND U9052 ( .A(n8764), .B(n8763), .Z(n8923) );
  XNOR U9053 ( .A(n8922), .B(n8923), .Z(n8866) );
  XNOR U9054 ( .A(n8867), .B(n8866), .Z(n8869) );
  NANDN U9055 ( .A(n8766), .B(n8765), .Z(n8770) );
  NANDN U9056 ( .A(n8768), .B(n8767), .Z(n8769) );
  AND U9057 ( .A(n8770), .B(n8769), .Z(n8868) );
  XOR U9058 ( .A(n8869), .B(n8868), .Z(n8983) );
  NANDN U9059 ( .A(n8772), .B(n8771), .Z(n8776) );
  NANDN U9060 ( .A(n8774), .B(n8773), .Z(n8775) );
  AND U9061 ( .A(n8776), .B(n8775), .Z(n8980) );
  NANDN U9062 ( .A(n8778), .B(n8777), .Z(n8782) );
  NANDN U9063 ( .A(n8780), .B(n8779), .Z(n8781) );
  AND U9064 ( .A(n8782), .B(n8781), .Z(n8863) );
  NANDN U9065 ( .A(n8784), .B(n8783), .Z(n8788) );
  OR U9066 ( .A(n8786), .B(n8785), .Z(n8787) );
  AND U9067 ( .A(n8788), .B(n8787), .Z(n8861) );
  NANDN U9068 ( .A(n8790), .B(n8789), .Z(n8794) );
  NANDN U9069 ( .A(n8792), .B(n8791), .Z(n8793) );
  AND U9070 ( .A(n8794), .B(n8793), .Z(n8927) );
  NANDN U9071 ( .A(n8796), .B(n8795), .Z(n8800) );
  NANDN U9072 ( .A(n8798), .B(n8797), .Z(n8799) );
  NAND U9073 ( .A(n8800), .B(n8799), .Z(n8926) );
  XNOR U9074 ( .A(n8927), .B(n8926), .Z(n8928) );
  NANDN U9075 ( .A(n19394), .B(n8801), .Z(n8803) );
  XOR U9076 ( .A(b[29]), .B(a[46]), .Z(n8953) );
  NANDN U9077 ( .A(n19395), .B(n8953), .Z(n8802) );
  AND U9078 ( .A(n8803), .B(n8802), .Z(n8873) );
  AND U9079 ( .A(b[31]), .B(a[42]), .Z(n8872) );
  XNOR U9080 ( .A(n8873), .B(n8872), .Z(n8874) );
  NAND U9081 ( .A(b[0]), .B(a[74]), .Z(n8804) );
  XNOR U9082 ( .A(b[1]), .B(n8804), .Z(n8806) );
  NANDN U9083 ( .A(b[0]), .B(a[73]), .Z(n8805) );
  NAND U9084 ( .A(n8806), .B(n8805), .Z(n8875) );
  XNOR U9085 ( .A(n8874), .B(n8875), .Z(n8914) );
  NANDN U9086 ( .A(n19005), .B(n8807), .Z(n8809) );
  XOR U9087 ( .A(b[23]), .B(a[52]), .Z(n8956) );
  NANDN U9088 ( .A(n19055), .B(n8956), .Z(n8808) );
  AND U9089 ( .A(n8809), .B(n8808), .Z(n8947) );
  NANDN U9090 ( .A(n17362), .B(n8810), .Z(n8812) );
  XOR U9091 ( .A(b[7]), .B(a[68]), .Z(n8959) );
  NANDN U9092 ( .A(n17522), .B(n8959), .Z(n8811) );
  AND U9093 ( .A(n8812), .B(n8811), .Z(n8945) );
  NANDN U9094 ( .A(n19116), .B(n8813), .Z(n8815) );
  XOR U9095 ( .A(b[25]), .B(a[50]), .Z(n8962) );
  NANDN U9096 ( .A(n19179), .B(n8962), .Z(n8814) );
  NAND U9097 ( .A(n8815), .B(n8814), .Z(n8944) );
  XNOR U9098 ( .A(n8945), .B(n8944), .Z(n8946) );
  XOR U9099 ( .A(n8947), .B(n8946), .Z(n8915) );
  XNOR U9100 ( .A(n8914), .B(n8915), .Z(n8916) );
  NANDN U9101 ( .A(n18113), .B(n8816), .Z(n8818) );
  XOR U9102 ( .A(b[13]), .B(a[62]), .Z(n8965) );
  NANDN U9103 ( .A(n18229), .B(n8965), .Z(n8817) );
  AND U9104 ( .A(n8818), .B(n8817), .Z(n8909) );
  NANDN U9105 ( .A(n17888), .B(n8819), .Z(n8821) );
  XOR U9106 ( .A(b[11]), .B(a[64]), .Z(n8968) );
  NANDN U9107 ( .A(n18025), .B(n8968), .Z(n8820) );
  NAND U9108 ( .A(n8821), .B(n8820), .Z(n8908) );
  XNOR U9109 ( .A(n8909), .B(n8908), .Z(n8910) );
  NANDN U9110 ( .A(n18487), .B(n8822), .Z(n8824) );
  XOR U9111 ( .A(b[15]), .B(a[60]), .Z(n8971) );
  NANDN U9112 ( .A(n18311), .B(n8971), .Z(n8823) );
  AND U9113 ( .A(n8824), .B(n8823), .Z(n8905) );
  NANDN U9114 ( .A(n18853), .B(n8825), .Z(n8827) );
  XOR U9115 ( .A(b[21]), .B(a[54]), .Z(n8974) );
  NANDN U9116 ( .A(n18926), .B(n8974), .Z(n8826) );
  AND U9117 ( .A(n8827), .B(n8826), .Z(n8903) );
  NANDN U9118 ( .A(n17613), .B(n8828), .Z(n8830) );
  XOR U9119 ( .A(b[9]), .B(a[66]), .Z(n8977) );
  NANDN U9120 ( .A(n17739), .B(n8977), .Z(n8829) );
  NAND U9121 ( .A(n8830), .B(n8829), .Z(n8902) );
  XNOR U9122 ( .A(n8903), .B(n8902), .Z(n8904) );
  XOR U9123 ( .A(n8905), .B(n8904), .Z(n8911) );
  XOR U9124 ( .A(n8910), .B(n8911), .Z(n8917) );
  XOR U9125 ( .A(n8916), .B(n8917), .Z(n8929) );
  XNOR U9126 ( .A(n8928), .B(n8929), .Z(n8860) );
  XNOR U9127 ( .A(n8861), .B(n8860), .Z(n8862) );
  XOR U9128 ( .A(n8863), .B(n8862), .Z(n8981) );
  XNOR U9129 ( .A(n8980), .B(n8981), .Z(n8982) );
  XNOR U9130 ( .A(n8983), .B(n8982), .Z(n8856) );
  XOR U9131 ( .A(n8857), .B(n8856), .Z(n8849) );
  NANDN U9132 ( .A(n8832), .B(n8831), .Z(n8836) );
  NANDN U9133 ( .A(n8834), .B(n8833), .Z(n8835) );
  AND U9134 ( .A(n8836), .B(n8835), .Z(n8848) );
  XOR U9135 ( .A(n8849), .B(n8848), .Z(n8851) );
  XNOR U9136 ( .A(n8850), .B(n8851), .Z(n8842) );
  XNOR U9137 ( .A(n8843), .B(n8842), .Z(n8844) );
  XNOR U9138 ( .A(n8845), .B(n8844), .Z(n8986) );
  XNOR U9139 ( .A(sreg[170]), .B(n8986), .Z(n8988) );
  NANDN U9140 ( .A(sreg[169]), .B(n8837), .Z(n8841) );
  NAND U9141 ( .A(n8839), .B(n8838), .Z(n8840) );
  NAND U9142 ( .A(n8841), .B(n8840), .Z(n8987) );
  XNOR U9143 ( .A(n8988), .B(n8987), .Z(c[170]) );
  NANDN U9144 ( .A(n8843), .B(n8842), .Z(n8847) );
  NANDN U9145 ( .A(n8845), .B(n8844), .Z(n8846) );
  AND U9146 ( .A(n8847), .B(n8846), .Z(n8994) );
  NANDN U9147 ( .A(n8849), .B(n8848), .Z(n8853) );
  NANDN U9148 ( .A(n8851), .B(n8850), .Z(n8852) );
  AND U9149 ( .A(n8853), .B(n8852), .Z(n8992) );
  NANDN U9150 ( .A(n8855), .B(n8854), .Z(n8859) );
  NAND U9151 ( .A(n8857), .B(n8856), .Z(n8858) );
  AND U9152 ( .A(n8859), .B(n8858), .Z(n8999) );
  NANDN U9153 ( .A(n8861), .B(n8860), .Z(n8865) );
  NANDN U9154 ( .A(n8863), .B(n8862), .Z(n8864) );
  AND U9155 ( .A(n8865), .B(n8864), .Z(n9004) );
  NANDN U9156 ( .A(n8867), .B(n8866), .Z(n8871) );
  NAND U9157 ( .A(n8869), .B(n8868), .Z(n8870) );
  AND U9158 ( .A(n8871), .B(n8870), .Z(n9003) );
  XNOR U9159 ( .A(n9004), .B(n9003), .Z(n9006) );
  NANDN U9160 ( .A(n8873), .B(n8872), .Z(n8877) );
  NANDN U9161 ( .A(n8875), .B(n8874), .Z(n8876) );
  AND U9162 ( .A(n8877), .B(n8876), .Z(n9083) );
  NANDN U9163 ( .A(n19237), .B(n8878), .Z(n8880) );
  XOR U9164 ( .A(b[27]), .B(a[49]), .Z(n9027) );
  NANDN U9165 ( .A(n19277), .B(n9027), .Z(n8879) );
  AND U9166 ( .A(n8880), .B(n8879), .Z(n9090) );
  NANDN U9167 ( .A(n17072), .B(n8881), .Z(n8883) );
  XOR U9168 ( .A(b[5]), .B(a[71]), .Z(n9030) );
  NANDN U9169 ( .A(n17223), .B(n9030), .Z(n8882) );
  AND U9170 ( .A(n8883), .B(n8882), .Z(n9088) );
  NANDN U9171 ( .A(n18673), .B(n8884), .Z(n8886) );
  XOR U9172 ( .A(b[19]), .B(a[57]), .Z(n9033) );
  NANDN U9173 ( .A(n18758), .B(n9033), .Z(n8885) );
  NAND U9174 ( .A(n8886), .B(n8885), .Z(n9087) );
  XNOR U9175 ( .A(n9088), .B(n9087), .Z(n9089) );
  XNOR U9176 ( .A(n9090), .B(n9089), .Z(n9081) );
  NANDN U9177 ( .A(n19425), .B(n8887), .Z(n8889) );
  XOR U9178 ( .A(b[31]), .B(a[45]), .Z(n9036) );
  NANDN U9179 ( .A(n19426), .B(n9036), .Z(n8888) );
  AND U9180 ( .A(n8889), .B(n8888), .Z(n9048) );
  NANDN U9181 ( .A(n17067), .B(n8890), .Z(n8892) );
  XOR U9182 ( .A(b[3]), .B(a[73]), .Z(n9039) );
  NANDN U9183 ( .A(n17068), .B(n9039), .Z(n8891) );
  AND U9184 ( .A(n8892), .B(n8891), .Z(n9046) );
  NANDN U9185 ( .A(n18514), .B(n8893), .Z(n8895) );
  XOR U9186 ( .A(b[17]), .B(a[59]), .Z(n9042) );
  NANDN U9187 ( .A(n18585), .B(n9042), .Z(n8894) );
  NAND U9188 ( .A(n8895), .B(n8894), .Z(n9045) );
  XNOR U9189 ( .A(n9046), .B(n9045), .Z(n9047) );
  XOR U9190 ( .A(n9048), .B(n9047), .Z(n9082) );
  XOR U9191 ( .A(n9081), .B(n9082), .Z(n9084) );
  XOR U9192 ( .A(n9083), .B(n9084), .Z(n9016) );
  NANDN U9193 ( .A(n8897), .B(n8896), .Z(n8901) );
  NANDN U9194 ( .A(n8899), .B(n8898), .Z(n8900) );
  AND U9195 ( .A(n8901), .B(n8900), .Z(n9069) );
  NANDN U9196 ( .A(n8903), .B(n8902), .Z(n8907) );
  NANDN U9197 ( .A(n8905), .B(n8904), .Z(n8906) );
  NAND U9198 ( .A(n8907), .B(n8906), .Z(n9070) );
  XNOR U9199 ( .A(n9069), .B(n9070), .Z(n9071) );
  NANDN U9200 ( .A(n8909), .B(n8908), .Z(n8913) );
  NANDN U9201 ( .A(n8911), .B(n8910), .Z(n8912) );
  NAND U9202 ( .A(n8913), .B(n8912), .Z(n9072) );
  XNOR U9203 ( .A(n9071), .B(n9072), .Z(n9015) );
  XNOR U9204 ( .A(n9016), .B(n9015), .Z(n9018) );
  NANDN U9205 ( .A(n8915), .B(n8914), .Z(n8919) );
  NANDN U9206 ( .A(n8917), .B(n8916), .Z(n8918) );
  AND U9207 ( .A(n8919), .B(n8918), .Z(n9017) );
  XOR U9208 ( .A(n9018), .B(n9017), .Z(n9132) );
  NANDN U9209 ( .A(n8921), .B(n8920), .Z(n8925) );
  NANDN U9210 ( .A(n8923), .B(n8922), .Z(n8924) );
  AND U9211 ( .A(n8925), .B(n8924), .Z(n9129) );
  NANDN U9212 ( .A(n8927), .B(n8926), .Z(n8931) );
  NANDN U9213 ( .A(n8929), .B(n8928), .Z(n8930) );
  AND U9214 ( .A(n8931), .B(n8930), .Z(n9012) );
  NANDN U9215 ( .A(n8933), .B(n8932), .Z(n8937) );
  OR U9216 ( .A(n8935), .B(n8934), .Z(n8936) );
  AND U9217 ( .A(n8937), .B(n8936), .Z(n9010) );
  NANDN U9218 ( .A(n8939), .B(n8938), .Z(n8943) );
  NANDN U9219 ( .A(n8941), .B(n8940), .Z(n8942) );
  AND U9220 ( .A(n8943), .B(n8942), .Z(n9076) );
  NANDN U9221 ( .A(n8945), .B(n8944), .Z(n8949) );
  NANDN U9222 ( .A(n8947), .B(n8946), .Z(n8948) );
  NAND U9223 ( .A(n8949), .B(n8948), .Z(n9075) );
  XNOR U9224 ( .A(n9076), .B(n9075), .Z(n9077) );
  NAND U9225 ( .A(b[0]), .B(a[75]), .Z(n8950) );
  XNOR U9226 ( .A(b[1]), .B(n8950), .Z(n8952) );
  NANDN U9227 ( .A(b[0]), .B(a[74]), .Z(n8951) );
  NAND U9228 ( .A(n8952), .B(n8951), .Z(n9024) );
  NANDN U9229 ( .A(n19394), .B(n8953), .Z(n8955) );
  XOR U9230 ( .A(b[29]), .B(a[47]), .Z(n9102) );
  NANDN U9231 ( .A(n19395), .B(n9102), .Z(n8954) );
  AND U9232 ( .A(n8955), .B(n8954), .Z(n9022) );
  AND U9233 ( .A(b[31]), .B(a[43]), .Z(n9021) );
  XNOR U9234 ( .A(n9022), .B(n9021), .Z(n9023) );
  XNOR U9235 ( .A(n9024), .B(n9023), .Z(n9063) );
  NANDN U9236 ( .A(n19005), .B(n8956), .Z(n8958) );
  XOR U9237 ( .A(b[23]), .B(a[53]), .Z(n9105) );
  NANDN U9238 ( .A(n19055), .B(n9105), .Z(n8957) );
  AND U9239 ( .A(n8958), .B(n8957), .Z(n9096) );
  NANDN U9240 ( .A(n17362), .B(n8959), .Z(n8961) );
  XOR U9241 ( .A(b[7]), .B(a[69]), .Z(n9108) );
  NANDN U9242 ( .A(n17522), .B(n9108), .Z(n8960) );
  AND U9243 ( .A(n8961), .B(n8960), .Z(n9094) );
  NANDN U9244 ( .A(n19116), .B(n8962), .Z(n8964) );
  XOR U9245 ( .A(b[25]), .B(a[51]), .Z(n9111) );
  NANDN U9246 ( .A(n19179), .B(n9111), .Z(n8963) );
  NAND U9247 ( .A(n8964), .B(n8963), .Z(n9093) );
  XNOR U9248 ( .A(n9094), .B(n9093), .Z(n9095) );
  XOR U9249 ( .A(n9096), .B(n9095), .Z(n9064) );
  XNOR U9250 ( .A(n9063), .B(n9064), .Z(n9065) );
  NANDN U9251 ( .A(n18113), .B(n8965), .Z(n8967) );
  XOR U9252 ( .A(b[13]), .B(a[63]), .Z(n9114) );
  NANDN U9253 ( .A(n18229), .B(n9114), .Z(n8966) );
  AND U9254 ( .A(n8967), .B(n8966), .Z(n9058) );
  NANDN U9255 ( .A(n17888), .B(n8968), .Z(n8970) );
  XOR U9256 ( .A(b[11]), .B(a[65]), .Z(n9117) );
  NANDN U9257 ( .A(n18025), .B(n9117), .Z(n8969) );
  NAND U9258 ( .A(n8970), .B(n8969), .Z(n9057) );
  XNOR U9259 ( .A(n9058), .B(n9057), .Z(n9059) );
  NANDN U9260 ( .A(n18487), .B(n8971), .Z(n8973) );
  XOR U9261 ( .A(b[15]), .B(a[61]), .Z(n9120) );
  NANDN U9262 ( .A(n18311), .B(n9120), .Z(n8972) );
  AND U9263 ( .A(n8973), .B(n8972), .Z(n9054) );
  NANDN U9264 ( .A(n18853), .B(n8974), .Z(n8976) );
  XOR U9265 ( .A(b[21]), .B(a[55]), .Z(n9123) );
  NANDN U9266 ( .A(n18926), .B(n9123), .Z(n8975) );
  AND U9267 ( .A(n8976), .B(n8975), .Z(n9052) );
  NANDN U9268 ( .A(n17613), .B(n8977), .Z(n8979) );
  XOR U9269 ( .A(b[9]), .B(a[67]), .Z(n9126) );
  NANDN U9270 ( .A(n17739), .B(n9126), .Z(n8978) );
  NAND U9271 ( .A(n8979), .B(n8978), .Z(n9051) );
  XNOR U9272 ( .A(n9052), .B(n9051), .Z(n9053) );
  XOR U9273 ( .A(n9054), .B(n9053), .Z(n9060) );
  XOR U9274 ( .A(n9059), .B(n9060), .Z(n9066) );
  XOR U9275 ( .A(n9065), .B(n9066), .Z(n9078) );
  XNOR U9276 ( .A(n9077), .B(n9078), .Z(n9009) );
  XNOR U9277 ( .A(n9010), .B(n9009), .Z(n9011) );
  XOR U9278 ( .A(n9012), .B(n9011), .Z(n9130) );
  XNOR U9279 ( .A(n9129), .B(n9130), .Z(n9131) );
  XNOR U9280 ( .A(n9132), .B(n9131), .Z(n9005) );
  XOR U9281 ( .A(n9006), .B(n9005), .Z(n8998) );
  NANDN U9282 ( .A(n8981), .B(n8980), .Z(n8985) );
  NANDN U9283 ( .A(n8983), .B(n8982), .Z(n8984) );
  AND U9284 ( .A(n8985), .B(n8984), .Z(n8997) );
  XOR U9285 ( .A(n8998), .B(n8997), .Z(n9000) );
  XNOR U9286 ( .A(n8999), .B(n9000), .Z(n8991) );
  XNOR U9287 ( .A(n8992), .B(n8991), .Z(n8993) );
  XNOR U9288 ( .A(n8994), .B(n8993), .Z(n9135) );
  XNOR U9289 ( .A(sreg[171]), .B(n9135), .Z(n9137) );
  NANDN U9290 ( .A(sreg[170]), .B(n8986), .Z(n8990) );
  NAND U9291 ( .A(n8988), .B(n8987), .Z(n8989) );
  NAND U9292 ( .A(n8990), .B(n8989), .Z(n9136) );
  XNOR U9293 ( .A(n9137), .B(n9136), .Z(c[171]) );
  NANDN U9294 ( .A(n8992), .B(n8991), .Z(n8996) );
  NANDN U9295 ( .A(n8994), .B(n8993), .Z(n8995) );
  AND U9296 ( .A(n8996), .B(n8995), .Z(n9143) );
  NANDN U9297 ( .A(n8998), .B(n8997), .Z(n9002) );
  NANDN U9298 ( .A(n9000), .B(n8999), .Z(n9001) );
  AND U9299 ( .A(n9002), .B(n9001), .Z(n9141) );
  NANDN U9300 ( .A(n9004), .B(n9003), .Z(n9008) );
  NAND U9301 ( .A(n9006), .B(n9005), .Z(n9007) );
  AND U9302 ( .A(n9008), .B(n9007), .Z(n9148) );
  NANDN U9303 ( .A(n9010), .B(n9009), .Z(n9014) );
  NANDN U9304 ( .A(n9012), .B(n9011), .Z(n9013) );
  AND U9305 ( .A(n9014), .B(n9013), .Z(n9153) );
  NANDN U9306 ( .A(n9016), .B(n9015), .Z(n9020) );
  NAND U9307 ( .A(n9018), .B(n9017), .Z(n9019) );
  AND U9308 ( .A(n9020), .B(n9019), .Z(n9152) );
  XNOR U9309 ( .A(n9153), .B(n9152), .Z(n9155) );
  NANDN U9310 ( .A(n9022), .B(n9021), .Z(n9026) );
  NANDN U9311 ( .A(n9024), .B(n9023), .Z(n9025) );
  AND U9312 ( .A(n9026), .B(n9025), .Z(n9232) );
  NANDN U9313 ( .A(n19237), .B(n9027), .Z(n9029) );
  XOR U9314 ( .A(b[27]), .B(a[50]), .Z(n9176) );
  NANDN U9315 ( .A(n19277), .B(n9176), .Z(n9028) );
  AND U9316 ( .A(n9029), .B(n9028), .Z(n9239) );
  NANDN U9317 ( .A(n17072), .B(n9030), .Z(n9032) );
  XOR U9318 ( .A(b[5]), .B(a[72]), .Z(n9179) );
  NANDN U9319 ( .A(n17223), .B(n9179), .Z(n9031) );
  AND U9320 ( .A(n9032), .B(n9031), .Z(n9237) );
  NANDN U9321 ( .A(n18673), .B(n9033), .Z(n9035) );
  XOR U9322 ( .A(b[19]), .B(a[58]), .Z(n9182) );
  NANDN U9323 ( .A(n18758), .B(n9182), .Z(n9034) );
  NAND U9324 ( .A(n9035), .B(n9034), .Z(n9236) );
  XNOR U9325 ( .A(n9237), .B(n9236), .Z(n9238) );
  XNOR U9326 ( .A(n9239), .B(n9238), .Z(n9230) );
  NANDN U9327 ( .A(n19425), .B(n9036), .Z(n9038) );
  XOR U9328 ( .A(b[31]), .B(a[46]), .Z(n9185) );
  NANDN U9329 ( .A(n19426), .B(n9185), .Z(n9037) );
  AND U9330 ( .A(n9038), .B(n9037), .Z(n9197) );
  NANDN U9331 ( .A(n17067), .B(n9039), .Z(n9041) );
  XOR U9332 ( .A(b[3]), .B(a[74]), .Z(n9188) );
  NANDN U9333 ( .A(n17068), .B(n9188), .Z(n9040) );
  AND U9334 ( .A(n9041), .B(n9040), .Z(n9195) );
  NANDN U9335 ( .A(n18514), .B(n9042), .Z(n9044) );
  XOR U9336 ( .A(b[17]), .B(a[60]), .Z(n9191) );
  NANDN U9337 ( .A(n18585), .B(n9191), .Z(n9043) );
  NAND U9338 ( .A(n9044), .B(n9043), .Z(n9194) );
  XNOR U9339 ( .A(n9195), .B(n9194), .Z(n9196) );
  XOR U9340 ( .A(n9197), .B(n9196), .Z(n9231) );
  XOR U9341 ( .A(n9230), .B(n9231), .Z(n9233) );
  XOR U9342 ( .A(n9232), .B(n9233), .Z(n9165) );
  NANDN U9343 ( .A(n9046), .B(n9045), .Z(n9050) );
  NANDN U9344 ( .A(n9048), .B(n9047), .Z(n9049) );
  AND U9345 ( .A(n9050), .B(n9049), .Z(n9218) );
  NANDN U9346 ( .A(n9052), .B(n9051), .Z(n9056) );
  NANDN U9347 ( .A(n9054), .B(n9053), .Z(n9055) );
  NAND U9348 ( .A(n9056), .B(n9055), .Z(n9219) );
  XNOR U9349 ( .A(n9218), .B(n9219), .Z(n9220) );
  NANDN U9350 ( .A(n9058), .B(n9057), .Z(n9062) );
  NANDN U9351 ( .A(n9060), .B(n9059), .Z(n9061) );
  NAND U9352 ( .A(n9062), .B(n9061), .Z(n9221) );
  XNOR U9353 ( .A(n9220), .B(n9221), .Z(n9164) );
  XNOR U9354 ( .A(n9165), .B(n9164), .Z(n9167) );
  NANDN U9355 ( .A(n9064), .B(n9063), .Z(n9068) );
  NANDN U9356 ( .A(n9066), .B(n9065), .Z(n9067) );
  AND U9357 ( .A(n9068), .B(n9067), .Z(n9166) );
  XOR U9358 ( .A(n9167), .B(n9166), .Z(n9281) );
  NANDN U9359 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U9360 ( .A(n9072), .B(n9071), .Z(n9073) );
  AND U9361 ( .A(n9074), .B(n9073), .Z(n9278) );
  NANDN U9362 ( .A(n9076), .B(n9075), .Z(n9080) );
  NANDN U9363 ( .A(n9078), .B(n9077), .Z(n9079) );
  AND U9364 ( .A(n9080), .B(n9079), .Z(n9161) );
  NANDN U9365 ( .A(n9082), .B(n9081), .Z(n9086) );
  OR U9366 ( .A(n9084), .B(n9083), .Z(n9085) );
  AND U9367 ( .A(n9086), .B(n9085), .Z(n9159) );
  NANDN U9368 ( .A(n9088), .B(n9087), .Z(n9092) );
  NANDN U9369 ( .A(n9090), .B(n9089), .Z(n9091) );
  AND U9370 ( .A(n9092), .B(n9091), .Z(n9225) );
  NANDN U9371 ( .A(n9094), .B(n9093), .Z(n9098) );
  NANDN U9372 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U9373 ( .A(n9098), .B(n9097), .Z(n9224) );
  XNOR U9374 ( .A(n9225), .B(n9224), .Z(n9226) );
  NAND U9375 ( .A(b[0]), .B(a[76]), .Z(n9099) );
  XNOR U9376 ( .A(b[1]), .B(n9099), .Z(n9101) );
  NANDN U9377 ( .A(b[0]), .B(a[75]), .Z(n9100) );
  NAND U9378 ( .A(n9101), .B(n9100), .Z(n9173) );
  NANDN U9379 ( .A(n19394), .B(n9102), .Z(n9104) );
  XOR U9380 ( .A(b[29]), .B(a[48]), .Z(n9248) );
  NANDN U9381 ( .A(n19395), .B(n9248), .Z(n9103) );
  AND U9382 ( .A(n9104), .B(n9103), .Z(n9171) );
  AND U9383 ( .A(b[31]), .B(a[44]), .Z(n9170) );
  XNOR U9384 ( .A(n9171), .B(n9170), .Z(n9172) );
  XNOR U9385 ( .A(n9173), .B(n9172), .Z(n9212) );
  NANDN U9386 ( .A(n19005), .B(n9105), .Z(n9107) );
  XOR U9387 ( .A(b[23]), .B(a[54]), .Z(n9254) );
  NANDN U9388 ( .A(n19055), .B(n9254), .Z(n9106) );
  AND U9389 ( .A(n9107), .B(n9106), .Z(n9245) );
  NANDN U9390 ( .A(n17362), .B(n9108), .Z(n9110) );
  XOR U9391 ( .A(b[7]), .B(a[70]), .Z(n9257) );
  NANDN U9392 ( .A(n17522), .B(n9257), .Z(n9109) );
  AND U9393 ( .A(n9110), .B(n9109), .Z(n9243) );
  NANDN U9394 ( .A(n19116), .B(n9111), .Z(n9113) );
  XOR U9395 ( .A(b[25]), .B(a[52]), .Z(n9260) );
  NANDN U9396 ( .A(n19179), .B(n9260), .Z(n9112) );
  NAND U9397 ( .A(n9113), .B(n9112), .Z(n9242) );
  XNOR U9398 ( .A(n9243), .B(n9242), .Z(n9244) );
  XOR U9399 ( .A(n9245), .B(n9244), .Z(n9213) );
  XNOR U9400 ( .A(n9212), .B(n9213), .Z(n9214) );
  NANDN U9401 ( .A(n18113), .B(n9114), .Z(n9116) );
  XOR U9402 ( .A(b[13]), .B(a[64]), .Z(n9263) );
  NANDN U9403 ( .A(n18229), .B(n9263), .Z(n9115) );
  AND U9404 ( .A(n9116), .B(n9115), .Z(n9207) );
  NANDN U9405 ( .A(n17888), .B(n9117), .Z(n9119) );
  XOR U9406 ( .A(b[11]), .B(a[66]), .Z(n9266) );
  NANDN U9407 ( .A(n18025), .B(n9266), .Z(n9118) );
  NAND U9408 ( .A(n9119), .B(n9118), .Z(n9206) );
  XNOR U9409 ( .A(n9207), .B(n9206), .Z(n9208) );
  NANDN U9410 ( .A(n18487), .B(n9120), .Z(n9122) );
  XOR U9411 ( .A(b[15]), .B(a[62]), .Z(n9269) );
  NANDN U9412 ( .A(n18311), .B(n9269), .Z(n9121) );
  AND U9413 ( .A(n9122), .B(n9121), .Z(n9203) );
  NANDN U9414 ( .A(n18853), .B(n9123), .Z(n9125) );
  XOR U9415 ( .A(b[21]), .B(a[56]), .Z(n9272) );
  NANDN U9416 ( .A(n18926), .B(n9272), .Z(n9124) );
  AND U9417 ( .A(n9125), .B(n9124), .Z(n9201) );
  NANDN U9418 ( .A(n17613), .B(n9126), .Z(n9128) );
  XOR U9419 ( .A(b[9]), .B(a[68]), .Z(n9275) );
  NANDN U9420 ( .A(n17739), .B(n9275), .Z(n9127) );
  NAND U9421 ( .A(n9128), .B(n9127), .Z(n9200) );
  XNOR U9422 ( .A(n9201), .B(n9200), .Z(n9202) );
  XOR U9423 ( .A(n9203), .B(n9202), .Z(n9209) );
  XOR U9424 ( .A(n9208), .B(n9209), .Z(n9215) );
  XOR U9425 ( .A(n9214), .B(n9215), .Z(n9227) );
  XNOR U9426 ( .A(n9226), .B(n9227), .Z(n9158) );
  XNOR U9427 ( .A(n9159), .B(n9158), .Z(n9160) );
  XOR U9428 ( .A(n9161), .B(n9160), .Z(n9279) );
  XNOR U9429 ( .A(n9278), .B(n9279), .Z(n9280) );
  XNOR U9430 ( .A(n9281), .B(n9280), .Z(n9154) );
  XOR U9431 ( .A(n9155), .B(n9154), .Z(n9147) );
  NANDN U9432 ( .A(n9130), .B(n9129), .Z(n9134) );
  NANDN U9433 ( .A(n9132), .B(n9131), .Z(n9133) );
  AND U9434 ( .A(n9134), .B(n9133), .Z(n9146) );
  XOR U9435 ( .A(n9147), .B(n9146), .Z(n9149) );
  XNOR U9436 ( .A(n9148), .B(n9149), .Z(n9140) );
  XNOR U9437 ( .A(n9141), .B(n9140), .Z(n9142) );
  XNOR U9438 ( .A(n9143), .B(n9142), .Z(n9284) );
  XNOR U9439 ( .A(sreg[172]), .B(n9284), .Z(n9286) );
  NANDN U9440 ( .A(sreg[171]), .B(n9135), .Z(n9139) );
  NAND U9441 ( .A(n9137), .B(n9136), .Z(n9138) );
  NAND U9442 ( .A(n9139), .B(n9138), .Z(n9285) );
  XNOR U9443 ( .A(n9286), .B(n9285), .Z(c[172]) );
  NANDN U9444 ( .A(n9141), .B(n9140), .Z(n9145) );
  NANDN U9445 ( .A(n9143), .B(n9142), .Z(n9144) );
  AND U9446 ( .A(n9145), .B(n9144), .Z(n9292) );
  NANDN U9447 ( .A(n9147), .B(n9146), .Z(n9151) );
  NANDN U9448 ( .A(n9149), .B(n9148), .Z(n9150) );
  AND U9449 ( .A(n9151), .B(n9150), .Z(n9290) );
  NANDN U9450 ( .A(n9153), .B(n9152), .Z(n9157) );
  NAND U9451 ( .A(n9155), .B(n9154), .Z(n9156) );
  AND U9452 ( .A(n9157), .B(n9156), .Z(n9297) );
  NANDN U9453 ( .A(n9159), .B(n9158), .Z(n9163) );
  NANDN U9454 ( .A(n9161), .B(n9160), .Z(n9162) );
  AND U9455 ( .A(n9163), .B(n9162), .Z(n9302) );
  NANDN U9456 ( .A(n9165), .B(n9164), .Z(n9169) );
  NAND U9457 ( .A(n9167), .B(n9166), .Z(n9168) );
  AND U9458 ( .A(n9169), .B(n9168), .Z(n9301) );
  XNOR U9459 ( .A(n9302), .B(n9301), .Z(n9304) );
  NANDN U9460 ( .A(n9171), .B(n9170), .Z(n9175) );
  NANDN U9461 ( .A(n9173), .B(n9172), .Z(n9174) );
  AND U9462 ( .A(n9175), .B(n9174), .Z(n9379) );
  NANDN U9463 ( .A(n19237), .B(n9176), .Z(n9178) );
  XOR U9464 ( .A(b[27]), .B(a[51]), .Z(n9325) );
  NANDN U9465 ( .A(n19277), .B(n9325), .Z(n9177) );
  AND U9466 ( .A(n9178), .B(n9177), .Z(n9386) );
  NANDN U9467 ( .A(n17072), .B(n9179), .Z(n9181) );
  XOR U9468 ( .A(b[5]), .B(a[73]), .Z(n9328) );
  NANDN U9469 ( .A(n17223), .B(n9328), .Z(n9180) );
  AND U9470 ( .A(n9181), .B(n9180), .Z(n9384) );
  NANDN U9471 ( .A(n18673), .B(n9182), .Z(n9184) );
  XOR U9472 ( .A(b[19]), .B(a[59]), .Z(n9331) );
  NANDN U9473 ( .A(n18758), .B(n9331), .Z(n9183) );
  NAND U9474 ( .A(n9184), .B(n9183), .Z(n9383) );
  XNOR U9475 ( .A(n9384), .B(n9383), .Z(n9385) );
  XNOR U9476 ( .A(n9386), .B(n9385), .Z(n9377) );
  NANDN U9477 ( .A(n19425), .B(n9185), .Z(n9187) );
  XOR U9478 ( .A(b[31]), .B(a[47]), .Z(n9334) );
  NANDN U9479 ( .A(n19426), .B(n9334), .Z(n9186) );
  AND U9480 ( .A(n9187), .B(n9186), .Z(n9346) );
  NANDN U9481 ( .A(n17067), .B(n9188), .Z(n9190) );
  XOR U9482 ( .A(b[3]), .B(a[75]), .Z(n9337) );
  NANDN U9483 ( .A(n17068), .B(n9337), .Z(n9189) );
  AND U9484 ( .A(n9190), .B(n9189), .Z(n9344) );
  NANDN U9485 ( .A(n18514), .B(n9191), .Z(n9193) );
  XOR U9486 ( .A(b[17]), .B(a[61]), .Z(n9340) );
  NANDN U9487 ( .A(n18585), .B(n9340), .Z(n9192) );
  NAND U9488 ( .A(n9193), .B(n9192), .Z(n9343) );
  XNOR U9489 ( .A(n9344), .B(n9343), .Z(n9345) );
  XOR U9490 ( .A(n9346), .B(n9345), .Z(n9378) );
  XOR U9491 ( .A(n9377), .B(n9378), .Z(n9380) );
  XOR U9492 ( .A(n9379), .B(n9380), .Z(n9314) );
  NANDN U9493 ( .A(n9195), .B(n9194), .Z(n9199) );
  NANDN U9494 ( .A(n9197), .B(n9196), .Z(n9198) );
  AND U9495 ( .A(n9199), .B(n9198), .Z(n9367) );
  NANDN U9496 ( .A(n9201), .B(n9200), .Z(n9205) );
  NANDN U9497 ( .A(n9203), .B(n9202), .Z(n9204) );
  NAND U9498 ( .A(n9205), .B(n9204), .Z(n9368) );
  XNOR U9499 ( .A(n9367), .B(n9368), .Z(n9369) );
  NANDN U9500 ( .A(n9207), .B(n9206), .Z(n9211) );
  NANDN U9501 ( .A(n9209), .B(n9208), .Z(n9210) );
  NAND U9502 ( .A(n9211), .B(n9210), .Z(n9370) );
  XNOR U9503 ( .A(n9369), .B(n9370), .Z(n9313) );
  XNOR U9504 ( .A(n9314), .B(n9313), .Z(n9316) );
  NANDN U9505 ( .A(n9213), .B(n9212), .Z(n9217) );
  NANDN U9506 ( .A(n9215), .B(n9214), .Z(n9216) );
  AND U9507 ( .A(n9217), .B(n9216), .Z(n9315) );
  XOR U9508 ( .A(n9316), .B(n9315), .Z(n9428) );
  NANDN U9509 ( .A(n9219), .B(n9218), .Z(n9223) );
  NANDN U9510 ( .A(n9221), .B(n9220), .Z(n9222) );
  AND U9511 ( .A(n9223), .B(n9222), .Z(n9425) );
  NANDN U9512 ( .A(n9225), .B(n9224), .Z(n9229) );
  NANDN U9513 ( .A(n9227), .B(n9226), .Z(n9228) );
  AND U9514 ( .A(n9229), .B(n9228), .Z(n9310) );
  NANDN U9515 ( .A(n9231), .B(n9230), .Z(n9235) );
  OR U9516 ( .A(n9233), .B(n9232), .Z(n9234) );
  AND U9517 ( .A(n9235), .B(n9234), .Z(n9308) );
  NANDN U9518 ( .A(n9237), .B(n9236), .Z(n9241) );
  NANDN U9519 ( .A(n9239), .B(n9238), .Z(n9240) );
  AND U9520 ( .A(n9241), .B(n9240), .Z(n9374) );
  NANDN U9521 ( .A(n9243), .B(n9242), .Z(n9247) );
  NANDN U9522 ( .A(n9245), .B(n9244), .Z(n9246) );
  NAND U9523 ( .A(n9247), .B(n9246), .Z(n9373) );
  XNOR U9524 ( .A(n9374), .B(n9373), .Z(n9376) );
  NANDN U9525 ( .A(n19394), .B(n9248), .Z(n9250) );
  XOR U9526 ( .A(b[29]), .B(a[49]), .Z(n9398) );
  NANDN U9527 ( .A(n19395), .B(n9398), .Z(n9249) );
  AND U9528 ( .A(n9250), .B(n9249), .Z(n9320) );
  AND U9529 ( .A(b[31]), .B(a[45]), .Z(n9319) );
  XNOR U9530 ( .A(n9320), .B(n9319), .Z(n9321) );
  NAND U9531 ( .A(b[0]), .B(a[77]), .Z(n9251) );
  XNOR U9532 ( .A(b[1]), .B(n9251), .Z(n9253) );
  NANDN U9533 ( .A(b[0]), .B(a[76]), .Z(n9252) );
  NAND U9534 ( .A(n9253), .B(n9252), .Z(n9322) );
  XNOR U9535 ( .A(n9321), .B(n9322), .Z(n9362) );
  NANDN U9536 ( .A(n19005), .B(n9254), .Z(n9256) );
  XOR U9537 ( .A(b[23]), .B(a[55]), .Z(n9401) );
  NANDN U9538 ( .A(n19055), .B(n9401), .Z(n9255) );
  AND U9539 ( .A(n9256), .B(n9255), .Z(n9391) );
  NANDN U9540 ( .A(n17362), .B(n9257), .Z(n9259) );
  XOR U9541 ( .A(b[7]), .B(a[71]), .Z(n9404) );
  NANDN U9542 ( .A(n17522), .B(n9404), .Z(n9258) );
  AND U9543 ( .A(n9259), .B(n9258), .Z(n9390) );
  NANDN U9544 ( .A(n19116), .B(n9260), .Z(n9262) );
  XOR U9545 ( .A(b[25]), .B(a[53]), .Z(n9407) );
  NANDN U9546 ( .A(n19179), .B(n9407), .Z(n9261) );
  NAND U9547 ( .A(n9262), .B(n9261), .Z(n9389) );
  XOR U9548 ( .A(n9390), .B(n9389), .Z(n9392) );
  XOR U9549 ( .A(n9391), .B(n9392), .Z(n9361) );
  XOR U9550 ( .A(n9362), .B(n9361), .Z(n9364) );
  NANDN U9551 ( .A(n18113), .B(n9263), .Z(n9265) );
  XOR U9552 ( .A(b[13]), .B(a[65]), .Z(n9410) );
  NANDN U9553 ( .A(n18229), .B(n9410), .Z(n9264) );
  AND U9554 ( .A(n9265), .B(n9264), .Z(n9356) );
  NANDN U9555 ( .A(n17888), .B(n9266), .Z(n9268) );
  XOR U9556 ( .A(b[11]), .B(a[67]), .Z(n9413) );
  NANDN U9557 ( .A(n18025), .B(n9413), .Z(n9267) );
  NAND U9558 ( .A(n9268), .B(n9267), .Z(n9355) );
  XNOR U9559 ( .A(n9356), .B(n9355), .Z(n9358) );
  NANDN U9560 ( .A(n18487), .B(n9269), .Z(n9271) );
  XOR U9561 ( .A(b[15]), .B(a[63]), .Z(n9416) );
  NANDN U9562 ( .A(n18311), .B(n9416), .Z(n9270) );
  AND U9563 ( .A(n9271), .B(n9270), .Z(n9352) );
  NANDN U9564 ( .A(n18853), .B(n9272), .Z(n9274) );
  XOR U9565 ( .A(b[21]), .B(a[57]), .Z(n9419) );
  NANDN U9566 ( .A(n18926), .B(n9419), .Z(n9273) );
  AND U9567 ( .A(n9274), .B(n9273), .Z(n9350) );
  NANDN U9568 ( .A(n17613), .B(n9275), .Z(n9277) );
  XOR U9569 ( .A(b[9]), .B(a[69]), .Z(n9422) );
  NANDN U9570 ( .A(n17739), .B(n9422), .Z(n9276) );
  NAND U9571 ( .A(n9277), .B(n9276), .Z(n9349) );
  XNOR U9572 ( .A(n9350), .B(n9349), .Z(n9351) );
  XNOR U9573 ( .A(n9352), .B(n9351), .Z(n9357) );
  XOR U9574 ( .A(n9358), .B(n9357), .Z(n9363) );
  XOR U9575 ( .A(n9364), .B(n9363), .Z(n9375) );
  XOR U9576 ( .A(n9376), .B(n9375), .Z(n9307) );
  XNOR U9577 ( .A(n9308), .B(n9307), .Z(n9309) );
  XOR U9578 ( .A(n9310), .B(n9309), .Z(n9426) );
  XNOR U9579 ( .A(n9425), .B(n9426), .Z(n9427) );
  XNOR U9580 ( .A(n9428), .B(n9427), .Z(n9303) );
  XOR U9581 ( .A(n9304), .B(n9303), .Z(n9296) );
  NANDN U9582 ( .A(n9279), .B(n9278), .Z(n9283) );
  NANDN U9583 ( .A(n9281), .B(n9280), .Z(n9282) );
  AND U9584 ( .A(n9283), .B(n9282), .Z(n9295) );
  XOR U9585 ( .A(n9296), .B(n9295), .Z(n9298) );
  XNOR U9586 ( .A(n9297), .B(n9298), .Z(n9289) );
  XNOR U9587 ( .A(n9290), .B(n9289), .Z(n9291) );
  XNOR U9588 ( .A(n9292), .B(n9291), .Z(n9431) );
  XNOR U9589 ( .A(sreg[173]), .B(n9431), .Z(n9433) );
  NANDN U9590 ( .A(sreg[172]), .B(n9284), .Z(n9288) );
  NAND U9591 ( .A(n9286), .B(n9285), .Z(n9287) );
  NAND U9592 ( .A(n9288), .B(n9287), .Z(n9432) );
  XNOR U9593 ( .A(n9433), .B(n9432), .Z(c[173]) );
  NANDN U9594 ( .A(n9290), .B(n9289), .Z(n9294) );
  NANDN U9595 ( .A(n9292), .B(n9291), .Z(n9293) );
  AND U9596 ( .A(n9294), .B(n9293), .Z(n9438) );
  NANDN U9597 ( .A(n9296), .B(n9295), .Z(n9300) );
  NANDN U9598 ( .A(n9298), .B(n9297), .Z(n9299) );
  AND U9599 ( .A(n9300), .B(n9299), .Z(n9437) );
  NANDN U9600 ( .A(n9302), .B(n9301), .Z(n9306) );
  NAND U9601 ( .A(n9304), .B(n9303), .Z(n9305) );
  AND U9602 ( .A(n9306), .B(n9305), .Z(n9444) );
  NANDN U9603 ( .A(n9308), .B(n9307), .Z(n9312) );
  NANDN U9604 ( .A(n9310), .B(n9309), .Z(n9311) );
  AND U9605 ( .A(n9312), .B(n9311), .Z(n9573) );
  NANDN U9606 ( .A(n9314), .B(n9313), .Z(n9318) );
  NAND U9607 ( .A(n9316), .B(n9315), .Z(n9317) );
  AND U9608 ( .A(n9318), .B(n9317), .Z(n9572) );
  XNOR U9609 ( .A(n9573), .B(n9572), .Z(n9575) );
  NANDN U9610 ( .A(n9320), .B(n9319), .Z(n9324) );
  NANDN U9611 ( .A(n9322), .B(n9321), .Z(n9323) );
  AND U9612 ( .A(n9324), .B(n9323), .Z(n9508) );
  NANDN U9613 ( .A(n19237), .B(n9325), .Z(n9327) );
  XOR U9614 ( .A(b[27]), .B(a[52]), .Z(n9454) );
  NANDN U9615 ( .A(n19277), .B(n9454), .Z(n9326) );
  AND U9616 ( .A(n9327), .B(n9326), .Z(n9515) );
  NANDN U9617 ( .A(n17072), .B(n9328), .Z(n9330) );
  XOR U9618 ( .A(b[5]), .B(a[74]), .Z(n9457) );
  NANDN U9619 ( .A(n17223), .B(n9457), .Z(n9329) );
  AND U9620 ( .A(n9330), .B(n9329), .Z(n9513) );
  NANDN U9621 ( .A(n18673), .B(n9331), .Z(n9333) );
  XOR U9622 ( .A(b[19]), .B(a[60]), .Z(n9460) );
  NANDN U9623 ( .A(n18758), .B(n9460), .Z(n9332) );
  NAND U9624 ( .A(n9333), .B(n9332), .Z(n9512) );
  XNOR U9625 ( .A(n9513), .B(n9512), .Z(n9514) );
  XNOR U9626 ( .A(n9515), .B(n9514), .Z(n9506) );
  NANDN U9627 ( .A(n19425), .B(n9334), .Z(n9336) );
  XOR U9628 ( .A(b[31]), .B(a[48]), .Z(n9463) );
  NANDN U9629 ( .A(n19426), .B(n9463), .Z(n9335) );
  AND U9630 ( .A(n9336), .B(n9335), .Z(n9475) );
  NANDN U9631 ( .A(n17067), .B(n9337), .Z(n9339) );
  XOR U9632 ( .A(b[3]), .B(a[76]), .Z(n9466) );
  NANDN U9633 ( .A(n17068), .B(n9466), .Z(n9338) );
  AND U9634 ( .A(n9339), .B(n9338), .Z(n9473) );
  NANDN U9635 ( .A(n18514), .B(n9340), .Z(n9342) );
  XOR U9636 ( .A(b[17]), .B(a[62]), .Z(n9469) );
  NANDN U9637 ( .A(n18585), .B(n9469), .Z(n9341) );
  NAND U9638 ( .A(n9342), .B(n9341), .Z(n9472) );
  XNOR U9639 ( .A(n9473), .B(n9472), .Z(n9474) );
  XOR U9640 ( .A(n9475), .B(n9474), .Z(n9507) );
  XOR U9641 ( .A(n9506), .B(n9507), .Z(n9509) );
  XOR U9642 ( .A(n9508), .B(n9509), .Z(n9555) );
  NANDN U9643 ( .A(n9344), .B(n9343), .Z(n9348) );
  NANDN U9644 ( .A(n9346), .B(n9345), .Z(n9347) );
  AND U9645 ( .A(n9348), .B(n9347), .Z(n9496) );
  NANDN U9646 ( .A(n9350), .B(n9349), .Z(n9354) );
  NANDN U9647 ( .A(n9352), .B(n9351), .Z(n9353) );
  NAND U9648 ( .A(n9354), .B(n9353), .Z(n9497) );
  XNOR U9649 ( .A(n9496), .B(n9497), .Z(n9498) );
  NANDN U9650 ( .A(n9356), .B(n9355), .Z(n9360) );
  NAND U9651 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U9652 ( .A(n9360), .B(n9359), .Z(n9499) );
  XNOR U9653 ( .A(n9498), .B(n9499), .Z(n9554) );
  XNOR U9654 ( .A(n9555), .B(n9554), .Z(n9557) );
  NAND U9655 ( .A(n9362), .B(n9361), .Z(n9366) );
  NAND U9656 ( .A(n9364), .B(n9363), .Z(n9365) );
  AND U9657 ( .A(n9366), .B(n9365), .Z(n9556) );
  XOR U9658 ( .A(n9557), .B(n9556), .Z(n9569) );
  NANDN U9659 ( .A(n9368), .B(n9367), .Z(n9372) );
  NANDN U9660 ( .A(n9370), .B(n9369), .Z(n9371) );
  AND U9661 ( .A(n9372), .B(n9371), .Z(n9566) );
  NANDN U9662 ( .A(n9378), .B(n9377), .Z(n9382) );
  OR U9663 ( .A(n9380), .B(n9379), .Z(n9381) );
  AND U9664 ( .A(n9382), .B(n9381), .Z(n9561) );
  NANDN U9665 ( .A(n9384), .B(n9383), .Z(n9388) );
  NANDN U9666 ( .A(n9386), .B(n9385), .Z(n9387) );
  AND U9667 ( .A(n9388), .B(n9387), .Z(n9503) );
  NANDN U9668 ( .A(n9390), .B(n9389), .Z(n9394) );
  OR U9669 ( .A(n9392), .B(n9391), .Z(n9393) );
  NAND U9670 ( .A(n9394), .B(n9393), .Z(n9502) );
  XNOR U9671 ( .A(n9503), .B(n9502), .Z(n9505) );
  NAND U9672 ( .A(b[0]), .B(a[78]), .Z(n9395) );
  XNOR U9673 ( .A(b[1]), .B(n9395), .Z(n9397) );
  NANDN U9674 ( .A(b[0]), .B(a[77]), .Z(n9396) );
  NAND U9675 ( .A(n9397), .B(n9396), .Z(n9451) );
  NANDN U9676 ( .A(n19394), .B(n9398), .Z(n9400) );
  XOR U9677 ( .A(b[29]), .B(a[50]), .Z(n9527) );
  NANDN U9678 ( .A(n19395), .B(n9527), .Z(n9399) );
  AND U9679 ( .A(n9400), .B(n9399), .Z(n9449) );
  AND U9680 ( .A(b[31]), .B(a[46]), .Z(n9448) );
  XNOR U9681 ( .A(n9449), .B(n9448), .Z(n9450) );
  XNOR U9682 ( .A(n9451), .B(n9450), .Z(n9491) );
  NANDN U9683 ( .A(n19005), .B(n9401), .Z(n9403) );
  XOR U9684 ( .A(b[23]), .B(a[56]), .Z(n9530) );
  NANDN U9685 ( .A(n19055), .B(n9530), .Z(n9402) );
  AND U9686 ( .A(n9403), .B(n9402), .Z(n9520) );
  NANDN U9687 ( .A(n17362), .B(n9404), .Z(n9406) );
  XOR U9688 ( .A(b[7]), .B(a[72]), .Z(n9533) );
  NANDN U9689 ( .A(n17522), .B(n9533), .Z(n9405) );
  AND U9690 ( .A(n9406), .B(n9405), .Z(n9519) );
  NANDN U9691 ( .A(n19116), .B(n9407), .Z(n9409) );
  XOR U9692 ( .A(b[25]), .B(a[54]), .Z(n9536) );
  NANDN U9693 ( .A(n19179), .B(n9536), .Z(n9408) );
  NAND U9694 ( .A(n9409), .B(n9408), .Z(n9518) );
  XOR U9695 ( .A(n9519), .B(n9518), .Z(n9521) );
  XOR U9696 ( .A(n9520), .B(n9521), .Z(n9490) );
  XOR U9697 ( .A(n9491), .B(n9490), .Z(n9493) );
  NANDN U9698 ( .A(n18113), .B(n9410), .Z(n9412) );
  XOR U9699 ( .A(b[13]), .B(a[66]), .Z(n9539) );
  NANDN U9700 ( .A(n18229), .B(n9539), .Z(n9411) );
  AND U9701 ( .A(n9412), .B(n9411), .Z(n9485) );
  NANDN U9702 ( .A(n17888), .B(n9413), .Z(n9415) );
  XOR U9703 ( .A(b[11]), .B(a[68]), .Z(n9542) );
  NANDN U9704 ( .A(n18025), .B(n9542), .Z(n9414) );
  NAND U9705 ( .A(n9415), .B(n9414), .Z(n9484) );
  XNOR U9706 ( .A(n9485), .B(n9484), .Z(n9487) );
  NANDN U9707 ( .A(n18487), .B(n9416), .Z(n9418) );
  XOR U9708 ( .A(b[15]), .B(a[64]), .Z(n9545) );
  NANDN U9709 ( .A(n18311), .B(n9545), .Z(n9417) );
  AND U9710 ( .A(n9418), .B(n9417), .Z(n9481) );
  NANDN U9711 ( .A(n18853), .B(n9419), .Z(n9421) );
  XOR U9712 ( .A(b[21]), .B(a[58]), .Z(n9548) );
  NANDN U9713 ( .A(n18926), .B(n9548), .Z(n9420) );
  AND U9714 ( .A(n9421), .B(n9420), .Z(n9479) );
  NANDN U9715 ( .A(n17613), .B(n9422), .Z(n9424) );
  XOR U9716 ( .A(b[9]), .B(a[70]), .Z(n9551) );
  NANDN U9717 ( .A(n17739), .B(n9551), .Z(n9423) );
  NAND U9718 ( .A(n9424), .B(n9423), .Z(n9478) );
  XNOR U9719 ( .A(n9479), .B(n9478), .Z(n9480) );
  XNOR U9720 ( .A(n9481), .B(n9480), .Z(n9486) );
  XOR U9721 ( .A(n9487), .B(n9486), .Z(n9492) );
  XOR U9722 ( .A(n9493), .B(n9492), .Z(n9504) );
  XOR U9723 ( .A(n9505), .B(n9504), .Z(n9560) );
  XNOR U9724 ( .A(n9561), .B(n9560), .Z(n9562) );
  XOR U9725 ( .A(n9563), .B(n9562), .Z(n9567) );
  XNOR U9726 ( .A(n9566), .B(n9567), .Z(n9568) );
  XNOR U9727 ( .A(n9569), .B(n9568), .Z(n9574) );
  XOR U9728 ( .A(n9575), .B(n9574), .Z(n9443) );
  NANDN U9729 ( .A(n9426), .B(n9425), .Z(n9430) );
  NANDN U9730 ( .A(n9428), .B(n9427), .Z(n9429) );
  AND U9731 ( .A(n9430), .B(n9429), .Z(n9442) );
  XOR U9732 ( .A(n9443), .B(n9442), .Z(n9445) );
  XNOR U9733 ( .A(n9444), .B(n9445), .Z(n9436) );
  XOR U9734 ( .A(n9437), .B(n9436), .Z(n9439) );
  XOR U9735 ( .A(n9438), .B(n9439), .Z(n9578) );
  XNOR U9736 ( .A(n9578), .B(sreg[174]), .Z(n9580) );
  NANDN U9737 ( .A(sreg[173]), .B(n9431), .Z(n9435) );
  NAND U9738 ( .A(n9433), .B(n9432), .Z(n9434) );
  AND U9739 ( .A(n9435), .B(n9434), .Z(n9579) );
  XOR U9740 ( .A(n9580), .B(n9579), .Z(c[174]) );
  NANDN U9741 ( .A(n9437), .B(n9436), .Z(n9441) );
  OR U9742 ( .A(n9439), .B(n9438), .Z(n9440) );
  AND U9743 ( .A(n9441), .B(n9440), .Z(n9586) );
  NANDN U9744 ( .A(n9443), .B(n9442), .Z(n9447) );
  NANDN U9745 ( .A(n9445), .B(n9444), .Z(n9446) );
  AND U9746 ( .A(n9447), .B(n9446), .Z(n9584) );
  NANDN U9747 ( .A(n9449), .B(n9448), .Z(n9453) );
  NANDN U9748 ( .A(n9451), .B(n9450), .Z(n9452) );
  AND U9749 ( .A(n9453), .B(n9452), .Z(n9661) );
  NANDN U9750 ( .A(n19237), .B(n9454), .Z(n9456) );
  XOR U9751 ( .A(b[27]), .B(a[53]), .Z(n9607) );
  NANDN U9752 ( .A(n19277), .B(n9607), .Z(n9455) );
  AND U9753 ( .A(n9456), .B(n9455), .Z(n9668) );
  NANDN U9754 ( .A(n17072), .B(n9457), .Z(n9459) );
  XOR U9755 ( .A(b[5]), .B(a[75]), .Z(n9610) );
  NANDN U9756 ( .A(n17223), .B(n9610), .Z(n9458) );
  AND U9757 ( .A(n9459), .B(n9458), .Z(n9666) );
  NANDN U9758 ( .A(n18673), .B(n9460), .Z(n9462) );
  XOR U9759 ( .A(b[19]), .B(a[61]), .Z(n9613) );
  NANDN U9760 ( .A(n18758), .B(n9613), .Z(n9461) );
  NAND U9761 ( .A(n9462), .B(n9461), .Z(n9665) );
  XNOR U9762 ( .A(n9666), .B(n9665), .Z(n9667) );
  XNOR U9763 ( .A(n9668), .B(n9667), .Z(n9659) );
  NANDN U9764 ( .A(n19425), .B(n9463), .Z(n9465) );
  XOR U9765 ( .A(b[31]), .B(a[49]), .Z(n9616) );
  NANDN U9766 ( .A(n19426), .B(n9616), .Z(n9464) );
  AND U9767 ( .A(n9465), .B(n9464), .Z(n9628) );
  NANDN U9768 ( .A(n17067), .B(n9466), .Z(n9468) );
  XOR U9769 ( .A(b[3]), .B(a[77]), .Z(n9619) );
  NANDN U9770 ( .A(n17068), .B(n9619), .Z(n9467) );
  AND U9771 ( .A(n9468), .B(n9467), .Z(n9626) );
  NANDN U9772 ( .A(n18514), .B(n9469), .Z(n9471) );
  XOR U9773 ( .A(b[17]), .B(a[63]), .Z(n9622) );
  NANDN U9774 ( .A(n18585), .B(n9622), .Z(n9470) );
  NAND U9775 ( .A(n9471), .B(n9470), .Z(n9625) );
  XNOR U9776 ( .A(n9626), .B(n9625), .Z(n9627) );
  XOR U9777 ( .A(n9628), .B(n9627), .Z(n9660) );
  XOR U9778 ( .A(n9659), .B(n9660), .Z(n9662) );
  XOR U9779 ( .A(n9661), .B(n9662), .Z(n9708) );
  NANDN U9780 ( .A(n9473), .B(n9472), .Z(n9477) );
  NANDN U9781 ( .A(n9475), .B(n9474), .Z(n9476) );
  AND U9782 ( .A(n9477), .B(n9476), .Z(n9649) );
  NANDN U9783 ( .A(n9479), .B(n9478), .Z(n9483) );
  NANDN U9784 ( .A(n9481), .B(n9480), .Z(n9482) );
  NAND U9785 ( .A(n9483), .B(n9482), .Z(n9650) );
  XNOR U9786 ( .A(n9649), .B(n9650), .Z(n9651) );
  NANDN U9787 ( .A(n9485), .B(n9484), .Z(n9489) );
  NAND U9788 ( .A(n9487), .B(n9486), .Z(n9488) );
  NAND U9789 ( .A(n9489), .B(n9488), .Z(n9652) );
  XNOR U9790 ( .A(n9651), .B(n9652), .Z(n9707) );
  XNOR U9791 ( .A(n9708), .B(n9707), .Z(n9710) );
  NAND U9792 ( .A(n9491), .B(n9490), .Z(n9495) );
  NAND U9793 ( .A(n9493), .B(n9492), .Z(n9494) );
  AND U9794 ( .A(n9495), .B(n9494), .Z(n9709) );
  XOR U9795 ( .A(n9710), .B(n9709), .Z(n9721) );
  NANDN U9796 ( .A(n9497), .B(n9496), .Z(n9501) );
  NANDN U9797 ( .A(n9499), .B(n9498), .Z(n9500) );
  AND U9798 ( .A(n9501), .B(n9500), .Z(n9719) );
  NANDN U9799 ( .A(n9507), .B(n9506), .Z(n9511) );
  OR U9800 ( .A(n9509), .B(n9508), .Z(n9510) );
  AND U9801 ( .A(n9511), .B(n9510), .Z(n9714) );
  NANDN U9802 ( .A(n9513), .B(n9512), .Z(n9517) );
  NANDN U9803 ( .A(n9515), .B(n9514), .Z(n9516) );
  AND U9804 ( .A(n9517), .B(n9516), .Z(n9656) );
  NANDN U9805 ( .A(n9519), .B(n9518), .Z(n9523) );
  OR U9806 ( .A(n9521), .B(n9520), .Z(n9522) );
  NAND U9807 ( .A(n9523), .B(n9522), .Z(n9655) );
  XNOR U9808 ( .A(n9656), .B(n9655), .Z(n9658) );
  NAND U9809 ( .A(b[0]), .B(a[79]), .Z(n9524) );
  XNOR U9810 ( .A(b[1]), .B(n9524), .Z(n9526) );
  NANDN U9811 ( .A(b[0]), .B(a[78]), .Z(n9525) );
  NAND U9812 ( .A(n9526), .B(n9525), .Z(n9604) );
  NANDN U9813 ( .A(n19394), .B(n9527), .Z(n9529) );
  XOR U9814 ( .A(b[29]), .B(a[51]), .Z(n9680) );
  NANDN U9815 ( .A(n19395), .B(n9680), .Z(n9528) );
  AND U9816 ( .A(n9529), .B(n9528), .Z(n9602) );
  AND U9817 ( .A(b[31]), .B(a[47]), .Z(n9601) );
  XNOR U9818 ( .A(n9602), .B(n9601), .Z(n9603) );
  XNOR U9819 ( .A(n9604), .B(n9603), .Z(n9644) );
  NANDN U9820 ( .A(n19005), .B(n9530), .Z(n9532) );
  XOR U9821 ( .A(b[23]), .B(a[57]), .Z(n9683) );
  NANDN U9822 ( .A(n19055), .B(n9683), .Z(n9531) );
  AND U9823 ( .A(n9532), .B(n9531), .Z(n9673) );
  NANDN U9824 ( .A(n17362), .B(n9533), .Z(n9535) );
  XOR U9825 ( .A(b[7]), .B(a[73]), .Z(n9686) );
  NANDN U9826 ( .A(n17522), .B(n9686), .Z(n9534) );
  AND U9827 ( .A(n9535), .B(n9534), .Z(n9672) );
  NANDN U9828 ( .A(n19116), .B(n9536), .Z(n9538) );
  XOR U9829 ( .A(b[25]), .B(a[55]), .Z(n9689) );
  NANDN U9830 ( .A(n19179), .B(n9689), .Z(n9537) );
  NAND U9831 ( .A(n9538), .B(n9537), .Z(n9671) );
  XOR U9832 ( .A(n9672), .B(n9671), .Z(n9674) );
  XOR U9833 ( .A(n9673), .B(n9674), .Z(n9643) );
  XOR U9834 ( .A(n9644), .B(n9643), .Z(n9646) );
  NANDN U9835 ( .A(n18113), .B(n9539), .Z(n9541) );
  XOR U9836 ( .A(b[13]), .B(a[67]), .Z(n9692) );
  NANDN U9837 ( .A(n18229), .B(n9692), .Z(n9540) );
  AND U9838 ( .A(n9541), .B(n9540), .Z(n9638) );
  NANDN U9839 ( .A(n17888), .B(n9542), .Z(n9544) );
  XOR U9840 ( .A(b[11]), .B(a[69]), .Z(n9695) );
  NANDN U9841 ( .A(n18025), .B(n9695), .Z(n9543) );
  NAND U9842 ( .A(n9544), .B(n9543), .Z(n9637) );
  XNOR U9843 ( .A(n9638), .B(n9637), .Z(n9640) );
  NANDN U9844 ( .A(n18487), .B(n9545), .Z(n9547) );
  XOR U9845 ( .A(b[15]), .B(a[65]), .Z(n9698) );
  NANDN U9846 ( .A(n18311), .B(n9698), .Z(n9546) );
  AND U9847 ( .A(n9547), .B(n9546), .Z(n9634) );
  NANDN U9848 ( .A(n18853), .B(n9548), .Z(n9550) );
  XOR U9849 ( .A(b[21]), .B(a[59]), .Z(n9701) );
  NANDN U9850 ( .A(n18926), .B(n9701), .Z(n9549) );
  AND U9851 ( .A(n9550), .B(n9549), .Z(n9632) );
  NANDN U9852 ( .A(n17613), .B(n9551), .Z(n9553) );
  XOR U9853 ( .A(b[9]), .B(a[71]), .Z(n9704) );
  NANDN U9854 ( .A(n17739), .B(n9704), .Z(n9552) );
  NAND U9855 ( .A(n9553), .B(n9552), .Z(n9631) );
  XNOR U9856 ( .A(n9632), .B(n9631), .Z(n9633) );
  XNOR U9857 ( .A(n9634), .B(n9633), .Z(n9639) );
  XOR U9858 ( .A(n9640), .B(n9639), .Z(n9645) );
  XOR U9859 ( .A(n9646), .B(n9645), .Z(n9657) );
  XOR U9860 ( .A(n9658), .B(n9657), .Z(n9713) );
  XNOR U9861 ( .A(n9714), .B(n9713), .Z(n9715) );
  XOR U9862 ( .A(n9716), .B(n9715), .Z(n9720) );
  XOR U9863 ( .A(n9719), .B(n9720), .Z(n9722) );
  XOR U9864 ( .A(n9721), .B(n9722), .Z(n9598) );
  NANDN U9865 ( .A(n9555), .B(n9554), .Z(n9559) );
  NAND U9866 ( .A(n9557), .B(n9556), .Z(n9558) );
  AND U9867 ( .A(n9559), .B(n9558), .Z(n9596) );
  NANDN U9868 ( .A(n9561), .B(n9560), .Z(n9565) );
  NANDN U9869 ( .A(n9563), .B(n9562), .Z(n9564) );
  AND U9870 ( .A(n9565), .B(n9564), .Z(n9595) );
  XNOR U9871 ( .A(n9596), .B(n9595), .Z(n9597) );
  XNOR U9872 ( .A(n9598), .B(n9597), .Z(n9589) );
  NANDN U9873 ( .A(n9567), .B(n9566), .Z(n9571) );
  NANDN U9874 ( .A(n9569), .B(n9568), .Z(n9570) );
  NAND U9875 ( .A(n9571), .B(n9570), .Z(n9590) );
  XNOR U9876 ( .A(n9589), .B(n9590), .Z(n9591) );
  NANDN U9877 ( .A(n9573), .B(n9572), .Z(n9577) );
  NAND U9878 ( .A(n9575), .B(n9574), .Z(n9576) );
  NAND U9879 ( .A(n9577), .B(n9576), .Z(n9592) );
  XNOR U9880 ( .A(n9591), .B(n9592), .Z(n9583) );
  XNOR U9881 ( .A(n9584), .B(n9583), .Z(n9585) );
  XNOR U9882 ( .A(n9586), .B(n9585), .Z(n9725) );
  XNOR U9883 ( .A(sreg[175]), .B(n9725), .Z(n9727) );
  NANDN U9884 ( .A(n9578), .B(sreg[174]), .Z(n9582) );
  NAND U9885 ( .A(n9580), .B(n9579), .Z(n9581) );
  AND U9886 ( .A(n9582), .B(n9581), .Z(n9726) );
  XNOR U9887 ( .A(n9727), .B(n9726), .Z(c[175]) );
  NANDN U9888 ( .A(n9584), .B(n9583), .Z(n9588) );
  NANDN U9889 ( .A(n9586), .B(n9585), .Z(n9587) );
  AND U9890 ( .A(n9588), .B(n9587), .Z(n9733) );
  NANDN U9891 ( .A(n9590), .B(n9589), .Z(n9594) );
  NANDN U9892 ( .A(n9592), .B(n9591), .Z(n9593) );
  AND U9893 ( .A(n9594), .B(n9593), .Z(n9731) );
  NANDN U9894 ( .A(n9596), .B(n9595), .Z(n9600) );
  NANDN U9895 ( .A(n9598), .B(n9597), .Z(n9599) );
  AND U9896 ( .A(n9600), .B(n9599), .Z(n9739) );
  NANDN U9897 ( .A(n9602), .B(n9601), .Z(n9606) );
  NANDN U9898 ( .A(n9604), .B(n9603), .Z(n9605) );
  AND U9899 ( .A(n9606), .B(n9605), .Z(n9810) );
  NANDN U9900 ( .A(n19237), .B(n9607), .Z(n9609) );
  XOR U9901 ( .A(b[27]), .B(a[54]), .Z(n9754) );
  NANDN U9902 ( .A(n19277), .B(n9754), .Z(n9608) );
  AND U9903 ( .A(n9609), .B(n9608), .Z(n9817) );
  NANDN U9904 ( .A(n17072), .B(n9610), .Z(n9612) );
  XOR U9905 ( .A(b[5]), .B(a[76]), .Z(n9757) );
  NANDN U9906 ( .A(n17223), .B(n9757), .Z(n9611) );
  AND U9907 ( .A(n9612), .B(n9611), .Z(n9815) );
  NANDN U9908 ( .A(n18673), .B(n9613), .Z(n9615) );
  XOR U9909 ( .A(b[19]), .B(a[62]), .Z(n9760) );
  NANDN U9910 ( .A(n18758), .B(n9760), .Z(n9614) );
  NAND U9911 ( .A(n9615), .B(n9614), .Z(n9814) );
  XNOR U9912 ( .A(n9815), .B(n9814), .Z(n9816) );
  XNOR U9913 ( .A(n9817), .B(n9816), .Z(n9808) );
  NANDN U9914 ( .A(n19425), .B(n9616), .Z(n9618) );
  XOR U9915 ( .A(b[31]), .B(a[50]), .Z(n9763) );
  NANDN U9916 ( .A(n19426), .B(n9763), .Z(n9617) );
  AND U9917 ( .A(n9618), .B(n9617), .Z(n9775) );
  NANDN U9918 ( .A(n17067), .B(n9619), .Z(n9621) );
  XOR U9919 ( .A(b[3]), .B(a[78]), .Z(n9766) );
  NANDN U9920 ( .A(n17068), .B(n9766), .Z(n9620) );
  AND U9921 ( .A(n9621), .B(n9620), .Z(n9773) );
  NANDN U9922 ( .A(n18514), .B(n9622), .Z(n9624) );
  XOR U9923 ( .A(b[17]), .B(a[64]), .Z(n9769) );
  NANDN U9924 ( .A(n18585), .B(n9769), .Z(n9623) );
  NAND U9925 ( .A(n9624), .B(n9623), .Z(n9772) );
  XNOR U9926 ( .A(n9773), .B(n9772), .Z(n9774) );
  XOR U9927 ( .A(n9775), .B(n9774), .Z(n9809) );
  XOR U9928 ( .A(n9808), .B(n9809), .Z(n9811) );
  XOR U9929 ( .A(n9810), .B(n9811), .Z(n9857) );
  NANDN U9930 ( .A(n9626), .B(n9625), .Z(n9630) );
  NANDN U9931 ( .A(n9628), .B(n9627), .Z(n9629) );
  AND U9932 ( .A(n9630), .B(n9629), .Z(n9796) );
  NANDN U9933 ( .A(n9632), .B(n9631), .Z(n9636) );
  NANDN U9934 ( .A(n9634), .B(n9633), .Z(n9635) );
  NAND U9935 ( .A(n9636), .B(n9635), .Z(n9797) );
  XNOR U9936 ( .A(n9796), .B(n9797), .Z(n9798) );
  NANDN U9937 ( .A(n9638), .B(n9637), .Z(n9642) );
  NAND U9938 ( .A(n9640), .B(n9639), .Z(n9641) );
  NAND U9939 ( .A(n9642), .B(n9641), .Z(n9799) );
  XNOR U9940 ( .A(n9798), .B(n9799), .Z(n9856) );
  XNOR U9941 ( .A(n9857), .B(n9856), .Z(n9859) );
  NAND U9942 ( .A(n9644), .B(n9643), .Z(n9648) );
  NAND U9943 ( .A(n9646), .B(n9645), .Z(n9647) );
  AND U9944 ( .A(n9648), .B(n9647), .Z(n9858) );
  XOR U9945 ( .A(n9859), .B(n9858), .Z(n9870) );
  NANDN U9946 ( .A(n9650), .B(n9649), .Z(n9654) );
  NANDN U9947 ( .A(n9652), .B(n9651), .Z(n9653) );
  AND U9948 ( .A(n9654), .B(n9653), .Z(n9868) );
  NANDN U9949 ( .A(n9660), .B(n9659), .Z(n9664) );
  OR U9950 ( .A(n9662), .B(n9661), .Z(n9663) );
  AND U9951 ( .A(n9664), .B(n9663), .Z(n9863) );
  NANDN U9952 ( .A(n9666), .B(n9665), .Z(n9670) );
  NANDN U9953 ( .A(n9668), .B(n9667), .Z(n9669) );
  AND U9954 ( .A(n9670), .B(n9669), .Z(n9803) );
  NANDN U9955 ( .A(n9672), .B(n9671), .Z(n9676) );
  OR U9956 ( .A(n9674), .B(n9673), .Z(n9675) );
  NAND U9957 ( .A(n9676), .B(n9675), .Z(n9802) );
  XNOR U9958 ( .A(n9803), .B(n9802), .Z(n9804) );
  NAND U9959 ( .A(b[0]), .B(a[80]), .Z(n9677) );
  XNOR U9960 ( .A(b[1]), .B(n9677), .Z(n9679) );
  NANDN U9961 ( .A(b[0]), .B(a[79]), .Z(n9678) );
  NAND U9962 ( .A(n9679), .B(n9678), .Z(n9751) );
  NANDN U9963 ( .A(n19394), .B(n9680), .Z(n9682) );
  XOR U9964 ( .A(b[29]), .B(a[52]), .Z(n9826) );
  NANDN U9965 ( .A(n19395), .B(n9826), .Z(n9681) );
  AND U9966 ( .A(n9682), .B(n9681), .Z(n9749) );
  AND U9967 ( .A(b[31]), .B(a[48]), .Z(n9748) );
  XNOR U9968 ( .A(n9749), .B(n9748), .Z(n9750) );
  XNOR U9969 ( .A(n9751), .B(n9750), .Z(n9790) );
  NANDN U9970 ( .A(n19005), .B(n9683), .Z(n9685) );
  XOR U9971 ( .A(b[23]), .B(a[58]), .Z(n9832) );
  NANDN U9972 ( .A(n19055), .B(n9832), .Z(n9684) );
  AND U9973 ( .A(n9685), .B(n9684), .Z(n9823) );
  NANDN U9974 ( .A(n17362), .B(n9686), .Z(n9688) );
  XOR U9975 ( .A(b[7]), .B(a[74]), .Z(n9835) );
  NANDN U9976 ( .A(n17522), .B(n9835), .Z(n9687) );
  AND U9977 ( .A(n9688), .B(n9687), .Z(n9821) );
  NANDN U9978 ( .A(n19116), .B(n9689), .Z(n9691) );
  XOR U9979 ( .A(b[25]), .B(a[56]), .Z(n9838) );
  NANDN U9980 ( .A(n19179), .B(n9838), .Z(n9690) );
  NAND U9981 ( .A(n9691), .B(n9690), .Z(n9820) );
  XNOR U9982 ( .A(n9821), .B(n9820), .Z(n9822) );
  XOR U9983 ( .A(n9823), .B(n9822), .Z(n9791) );
  XNOR U9984 ( .A(n9790), .B(n9791), .Z(n9792) );
  NANDN U9985 ( .A(n18113), .B(n9692), .Z(n9694) );
  XOR U9986 ( .A(b[13]), .B(a[68]), .Z(n9841) );
  NANDN U9987 ( .A(n18229), .B(n9841), .Z(n9693) );
  AND U9988 ( .A(n9694), .B(n9693), .Z(n9785) );
  NANDN U9989 ( .A(n17888), .B(n9695), .Z(n9697) );
  XOR U9990 ( .A(b[11]), .B(a[70]), .Z(n9844) );
  NANDN U9991 ( .A(n18025), .B(n9844), .Z(n9696) );
  NAND U9992 ( .A(n9697), .B(n9696), .Z(n9784) );
  XNOR U9993 ( .A(n9785), .B(n9784), .Z(n9786) );
  NANDN U9994 ( .A(n18487), .B(n9698), .Z(n9700) );
  XOR U9995 ( .A(b[15]), .B(a[66]), .Z(n9847) );
  NANDN U9996 ( .A(n18311), .B(n9847), .Z(n9699) );
  AND U9997 ( .A(n9700), .B(n9699), .Z(n9781) );
  NANDN U9998 ( .A(n18853), .B(n9701), .Z(n9703) );
  XOR U9999 ( .A(b[21]), .B(a[60]), .Z(n9850) );
  NANDN U10000 ( .A(n18926), .B(n9850), .Z(n9702) );
  AND U10001 ( .A(n9703), .B(n9702), .Z(n9779) );
  NANDN U10002 ( .A(n17613), .B(n9704), .Z(n9706) );
  XOR U10003 ( .A(b[9]), .B(a[72]), .Z(n9853) );
  NANDN U10004 ( .A(n17739), .B(n9853), .Z(n9705) );
  NAND U10005 ( .A(n9706), .B(n9705), .Z(n9778) );
  XNOR U10006 ( .A(n9779), .B(n9778), .Z(n9780) );
  XOR U10007 ( .A(n9781), .B(n9780), .Z(n9787) );
  XOR U10008 ( .A(n9786), .B(n9787), .Z(n9793) );
  XOR U10009 ( .A(n9792), .B(n9793), .Z(n9805) );
  XNOR U10010 ( .A(n9804), .B(n9805), .Z(n9862) );
  XNOR U10011 ( .A(n9863), .B(n9862), .Z(n9864) );
  XOR U10012 ( .A(n9865), .B(n9864), .Z(n9869) );
  XOR U10013 ( .A(n9868), .B(n9869), .Z(n9871) );
  XOR U10014 ( .A(n9870), .B(n9871), .Z(n9745) );
  NANDN U10015 ( .A(n9708), .B(n9707), .Z(n9712) );
  NAND U10016 ( .A(n9710), .B(n9709), .Z(n9711) );
  AND U10017 ( .A(n9712), .B(n9711), .Z(n9743) );
  NANDN U10018 ( .A(n9714), .B(n9713), .Z(n9718) );
  NANDN U10019 ( .A(n9716), .B(n9715), .Z(n9717) );
  AND U10020 ( .A(n9718), .B(n9717), .Z(n9742) );
  XNOR U10021 ( .A(n9743), .B(n9742), .Z(n9744) );
  XNOR U10022 ( .A(n9745), .B(n9744), .Z(n9736) );
  NANDN U10023 ( .A(n9720), .B(n9719), .Z(n9724) );
  OR U10024 ( .A(n9722), .B(n9721), .Z(n9723) );
  NAND U10025 ( .A(n9724), .B(n9723), .Z(n9737) );
  XNOR U10026 ( .A(n9736), .B(n9737), .Z(n9738) );
  XNOR U10027 ( .A(n9739), .B(n9738), .Z(n9730) );
  XNOR U10028 ( .A(n9731), .B(n9730), .Z(n9732) );
  XNOR U10029 ( .A(n9733), .B(n9732), .Z(n9874) );
  XNOR U10030 ( .A(sreg[176]), .B(n9874), .Z(n9876) );
  NANDN U10031 ( .A(sreg[175]), .B(n9725), .Z(n9729) );
  NAND U10032 ( .A(n9727), .B(n9726), .Z(n9728) );
  NAND U10033 ( .A(n9729), .B(n9728), .Z(n9875) );
  XNOR U10034 ( .A(n9876), .B(n9875), .Z(c[176]) );
  NANDN U10035 ( .A(n9731), .B(n9730), .Z(n9735) );
  NANDN U10036 ( .A(n9733), .B(n9732), .Z(n9734) );
  AND U10037 ( .A(n9735), .B(n9734), .Z(n9882) );
  NANDN U10038 ( .A(n9737), .B(n9736), .Z(n9741) );
  NANDN U10039 ( .A(n9739), .B(n9738), .Z(n9740) );
  AND U10040 ( .A(n9741), .B(n9740), .Z(n9880) );
  NANDN U10041 ( .A(n9743), .B(n9742), .Z(n9747) );
  NANDN U10042 ( .A(n9745), .B(n9744), .Z(n9746) );
  AND U10043 ( .A(n9747), .B(n9746), .Z(n9888) );
  NANDN U10044 ( .A(n9749), .B(n9748), .Z(n9753) );
  NANDN U10045 ( .A(n9751), .B(n9750), .Z(n9752) );
  AND U10046 ( .A(n9753), .B(n9752), .Z(n9969) );
  NANDN U10047 ( .A(n19237), .B(n9754), .Z(n9756) );
  XOR U10048 ( .A(b[27]), .B(a[55]), .Z(n9915) );
  NANDN U10049 ( .A(n19277), .B(n9915), .Z(n9755) );
  AND U10050 ( .A(n9756), .B(n9755), .Z(n9976) );
  NANDN U10051 ( .A(n17072), .B(n9757), .Z(n9759) );
  XOR U10052 ( .A(b[5]), .B(a[77]), .Z(n9918) );
  NANDN U10053 ( .A(n17223), .B(n9918), .Z(n9758) );
  AND U10054 ( .A(n9759), .B(n9758), .Z(n9974) );
  NANDN U10055 ( .A(n18673), .B(n9760), .Z(n9762) );
  XOR U10056 ( .A(b[19]), .B(a[63]), .Z(n9921) );
  NANDN U10057 ( .A(n18758), .B(n9921), .Z(n9761) );
  NAND U10058 ( .A(n9762), .B(n9761), .Z(n9973) );
  XNOR U10059 ( .A(n9974), .B(n9973), .Z(n9975) );
  XNOR U10060 ( .A(n9976), .B(n9975), .Z(n9967) );
  NANDN U10061 ( .A(n19425), .B(n9763), .Z(n9765) );
  XOR U10062 ( .A(b[31]), .B(a[51]), .Z(n9924) );
  NANDN U10063 ( .A(n19426), .B(n9924), .Z(n9764) );
  AND U10064 ( .A(n9765), .B(n9764), .Z(n9936) );
  NANDN U10065 ( .A(n17067), .B(n9766), .Z(n9768) );
  XOR U10066 ( .A(b[3]), .B(a[79]), .Z(n9927) );
  NANDN U10067 ( .A(n17068), .B(n9927), .Z(n9767) );
  AND U10068 ( .A(n9768), .B(n9767), .Z(n9934) );
  NANDN U10069 ( .A(n18514), .B(n9769), .Z(n9771) );
  XOR U10070 ( .A(b[17]), .B(a[65]), .Z(n9930) );
  NANDN U10071 ( .A(n18585), .B(n9930), .Z(n9770) );
  NAND U10072 ( .A(n9771), .B(n9770), .Z(n9933) );
  XNOR U10073 ( .A(n9934), .B(n9933), .Z(n9935) );
  XOR U10074 ( .A(n9936), .B(n9935), .Z(n9968) );
  XOR U10075 ( .A(n9967), .B(n9968), .Z(n9970) );
  XOR U10076 ( .A(n9969), .B(n9970), .Z(n9904) );
  NANDN U10077 ( .A(n9773), .B(n9772), .Z(n9777) );
  NANDN U10078 ( .A(n9775), .B(n9774), .Z(n9776) );
  AND U10079 ( .A(n9777), .B(n9776), .Z(n9957) );
  NANDN U10080 ( .A(n9779), .B(n9778), .Z(n9783) );
  NANDN U10081 ( .A(n9781), .B(n9780), .Z(n9782) );
  NAND U10082 ( .A(n9783), .B(n9782), .Z(n9958) );
  XNOR U10083 ( .A(n9957), .B(n9958), .Z(n9959) );
  NANDN U10084 ( .A(n9785), .B(n9784), .Z(n9789) );
  NANDN U10085 ( .A(n9787), .B(n9786), .Z(n9788) );
  NAND U10086 ( .A(n9789), .B(n9788), .Z(n9960) );
  XNOR U10087 ( .A(n9959), .B(n9960), .Z(n9903) );
  XNOR U10088 ( .A(n9904), .B(n9903), .Z(n9906) );
  NANDN U10089 ( .A(n9791), .B(n9790), .Z(n9795) );
  NANDN U10090 ( .A(n9793), .B(n9792), .Z(n9794) );
  AND U10091 ( .A(n9795), .B(n9794), .Z(n9905) );
  XOR U10092 ( .A(n9906), .B(n9905), .Z(n10017) );
  NANDN U10093 ( .A(n9797), .B(n9796), .Z(n9801) );
  NANDN U10094 ( .A(n9799), .B(n9798), .Z(n9800) );
  AND U10095 ( .A(n9801), .B(n9800), .Z(n10015) );
  NANDN U10096 ( .A(n9803), .B(n9802), .Z(n9807) );
  NANDN U10097 ( .A(n9805), .B(n9804), .Z(n9806) );
  AND U10098 ( .A(n9807), .B(n9806), .Z(n9900) );
  NANDN U10099 ( .A(n9809), .B(n9808), .Z(n9813) );
  OR U10100 ( .A(n9811), .B(n9810), .Z(n9812) );
  AND U10101 ( .A(n9813), .B(n9812), .Z(n9898) );
  NANDN U10102 ( .A(n9815), .B(n9814), .Z(n9819) );
  NANDN U10103 ( .A(n9817), .B(n9816), .Z(n9818) );
  AND U10104 ( .A(n9819), .B(n9818), .Z(n9964) );
  NANDN U10105 ( .A(n9821), .B(n9820), .Z(n9825) );
  NANDN U10106 ( .A(n9823), .B(n9822), .Z(n9824) );
  NAND U10107 ( .A(n9825), .B(n9824), .Z(n9963) );
  XNOR U10108 ( .A(n9964), .B(n9963), .Z(n9966) );
  NANDN U10109 ( .A(n19394), .B(n9826), .Z(n9828) );
  XOR U10110 ( .A(b[29]), .B(a[53]), .Z(n9988) );
  NANDN U10111 ( .A(n19395), .B(n9988), .Z(n9827) );
  AND U10112 ( .A(n9828), .B(n9827), .Z(n9910) );
  AND U10113 ( .A(b[31]), .B(a[49]), .Z(n9909) );
  XNOR U10114 ( .A(n9910), .B(n9909), .Z(n9911) );
  NAND U10115 ( .A(b[0]), .B(a[81]), .Z(n9829) );
  XNOR U10116 ( .A(b[1]), .B(n9829), .Z(n9831) );
  NANDN U10117 ( .A(b[0]), .B(a[80]), .Z(n9830) );
  NAND U10118 ( .A(n9831), .B(n9830), .Z(n9912) );
  XNOR U10119 ( .A(n9911), .B(n9912), .Z(n9952) );
  NANDN U10120 ( .A(n19005), .B(n9832), .Z(n9834) );
  XOR U10121 ( .A(b[23]), .B(a[59]), .Z(n9991) );
  NANDN U10122 ( .A(n19055), .B(n9991), .Z(n9833) );
  AND U10123 ( .A(n9834), .B(n9833), .Z(n9981) );
  NANDN U10124 ( .A(n17362), .B(n9835), .Z(n9837) );
  XOR U10125 ( .A(b[7]), .B(a[75]), .Z(n9994) );
  NANDN U10126 ( .A(n17522), .B(n9994), .Z(n9836) );
  AND U10127 ( .A(n9837), .B(n9836), .Z(n9980) );
  NANDN U10128 ( .A(n19116), .B(n9838), .Z(n9840) );
  XOR U10129 ( .A(b[25]), .B(a[57]), .Z(n9997) );
  NANDN U10130 ( .A(n19179), .B(n9997), .Z(n9839) );
  NAND U10131 ( .A(n9840), .B(n9839), .Z(n9979) );
  XOR U10132 ( .A(n9980), .B(n9979), .Z(n9982) );
  XOR U10133 ( .A(n9981), .B(n9982), .Z(n9951) );
  XOR U10134 ( .A(n9952), .B(n9951), .Z(n9954) );
  NANDN U10135 ( .A(n18113), .B(n9841), .Z(n9843) );
  XOR U10136 ( .A(b[13]), .B(a[69]), .Z(n10000) );
  NANDN U10137 ( .A(n18229), .B(n10000), .Z(n9842) );
  AND U10138 ( .A(n9843), .B(n9842), .Z(n9946) );
  NANDN U10139 ( .A(n17888), .B(n9844), .Z(n9846) );
  XOR U10140 ( .A(b[11]), .B(a[71]), .Z(n10003) );
  NANDN U10141 ( .A(n18025), .B(n10003), .Z(n9845) );
  NAND U10142 ( .A(n9846), .B(n9845), .Z(n9945) );
  XNOR U10143 ( .A(n9946), .B(n9945), .Z(n9948) );
  NANDN U10144 ( .A(n18487), .B(n9847), .Z(n9849) );
  XOR U10145 ( .A(b[15]), .B(a[67]), .Z(n10006) );
  NANDN U10146 ( .A(n18311), .B(n10006), .Z(n9848) );
  AND U10147 ( .A(n9849), .B(n9848), .Z(n9942) );
  NANDN U10148 ( .A(n18853), .B(n9850), .Z(n9852) );
  XOR U10149 ( .A(b[21]), .B(a[61]), .Z(n10009) );
  NANDN U10150 ( .A(n18926), .B(n10009), .Z(n9851) );
  AND U10151 ( .A(n9852), .B(n9851), .Z(n9940) );
  NANDN U10152 ( .A(n17613), .B(n9853), .Z(n9855) );
  XOR U10153 ( .A(b[9]), .B(a[73]), .Z(n10012) );
  NANDN U10154 ( .A(n17739), .B(n10012), .Z(n9854) );
  NAND U10155 ( .A(n9855), .B(n9854), .Z(n9939) );
  XNOR U10156 ( .A(n9940), .B(n9939), .Z(n9941) );
  XNOR U10157 ( .A(n9942), .B(n9941), .Z(n9947) );
  XOR U10158 ( .A(n9948), .B(n9947), .Z(n9953) );
  XOR U10159 ( .A(n9954), .B(n9953), .Z(n9965) );
  XOR U10160 ( .A(n9966), .B(n9965), .Z(n9897) );
  XNOR U10161 ( .A(n9898), .B(n9897), .Z(n9899) );
  XOR U10162 ( .A(n9900), .B(n9899), .Z(n10016) );
  XOR U10163 ( .A(n10015), .B(n10016), .Z(n10018) );
  XOR U10164 ( .A(n10017), .B(n10018), .Z(n9894) );
  NANDN U10165 ( .A(n9857), .B(n9856), .Z(n9861) );
  NAND U10166 ( .A(n9859), .B(n9858), .Z(n9860) );
  AND U10167 ( .A(n9861), .B(n9860), .Z(n9892) );
  NANDN U10168 ( .A(n9863), .B(n9862), .Z(n9867) );
  NANDN U10169 ( .A(n9865), .B(n9864), .Z(n9866) );
  AND U10170 ( .A(n9867), .B(n9866), .Z(n9891) );
  XNOR U10171 ( .A(n9892), .B(n9891), .Z(n9893) );
  XNOR U10172 ( .A(n9894), .B(n9893), .Z(n9885) );
  NANDN U10173 ( .A(n9869), .B(n9868), .Z(n9873) );
  OR U10174 ( .A(n9871), .B(n9870), .Z(n9872) );
  NAND U10175 ( .A(n9873), .B(n9872), .Z(n9886) );
  XNOR U10176 ( .A(n9885), .B(n9886), .Z(n9887) );
  XNOR U10177 ( .A(n9888), .B(n9887), .Z(n9879) );
  XNOR U10178 ( .A(n9880), .B(n9879), .Z(n9881) );
  XNOR U10179 ( .A(n9882), .B(n9881), .Z(n10021) );
  XNOR U10180 ( .A(sreg[177]), .B(n10021), .Z(n10023) );
  NANDN U10181 ( .A(sreg[176]), .B(n9874), .Z(n9878) );
  NAND U10182 ( .A(n9876), .B(n9875), .Z(n9877) );
  NAND U10183 ( .A(n9878), .B(n9877), .Z(n10022) );
  XNOR U10184 ( .A(n10023), .B(n10022), .Z(c[177]) );
  NANDN U10185 ( .A(n9880), .B(n9879), .Z(n9884) );
  NANDN U10186 ( .A(n9882), .B(n9881), .Z(n9883) );
  AND U10187 ( .A(n9884), .B(n9883), .Z(n10029) );
  NANDN U10188 ( .A(n9886), .B(n9885), .Z(n9890) );
  NANDN U10189 ( .A(n9888), .B(n9887), .Z(n9889) );
  AND U10190 ( .A(n9890), .B(n9889), .Z(n10027) );
  NANDN U10191 ( .A(n9892), .B(n9891), .Z(n9896) );
  NANDN U10192 ( .A(n9894), .B(n9893), .Z(n9895) );
  AND U10193 ( .A(n9896), .B(n9895), .Z(n10035) );
  NANDN U10194 ( .A(n9898), .B(n9897), .Z(n9902) );
  NANDN U10195 ( .A(n9900), .B(n9899), .Z(n9901) );
  AND U10196 ( .A(n9902), .B(n9901), .Z(n10163) );
  NANDN U10197 ( .A(n9904), .B(n9903), .Z(n9908) );
  NAND U10198 ( .A(n9906), .B(n9905), .Z(n9907) );
  AND U10199 ( .A(n9908), .B(n9907), .Z(n10162) );
  XNOR U10200 ( .A(n10163), .B(n10162), .Z(n10165) );
  NANDN U10201 ( .A(n9910), .B(n9909), .Z(n9914) );
  NANDN U10202 ( .A(n9912), .B(n9911), .Z(n9913) );
  AND U10203 ( .A(n9914), .B(n9913), .Z(n10098) );
  NANDN U10204 ( .A(n19237), .B(n9915), .Z(n9917) );
  XOR U10205 ( .A(b[27]), .B(a[56]), .Z(n10044) );
  NANDN U10206 ( .A(n19277), .B(n10044), .Z(n9916) );
  AND U10207 ( .A(n9917), .B(n9916), .Z(n10105) );
  NANDN U10208 ( .A(n17072), .B(n9918), .Z(n9920) );
  XOR U10209 ( .A(b[5]), .B(a[78]), .Z(n10047) );
  NANDN U10210 ( .A(n17223), .B(n10047), .Z(n9919) );
  AND U10211 ( .A(n9920), .B(n9919), .Z(n10103) );
  NANDN U10212 ( .A(n18673), .B(n9921), .Z(n9923) );
  XOR U10213 ( .A(b[19]), .B(a[64]), .Z(n10050) );
  NANDN U10214 ( .A(n18758), .B(n10050), .Z(n9922) );
  NAND U10215 ( .A(n9923), .B(n9922), .Z(n10102) );
  XNOR U10216 ( .A(n10103), .B(n10102), .Z(n10104) );
  XNOR U10217 ( .A(n10105), .B(n10104), .Z(n10096) );
  NANDN U10218 ( .A(n19425), .B(n9924), .Z(n9926) );
  XOR U10219 ( .A(b[31]), .B(a[52]), .Z(n10053) );
  NANDN U10220 ( .A(n19426), .B(n10053), .Z(n9925) );
  AND U10221 ( .A(n9926), .B(n9925), .Z(n10065) );
  NANDN U10222 ( .A(n17067), .B(n9927), .Z(n9929) );
  XOR U10223 ( .A(b[3]), .B(a[80]), .Z(n10056) );
  NANDN U10224 ( .A(n17068), .B(n10056), .Z(n9928) );
  AND U10225 ( .A(n9929), .B(n9928), .Z(n10063) );
  NANDN U10226 ( .A(n18514), .B(n9930), .Z(n9932) );
  XOR U10227 ( .A(b[17]), .B(a[66]), .Z(n10059) );
  NANDN U10228 ( .A(n18585), .B(n10059), .Z(n9931) );
  NAND U10229 ( .A(n9932), .B(n9931), .Z(n10062) );
  XNOR U10230 ( .A(n10063), .B(n10062), .Z(n10064) );
  XOR U10231 ( .A(n10065), .B(n10064), .Z(n10097) );
  XOR U10232 ( .A(n10096), .B(n10097), .Z(n10099) );
  XOR U10233 ( .A(n10098), .B(n10099), .Z(n10145) );
  NANDN U10234 ( .A(n9934), .B(n9933), .Z(n9938) );
  NANDN U10235 ( .A(n9936), .B(n9935), .Z(n9937) );
  AND U10236 ( .A(n9938), .B(n9937), .Z(n10086) );
  NANDN U10237 ( .A(n9940), .B(n9939), .Z(n9944) );
  NANDN U10238 ( .A(n9942), .B(n9941), .Z(n9943) );
  NAND U10239 ( .A(n9944), .B(n9943), .Z(n10087) );
  XNOR U10240 ( .A(n10086), .B(n10087), .Z(n10088) );
  NANDN U10241 ( .A(n9946), .B(n9945), .Z(n9950) );
  NAND U10242 ( .A(n9948), .B(n9947), .Z(n9949) );
  NAND U10243 ( .A(n9950), .B(n9949), .Z(n10089) );
  XNOR U10244 ( .A(n10088), .B(n10089), .Z(n10144) );
  XNOR U10245 ( .A(n10145), .B(n10144), .Z(n10147) );
  NAND U10246 ( .A(n9952), .B(n9951), .Z(n9956) );
  NAND U10247 ( .A(n9954), .B(n9953), .Z(n9955) );
  AND U10248 ( .A(n9956), .B(n9955), .Z(n10146) );
  XOR U10249 ( .A(n10147), .B(n10146), .Z(n10159) );
  NANDN U10250 ( .A(n9958), .B(n9957), .Z(n9962) );
  NANDN U10251 ( .A(n9960), .B(n9959), .Z(n9961) );
  AND U10252 ( .A(n9962), .B(n9961), .Z(n10156) );
  NANDN U10253 ( .A(n9968), .B(n9967), .Z(n9972) );
  OR U10254 ( .A(n9970), .B(n9969), .Z(n9971) );
  AND U10255 ( .A(n9972), .B(n9971), .Z(n10151) );
  NANDN U10256 ( .A(n9974), .B(n9973), .Z(n9978) );
  NANDN U10257 ( .A(n9976), .B(n9975), .Z(n9977) );
  AND U10258 ( .A(n9978), .B(n9977), .Z(n10093) );
  NANDN U10259 ( .A(n9980), .B(n9979), .Z(n9984) );
  OR U10260 ( .A(n9982), .B(n9981), .Z(n9983) );
  NAND U10261 ( .A(n9984), .B(n9983), .Z(n10092) );
  XNOR U10262 ( .A(n10093), .B(n10092), .Z(n10095) );
  NAND U10263 ( .A(b[0]), .B(a[82]), .Z(n9985) );
  XNOR U10264 ( .A(b[1]), .B(n9985), .Z(n9987) );
  NANDN U10265 ( .A(b[0]), .B(a[81]), .Z(n9986) );
  NAND U10266 ( .A(n9987), .B(n9986), .Z(n10041) );
  NANDN U10267 ( .A(n19394), .B(n9988), .Z(n9990) );
  XOR U10268 ( .A(b[29]), .B(a[54]), .Z(n10117) );
  NANDN U10269 ( .A(n19395), .B(n10117), .Z(n9989) );
  AND U10270 ( .A(n9990), .B(n9989), .Z(n10039) );
  AND U10271 ( .A(b[31]), .B(a[50]), .Z(n10038) );
  XNOR U10272 ( .A(n10039), .B(n10038), .Z(n10040) );
  XNOR U10273 ( .A(n10041), .B(n10040), .Z(n10081) );
  NANDN U10274 ( .A(n19005), .B(n9991), .Z(n9993) );
  XOR U10275 ( .A(b[23]), .B(a[60]), .Z(n10120) );
  NANDN U10276 ( .A(n19055), .B(n10120), .Z(n9992) );
  AND U10277 ( .A(n9993), .B(n9992), .Z(n10110) );
  NANDN U10278 ( .A(n17362), .B(n9994), .Z(n9996) );
  XOR U10279 ( .A(b[7]), .B(a[76]), .Z(n10123) );
  NANDN U10280 ( .A(n17522), .B(n10123), .Z(n9995) );
  AND U10281 ( .A(n9996), .B(n9995), .Z(n10109) );
  NANDN U10282 ( .A(n19116), .B(n9997), .Z(n9999) );
  XOR U10283 ( .A(b[25]), .B(a[58]), .Z(n10126) );
  NANDN U10284 ( .A(n19179), .B(n10126), .Z(n9998) );
  NAND U10285 ( .A(n9999), .B(n9998), .Z(n10108) );
  XOR U10286 ( .A(n10109), .B(n10108), .Z(n10111) );
  XOR U10287 ( .A(n10110), .B(n10111), .Z(n10080) );
  XOR U10288 ( .A(n10081), .B(n10080), .Z(n10083) );
  NANDN U10289 ( .A(n18113), .B(n10000), .Z(n10002) );
  XOR U10290 ( .A(b[13]), .B(a[70]), .Z(n10129) );
  NANDN U10291 ( .A(n18229), .B(n10129), .Z(n10001) );
  AND U10292 ( .A(n10002), .B(n10001), .Z(n10075) );
  NANDN U10293 ( .A(n17888), .B(n10003), .Z(n10005) );
  XOR U10294 ( .A(b[11]), .B(a[72]), .Z(n10132) );
  NANDN U10295 ( .A(n18025), .B(n10132), .Z(n10004) );
  NAND U10296 ( .A(n10005), .B(n10004), .Z(n10074) );
  XNOR U10297 ( .A(n10075), .B(n10074), .Z(n10077) );
  NANDN U10298 ( .A(n18487), .B(n10006), .Z(n10008) );
  XOR U10299 ( .A(b[15]), .B(a[68]), .Z(n10135) );
  NANDN U10300 ( .A(n18311), .B(n10135), .Z(n10007) );
  AND U10301 ( .A(n10008), .B(n10007), .Z(n10071) );
  NANDN U10302 ( .A(n18853), .B(n10009), .Z(n10011) );
  XOR U10303 ( .A(b[21]), .B(a[62]), .Z(n10138) );
  NANDN U10304 ( .A(n18926), .B(n10138), .Z(n10010) );
  AND U10305 ( .A(n10011), .B(n10010), .Z(n10069) );
  NANDN U10306 ( .A(n17613), .B(n10012), .Z(n10014) );
  XOR U10307 ( .A(b[9]), .B(a[74]), .Z(n10141) );
  NANDN U10308 ( .A(n17739), .B(n10141), .Z(n10013) );
  NAND U10309 ( .A(n10014), .B(n10013), .Z(n10068) );
  XNOR U10310 ( .A(n10069), .B(n10068), .Z(n10070) );
  XNOR U10311 ( .A(n10071), .B(n10070), .Z(n10076) );
  XOR U10312 ( .A(n10077), .B(n10076), .Z(n10082) );
  XOR U10313 ( .A(n10083), .B(n10082), .Z(n10094) );
  XOR U10314 ( .A(n10095), .B(n10094), .Z(n10150) );
  XNOR U10315 ( .A(n10151), .B(n10150), .Z(n10152) );
  XOR U10316 ( .A(n10153), .B(n10152), .Z(n10157) );
  XNOR U10317 ( .A(n10156), .B(n10157), .Z(n10158) );
  XNOR U10318 ( .A(n10159), .B(n10158), .Z(n10164) );
  XOR U10319 ( .A(n10165), .B(n10164), .Z(n10033) );
  NANDN U10320 ( .A(n10016), .B(n10015), .Z(n10020) );
  OR U10321 ( .A(n10018), .B(n10017), .Z(n10019) );
  AND U10322 ( .A(n10020), .B(n10019), .Z(n10032) );
  XNOR U10323 ( .A(n10033), .B(n10032), .Z(n10034) );
  XNOR U10324 ( .A(n10035), .B(n10034), .Z(n10026) );
  XNOR U10325 ( .A(n10027), .B(n10026), .Z(n10028) );
  XNOR U10326 ( .A(n10029), .B(n10028), .Z(n10168) );
  XNOR U10327 ( .A(sreg[178]), .B(n10168), .Z(n10170) );
  NANDN U10328 ( .A(sreg[177]), .B(n10021), .Z(n10025) );
  NAND U10329 ( .A(n10023), .B(n10022), .Z(n10024) );
  NAND U10330 ( .A(n10025), .B(n10024), .Z(n10169) );
  XNOR U10331 ( .A(n10170), .B(n10169), .Z(c[178]) );
  NANDN U10332 ( .A(n10027), .B(n10026), .Z(n10031) );
  NANDN U10333 ( .A(n10029), .B(n10028), .Z(n10030) );
  AND U10334 ( .A(n10031), .B(n10030), .Z(n10176) );
  NANDN U10335 ( .A(n10033), .B(n10032), .Z(n10037) );
  NANDN U10336 ( .A(n10035), .B(n10034), .Z(n10036) );
  AND U10337 ( .A(n10037), .B(n10036), .Z(n10174) );
  NANDN U10338 ( .A(n10039), .B(n10038), .Z(n10043) );
  NANDN U10339 ( .A(n10041), .B(n10040), .Z(n10042) );
  AND U10340 ( .A(n10043), .B(n10042), .Z(n10251) );
  NANDN U10341 ( .A(n19237), .B(n10044), .Z(n10046) );
  XOR U10342 ( .A(b[27]), .B(a[57]), .Z(n10197) );
  NANDN U10343 ( .A(n19277), .B(n10197), .Z(n10045) );
  AND U10344 ( .A(n10046), .B(n10045), .Z(n10258) );
  NANDN U10345 ( .A(n17072), .B(n10047), .Z(n10049) );
  XOR U10346 ( .A(b[5]), .B(a[79]), .Z(n10200) );
  NANDN U10347 ( .A(n17223), .B(n10200), .Z(n10048) );
  AND U10348 ( .A(n10049), .B(n10048), .Z(n10256) );
  NANDN U10349 ( .A(n18673), .B(n10050), .Z(n10052) );
  XOR U10350 ( .A(b[19]), .B(a[65]), .Z(n10203) );
  NANDN U10351 ( .A(n18758), .B(n10203), .Z(n10051) );
  NAND U10352 ( .A(n10052), .B(n10051), .Z(n10255) );
  XNOR U10353 ( .A(n10256), .B(n10255), .Z(n10257) );
  XNOR U10354 ( .A(n10258), .B(n10257), .Z(n10249) );
  NANDN U10355 ( .A(n19425), .B(n10053), .Z(n10055) );
  XOR U10356 ( .A(b[31]), .B(a[53]), .Z(n10206) );
  NANDN U10357 ( .A(n19426), .B(n10206), .Z(n10054) );
  AND U10358 ( .A(n10055), .B(n10054), .Z(n10218) );
  NANDN U10359 ( .A(n17067), .B(n10056), .Z(n10058) );
  XOR U10360 ( .A(b[3]), .B(a[81]), .Z(n10209) );
  NANDN U10361 ( .A(n17068), .B(n10209), .Z(n10057) );
  AND U10362 ( .A(n10058), .B(n10057), .Z(n10216) );
  NANDN U10363 ( .A(n18514), .B(n10059), .Z(n10061) );
  XOR U10364 ( .A(b[17]), .B(a[67]), .Z(n10212) );
  NANDN U10365 ( .A(n18585), .B(n10212), .Z(n10060) );
  NAND U10366 ( .A(n10061), .B(n10060), .Z(n10215) );
  XNOR U10367 ( .A(n10216), .B(n10215), .Z(n10217) );
  XOR U10368 ( .A(n10218), .B(n10217), .Z(n10250) );
  XOR U10369 ( .A(n10249), .B(n10250), .Z(n10252) );
  XOR U10370 ( .A(n10251), .B(n10252), .Z(n10298) );
  NANDN U10371 ( .A(n10063), .B(n10062), .Z(n10067) );
  NANDN U10372 ( .A(n10065), .B(n10064), .Z(n10066) );
  AND U10373 ( .A(n10067), .B(n10066), .Z(n10239) );
  NANDN U10374 ( .A(n10069), .B(n10068), .Z(n10073) );
  NANDN U10375 ( .A(n10071), .B(n10070), .Z(n10072) );
  NAND U10376 ( .A(n10073), .B(n10072), .Z(n10240) );
  XNOR U10377 ( .A(n10239), .B(n10240), .Z(n10241) );
  NANDN U10378 ( .A(n10075), .B(n10074), .Z(n10079) );
  NAND U10379 ( .A(n10077), .B(n10076), .Z(n10078) );
  NAND U10380 ( .A(n10079), .B(n10078), .Z(n10242) );
  XNOR U10381 ( .A(n10241), .B(n10242), .Z(n10297) );
  XNOR U10382 ( .A(n10298), .B(n10297), .Z(n10300) );
  NAND U10383 ( .A(n10081), .B(n10080), .Z(n10085) );
  NAND U10384 ( .A(n10083), .B(n10082), .Z(n10084) );
  AND U10385 ( .A(n10085), .B(n10084), .Z(n10299) );
  XOR U10386 ( .A(n10300), .B(n10299), .Z(n10311) );
  NANDN U10387 ( .A(n10087), .B(n10086), .Z(n10091) );
  NANDN U10388 ( .A(n10089), .B(n10088), .Z(n10090) );
  AND U10389 ( .A(n10091), .B(n10090), .Z(n10309) );
  NANDN U10390 ( .A(n10097), .B(n10096), .Z(n10101) );
  OR U10391 ( .A(n10099), .B(n10098), .Z(n10100) );
  AND U10392 ( .A(n10101), .B(n10100), .Z(n10304) );
  NANDN U10393 ( .A(n10103), .B(n10102), .Z(n10107) );
  NANDN U10394 ( .A(n10105), .B(n10104), .Z(n10106) );
  AND U10395 ( .A(n10107), .B(n10106), .Z(n10246) );
  NANDN U10396 ( .A(n10109), .B(n10108), .Z(n10113) );
  OR U10397 ( .A(n10111), .B(n10110), .Z(n10112) );
  NAND U10398 ( .A(n10113), .B(n10112), .Z(n10245) );
  XNOR U10399 ( .A(n10246), .B(n10245), .Z(n10248) );
  NAND U10400 ( .A(b[0]), .B(a[83]), .Z(n10114) );
  XNOR U10401 ( .A(b[1]), .B(n10114), .Z(n10116) );
  NANDN U10402 ( .A(b[0]), .B(a[82]), .Z(n10115) );
  NAND U10403 ( .A(n10116), .B(n10115), .Z(n10194) );
  NANDN U10404 ( .A(n19394), .B(n10117), .Z(n10119) );
  XOR U10405 ( .A(b[29]), .B(a[55]), .Z(n10270) );
  NANDN U10406 ( .A(n19395), .B(n10270), .Z(n10118) );
  AND U10407 ( .A(n10119), .B(n10118), .Z(n10192) );
  AND U10408 ( .A(b[31]), .B(a[51]), .Z(n10191) );
  XNOR U10409 ( .A(n10192), .B(n10191), .Z(n10193) );
  XNOR U10410 ( .A(n10194), .B(n10193), .Z(n10234) );
  NANDN U10411 ( .A(n19005), .B(n10120), .Z(n10122) );
  XOR U10412 ( .A(b[23]), .B(a[61]), .Z(n10273) );
  NANDN U10413 ( .A(n19055), .B(n10273), .Z(n10121) );
  AND U10414 ( .A(n10122), .B(n10121), .Z(n10263) );
  NANDN U10415 ( .A(n17362), .B(n10123), .Z(n10125) );
  XOR U10416 ( .A(b[7]), .B(a[77]), .Z(n10276) );
  NANDN U10417 ( .A(n17522), .B(n10276), .Z(n10124) );
  AND U10418 ( .A(n10125), .B(n10124), .Z(n10262) );
  NANDN U10419 ( .A(n19116), .B(n10126), .Z(n10128) );
  XOR U10420 ( .A(b[25]), .B(a[59]), .Z(n10279) );
  NANDN U10421 ( .A(n19179), .B(n10279), .Z(n10127) );
  NAND U10422 ( .A(n10128), .B(n10127), .Z(n10261) );
  XOR U10423 ( .A(n10262), .B(n10261), .Z(n10264) );
  XOR U10424 ( .A(n10263), .B(n10264), .Z(n10233) );
  XOR U10425 ( .A(n10234), .B(n10233), .Z(n10236) );
  NANDN U10426 ( .A(n18113), .B(n10129), .Z(n10131) );
  XOR U10427 ( .A(b[13]), .B(a[71]), .Z(n10282) );
  NANDN U10428 ( .A(n18229), .B(n10282), .Z(n10130) );
  AND U10429 ( .A(n10131), .B(n10130), .Z(n10228) );
  NANDN U10430 ( .A(n17888), .B(n10132), .Z(n10134) );
  XOR U10431 ( .A(b[11]), .B(a[73]), .Z(n10285) );
  NANDN U10432 ( .A(n18025), .B(n10285), .Z(n10133) );
  NAND U10433 ( .A(n10134), .B(n10133), .Z(n10227) );
  XNOR U10434 ( .A(n10228), .B(n10227), .Z(n10230) );
  NANDN U10435 ( .A(n18487), .B(n10135), .Z(n10137) );
  XOR U10436 ( .A(b[15]), .B(a[69]), .Z(n10288) );
  NANDN U10437 ( .A(n18311), .B(n10288), .Z(n10136) );
  AND U10438 ( .A(n10137), .B(n10136), .Z(n10224) );
  NANDN U10439 ( .A(n18853), .B(n10138), .Z(n10140) );
  XOR U10440 ( .A(b[21]), .B(a[63]), .Z(n10291) );
  NANDN U10441 ( .A(n18926), .B(n10291), .Z(n10139) );
  AND U10442 ( .A(n10140), .B(n10139), .Z(n10222) );
  NANDN U10443 ( .A(n17613), .B(n10141), .Z(n10143) );
  XOR U10444 ( .A(b[9]), .B(a[75]), .Z(n10294) );
  NANDN U10445 ( .A(n17739), .B(n10294), .Z(n10142) );
  NAND U10446 ( .A(n10143), .B(n10142), .Z(n10221) );
  XNOR U10447 ( .A(n10222), .B(n10221), .Z(n10223) );
  XNOR U10448 ( .A(n10224), .B(n10223), .Z(n10229) );
  XOR U10449 ( .A(n10230), .B(n10229), .Z(n10235) );
  XOR U10450 ( .A(n10236), .B(n10235), .Z(n10247) );
  XOR U10451 ( .A(n10248), .B(n10247), .Z(n10303) );
  XNOR U10452 ( .A(n10304), .B(n10303), .Z(n10305) );
  XOR U10453 ( .A(n10306), .B(n10305), .Z(n10310) );
  XOR U10454 ( .A(n10309), .B(n10310), .Z(n10312) );
  XOR U10455 ( .A(n10311), .B(n10312), .Z(n10188) );
  NANDN U10456 ( .A(n10145), .B(n10144), .Z(n10149) );
  NAND U10457 ( .A(n10147), .B(n10146), .Z(n10148) );
  AND U10458 ( .A(n10149), .B(n10148), .Z(n10186) );
  NANDN U10459 ( .A(n10151), .B(n10150), .Z(n10155) );
  NANDN U10460 ( .A(n10153), .B(n10152), .Z(n10154) );
  AND U10461 ( .A(n10155), .B(n10154), .Z(n10185) );
  XNOR U10462 ( .A(n10186), .B(n10185), .Z(n10187) );
  XNOR U10463 ( .A(n10188), .B(n10187), .Z(n10179) );
  NANDN U10464 ( .A(n10157), .B(n10156), .Z(n10161) );
  NANDN U10465 ( .A(n10159), .B(n10158), .Z(n10160) );
  NAND U10466 ( .A(n10161), .B(n10160), .Z(n10180) );
  XNOR U10467 ( .A(n10179), .B(n10180), .Z(n10181) );
  NANDN U10468 ( .A(n10163), .B(n10162), .Z(n10167) );
  NAND U10469 ( .A(n10165), .B(n10164), .Z(n10166) );
  NAND U10470 ( .A(n10167), .B(n10166), .Z(n10182) );
  XNOR U10471 ( .A(n10181), .B(n10182), .Z(n10173) );
  XNOR U10472 ( .A(n10174), .B(n10173), .Z(n10175) );
  XNOR U10473 ( .A(n10176), .B(n10175), .Z(n10315) );
  XNOR U10474 ( .A(sreg[179]), .B(n10315), .Z(n10317) );
  NANDN U10475 ( .A(sreg[178]), .B(n10168), .Z(n10172) );
  NAND U10476 ( .A(n10170), .B(n10169), .Z(n10171) );
  NAND U10477 ( .A(n10172), .B(n10171), .Z(n10316) );
  XNOR U10478 ( .A(n10317), .B(n10316), .Z(c[179]) );
  NANDN U10479 ( .A(n10174), .B(n10173), .Z(n10178) );
  NANDN U10480 ( .A(n10176), .B(n10175), .Z(n10177) );
  AND U10481 ( .A(n10178), .B(n10177), .Z(n10323) );
  NANDN U10482 ( .A(n10180), .B(n10179), .Z(n10184) );
  NANDN U10483 ( .A(n10182), .B(n10181), .Z(n10183) );
  AND U10484 ( .A(n10184), .B(n10183), .Z(n10321) );
  NANDN U10485 ( .A(n10186), .B(n10185), .Z(n10190) );
  NANDN U10486 ( .A(n10188), .B(n10187), .Z(n10189) );
  AND U10487 ( .A(n10190), .B(n10189), .Z(n10329) );
  NANDN U10488 ( .A(n10192), .B(n10191), .Z(n10196) );
  NANDN U10489 ( .A(n10194), .B(n10193), .Z(n10195) );
  AND U10490 ( .A(n10196), .B(n10195), .Z(n10400) );
  NANDN U10491 ( .A(n19237), .B(n10197), .Z(n10199) );
  XOR U10492 ( .A(b[27]), .B(a[58]), .Z(n10344) );
  NANDN U10493 ( .A(n19277), .B(n10344), .Z(n10198) );
  AND U10494 ( .A(n10199), .B(n10198), .Z(n10407) );
  NANDN U10495 ( .A(n17072), .B(n10200), .Z(n10202) );
  XOR U10496 ( .A(b[5]), .B(a[80]), .Z(n10347) );
  NANDN U10497 ( .A(n17223), .B(n10347), .Z(n10201) );
  AND U10498 ( .A(n10202), .B(n10201), .Z(n10405) );
  NANDN U10499 ( .A(n18673), .B(n10203), .Z(n10205) );
  XOR U10500 ( .A(b[19]), .B(a[66]), .Z(n10350) );
  NANDN U10501 ( .A(n18758), .B(n10350), .Z(n10204) );
  NAND U10502 ( .A(n10205), .B(n10204), .Z(n10404) );
  XNOR U10503 ( .A(n10405), .B(n10404), .Z(n10406) );
  XNOR U10504 ( .A(n10407), .B(n10406), .Z(n10398) );
  NANDN U10505 ( .A(n19425), .B(n10206), .Z(n10208) );
  XOR U10506 ( .A(b[31]), .B(a[54]), .Z(n10353) );
  NANDN U10507 ( .A(n19426), .B(n10353), .Z(n10207) );
  AND U10508 ( .A(n10208), .B(n10207), .Z(n10365) );
  NANDN U10509 ( .A(n17067), .B(n10209), .Z(n10211) );
  XOR U10510 ( .A(b[3]), .B(a[82]), .Z(n10356) );
  NANDN U10511 ( .A(n17068), .B(n10356), .Z(n10210) );
  AND U10512 ( .A(n10211), .B(n10210), .Z(n10363) );
  NANDN U10513 ( .A(n18514), .B(n10212), .Z(n10214) );
  XOR U10514 ( .A(b[17]), .B(a[68]), .Z(n10359) );
  NANDN U10515 ( .A(n18585), .B(n10359), .Z(n10213) );
  NAND U10516 ( .A(n10214), .B(n10213), .Z(n10362) );
  XNOR U10517 ( .A(n10363), .B(n10362), .Z(n10364) );
  XOR U10518 ( .A(n10365), .B(n10364), .Z(n10399) );
  XOR U10519 ( .A(n10398), .B(n10399), .Z(n10401) );
  XOR U10520 ( .A(n10400), .B(n10401), .Z(n10447) );
  NANDN U10521 ( .A(n10216), .B(n10215), .Z(n10220) );
  NANDN U10522 ( .A(n10218), .B(n10217), .Z(n10219) );
  AND U10523 ( .A(n10220), .B(n10219), .Z(n10386) );
  NANDN U10524 ( .A(n10222), .B(n10221), .Z(n10226) );
  NANDN U10525 ( .A(n10224), .B(n10223), .Z(n10225) );
  NAND U10526 ( .A(n10226), .B(n10225), .Z(n10387) );
  XNOR U10527 ( .A(n10386), .B(n10387), .Z(n10388) );
  NANDN U10528 ( .A(n10228), .B(n10227), .Z(n10232) );
  NAND U10529 ( .A(n10230), .B(n10229), .Z(n10231) );
  NAND U10530 ( .A(n10232), .B(n10231), .Z(n10389) );
  XNOR U10531 ( .A(n10388), .B(n10389), .Z(n10446) );
  XNOR U10532 ( .A(n10447), .B(n10446), .Z(n10449) );
  NAND U10533 ( .A(n10234), .B(n10233), .Z(n10238) );
  NAND U10534 ( .A(n10236), .B(n10235), .Z(n10237) );
  AND U10535 ( .A(n10238), .B(n10237), .Z(n10448) );
  XOR U10536 ( .A(n10449), .B(n10448), .Z(n10460) );
  NANDN U10537 ( .A(n10240), .B(n10239), .Z(n10244) );
  NANDN U10538 ( .A(n10242), .B(n10241), .Z(n10243) );
  AND U10539 ( .A(n10244), .B(n10243), .Z(n10458) );
  NANDN U10540 ( .A(n10250), .B(n10249), .Z(n10254) );
  OR U10541 ( .A(n10252), .B(n10251), .Z(n10253) );
  AND U10542 ( .A(n10254), .B(n10253), .Z(n10453) );
  NANDN U10543 ( .A(n10256), .B(n10255), .Z(n10260) );
  NANDN U10544 ( .A(n10258), .B(n10257), .Z(n10259) );
  AND U10545 ( .A(n10260), .B(n10259), .Z(n10393) );
  NANDN U10546 ( .A(n10262), .B(n10261), .Z(n10266) );
  OR U10547 ( .A(n10264), .B(n10263), .Z(n10265) );
  NAND U10548 ( .A(n10266), .B(n10265), .Z(n10392) );
  XNOR U10549 ( .A(n10393), .B(n10392), .Z(n10394) );
  NAND U10550 ( .A(b[0]), .B(a[84]), .Z(n10267) );
  XNOR U10551 ( .A(b[1]), .B(n10267), .Z(n10269) );
  NANDN U10552 ( .A(b[0]), .B(a[83]), .Z(n10268) );
  NAND U10553 ( .A(n10269), .B(n10268), .Z(n10341) );
  NANDN U10554 ( .A(n19394), .B(n10270), .Z(n10272) );
  XOR U10555 ( .A(b[29]), .B(a[56]), .Z(n10419) );
  NANDN U10556 ( .A(n19395), .B(n10419), .Z(n10271) );
  AND U10557 ( .A(n10272), .B(n10271), .Z(n10339) );
  AND U10558 ( .A(b[31]), .B(a[52]), .Z(n10338) );
  XNOR U10559 ( .A(n10339), .B(n10338), .Z(n10340) );
  XNOR U10560 ( .A(n10341), .B(n10340), .Z(n10380) );
  NANDN U10561 ( .A(n19005), .B(n10273), .Z(n10275) );
  XOR U10562 ( .A(b[23]), .B(a[62]), .Z(n10422) );
  NANDN U10563 ( .A(n19055), .B(n10422), .Z(n10274) );
  AND U10564 ( .A(n10275), .B(n10274), .Z(n10413) );
  NANDN U10565 ( .A(n17362), .B(n10276), .Z(n10278) );
  XOR U10566 ( .A(b[7]), .B(a[78]), .Z(n10425) );
  NANDN U10567 ( .A(n17522), .B(n10425), .Z(n10277) );
  AND U10568 ( .A(n10278), .B(n10277), .Z(n10411) );
  NANDN U10569 ( .A(n19116), .B(n10279), .Z(n10281) );
  XOR U10570 ( .A(b[25]), .B(a[60]), .Z(n10428) );
  NANDN U10571 ( .A(n19179), .B(n10428), .Z(n10280) );
  NAND U10572 ( .A(n10281), .B(n10280), .Z(n10410) );
  XNOR U10573 ( .A(n10411), .B(n10410), .Z(n10412) );
  XOR U10574 ( .A(n10413), .B(n10412), .Z(n10381) );
  XNOR U10575 ( .A(n10380), .B(n10381), .Z(n10382) );
  NANDN U10576 ( .A(n18113), .B(n10282), .Z(n10284) );
  XOR U10577 ( .A(b[13]), .B(a[72]), .Z(n10431) );
  NANDN U10578 ( .A(n18229), .B(n10431), .Z(n10283) );
  AND U10579 ( .A(n10284), .B(n10283), .Z(n10375) );
  NANDN U10580 ( .A(n17888), .B(n10285), .Z(n10287) );
  XOR U10581 ( .A(b[11]), .B(a[74]), .Z(n10434) );
  NANDN U10582 ( .A(n18025), .B(n10434), .Z(n10286) );
  NAND U10583 ( .A(n10287), .B(n10286), .Z(n10374) );
  XNOR U10584 ( .A(n10375), .B(n10374), .Z(n10376) );
  NANDN U10585 ( .A(n18487), .B(n10288), .Z(n10290) );
  XOR U10586 ( .A(b[15]), .B(a[70]), .Z(n10437) );
  NANDN U10587 ( .A(n18311), .B(n10437), .Z(n10289) );
  AND U10588 ( .A(n10290), .B(n10289), .Z(n10371) );
  NANDN U10589 ( .A(n18853), .B(n10291), .Z(n10293) );
  XOR U10590 ( .A(b[21]), .B(a[64]), .Z(n10440) );
  NANDN U10591 ( .A(n18926), .B(n10440), .Z(n10292) );
  AND U10592 ( .A(n10293), .B(n10292), .Z(n10369) );
  NANDN U10593 ( .A(n17613), .B(n10294), .Z(n10296) );
  XOR U10594 ( .A(b[9]), .B(a[76]), .Z(n10443) );
  NANDN U10595 ( .A(n17739), .B(n10443), .Z(n10295) );
  NAND U10596 ( .A(n10296), .B(n10295), .Z(n10368) );
  XNOR U10597 ( .A(n10369), .B(n10368), .Z(n10370) );
  XOR U10598 ( .A(n10371), .B(n10370), .Z(n10377) );
  XOR U10599 ( .A(n10376), .B(n10377), .Z(n10383) );
  XOR U10600 ( .A(n10382), .B(n10383), .Z(n10395) );
  XNOR U10601 ( .A(n10394), .B(n10395), .Z(n10452) );
  XNOR U10602 ( .A(n10453), .B(n10452), .Z(n10454) );
  XOR U10603 ( .A(n10455), .B(n10454), .Z(n10459) );
  XOR U10604 ( .A(n10458), .B(n10459), .Z(n10461) );
  XOR U10605 ( .A(n10460), .B(n10461), .Z(n10335) );
  NANDN U10606 ( .A(n10298), .B(n10297), .Z(n10302) );
  NAND U10607 ( .A(n10300), .B(n10299), .Z(n10301) );
  AND U10608 ( .A(n10302), .B(n10301), .Z(n10333) );
  NANDN U10609 ( .A(n10304), .B(n10303), .Z(n10308) );
  NANDN U10610 ( .A(n10306), .B(n10305), .Z(n10307) );
  AND U10611 ( .A(n10308), .B(n10307), .Z(n10332) );
  XNOR U10612 ( .A(n10333), .B(n10332), .Z(n10334) );
  XNOR U10613 ( .A(n10335), .B(n10334), .Z(n10326) );
  NANDN U10614 ( .A(n10310), .B(n10309), .Z(n10314) );
  OR U10615 ( .A(n10312), .B(n10311), .Z(n10313) );
  NAND U10616 ( .A(n10314), .B(n10313), .Z(n10327) );
  XNOR U10617 ( .A(n10326), .B(n10327), .Z(n10328) );
  XNOR U10618 ( .A(n10329), .B(n10328), .Z(n10320) );
  XNOR U10619 ( .A(n10321), .B(n10320), .Z(n10322) );
  XNOR U10620 ( .A(n10323), .B(n10322), .Z(n10464) );
  XNOR U10621 ( .A(sreg[180]), .B(n10464), .Z(n10466) );
  NANDN U10622 ( .A(sreg[179]), .B(n10315), .Z(n10319) );
  NAND U10623 ( .A(n10317), .B(n10316), .Z(n10318) );
  NAND U10624 ( .A(n10319), .B(n10318), .Z(n10465) );
  XNOR U10625 ( .A(n10466), .B(n10465), .Z(c[180]) );
  NANDN U10626 ( .A(n10321), .B(n10320), .Z(n10325) );
  NANDN U10627 ( .A(n10323), .B(n10322), .Z(n10324) );
  AND U10628 ( .A(n10325), .B(n10324), .Z(n10472) );
  NANDN U10629 ( .A(n10327), .B(n10326), .Z(n10331) );
  NANDN U10630 ( .A(n10329), .B(n10328), .Z(n10330) );
  AND U10631 ( .A(n10331), .B(n10330), .Z(n10470) );
  NANDN U10632 ( .A(n10333), .B(n10332), .Z(n10337) );
  NANDN U10633 ( .A(n10335), .B(n10334), .Z(n10336) );
  AND U10634 ( .A(n10337), .B(n10336), .Z(n10478) );
  NANDN U10635 ( .A(n10339), .B(n10338), .Z(n10343) );
  NANDN U10636 ( .A(n10341), .B(n10340), .Z(n10342) );
  AND U10637 ( .A(n10343), .B(n10342), .Z(n10559) );
  NANDN U10638 ( .A(n19237), .B(n10344), .Z(n10346) );
  XOR U10639 ( .A(b[27]), .B(a[59]), .Z(n10505) );
  NANDN U10640 ( .A(n19277), .B(n10505), .Z(n10345) );
  AND U10641 ( .A(n10346), .B(n10345), .Z(n10566) );
  NANDN U10642 ( .A(n17072), .B(n10347), .Z(n10349) );
  XOR U10643 ( .A(b[5]), .B(a[81]), .Z(n10508) );
  NANDN U10644 ( .A(n17223), .B(n10508), .Z(n10348) );
  AND U10645 ( .A(n10349), .B(n10348), .Z(n10564) );
  NANDN U10646 ( .A(n18673), .B(n10350), .Z(n10352) );
  XOR U10647 ( .A(b[19]), .B(a[67]), .Z(n10511) );
  NANDN U10648 ( .A(n18758), .B(n10511), .Z(n10351) );
  NAND U10649 ( .A(n10352), .B(n10351), .Z(n10563) );
  XNOR U10650 ( .A(n10564), .B(n10563), .Z(n10565) );
  XNOR U10651 ( .A(n10566), .B(n10565), .Z(n10557) );
  NANDN U10652 ( .A(n19425), .B(n10353), .Z(n10355) );
  XOR U10653 ( .A(b[31]), .B(a[55]), .Z(n10514) );
  NANDN U10654 ( .A(n19426), .B(n10514), .Z(n10354) );
  AND U10655 ( .A(n10355), .B(n10354), .Z(n10526) );
  NANDN U10656 ( .A(n17067), .B(n10356), .Z(n10358) );
  XOR U10657 ( .A(b[3]), .B(a[83]), .Z(n10517) );
  NANDN U10658 ( .A(n17068), .B(n10517), .Z(n10357) );
  AND U10659 ( .A(n10358), .B(n10357), .Z(n10524) );
  NANDN U10660 ( .A(n18514), .B(n10359), .Z(n10361) );
  XOR U10661 ( .A(b[17]), .B(a[69]), .Z(n10520) );
  NANDN U10662 ( .A(n18585), .B(n10520), .Z(n10360) );
  NAND U10663 ( .A(n10361), .B(n10360), .Z(n10523) );
  XNOR U10664 ( .A(n10524), .B(n10523), .Z(n10525) );
  XOR U10665 ( .A(n10526), .B(n10525), .Z(n10558) );
  XOR U10666 ( .A(n10557), .B(n10558), .Z(n10560) );
  XOR U10667 ( .A(n10559), .B(n10560), .Z(n10494) );
  NANDN U10668 ( .A(n10363), .B(n10362), .Z(n10367) );
  NANDN U10669 ( .A(n10365), .B(n10364), .Z(n10366) );
  AND U10670 ( .A(n10367), .B(n10366), .Z(n10547) );
  NANDN U10671 ( .A(n10369), .B(n10368), .Z(n10373) );
  NANDN U10672 ( .A(n10371), .B(n10370), .Z(n10372) );
  NAND U10673 ( .A(n10373), .B(n10372), .Z(n10548) );
  XNOR U10674 ( .A(n10547), .B(n10548), .Z(n10549) );
  NANDN U10675 ( .A(n10375), .B(n10374), .Z(n10379) );
  NANDN U10676 ( .A(n10377), .B(n10376), .Z(n10378) );
  NAND U10677 ( .A(n10379), .B(n10378), .Z(n10550) );
  XNOR U10678 ( .A(n10549), .B(n10550), .Z(n10493) );
  XNOR U10679 ( .A(n10494), .B(n10493), .Z(n10496) );
  NANDN U10680 ( .A(n10381), .B(n10380), .Z(n10385) );
  NANDN U10681 ( .A(n10383), .B(n10382), .Z(n10384) );
  AND U10682 ( .A(n10385), .B(n10384), .Z(n10495) );
  XOR U10683 ( .A(n10496), .B(n10495), .Z(n10607) );
  NANDN U10684 ( .A(n10387), .B(n10386), .Z(n10391) );
  NANDN U10685 ( .A(n10389), .B(n10388), .Z(n10390) );
  AND U10686 ( .A(n10391), .B(n10390), .Z(n10605) );
  NANDN U10687 ( .A(n10393), .B(n10392), .Z(n10397) );
  NANDN U10688 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U10689 ( .A(n10397), .B(n10396), .Z(n10490) );
  NANDN U10690 ( .A(n10399), .B(n10398), .Z(n10403) );
  OR U10691 ( .A(n10401), .B(n10400), .Z(n10402) );
  AND U10692 ( .A(n10403), .B(n10402), .Z(n10488) );
  NANDN U10693 ( .A(n10405), .B(n10404), .Z(n10409) );
  NANDN U10694 ( .A(n10407), .B(n10406), .Z(n10408) );
  AND U10695 ( .A(n10409), .B(n10408), .Z(n10554) );
  NANDN U10696 ( .A(n10411), .B(n10410), .Z(n10415) );
  NANDN U10697 ( .A(n10413), .B(n10412), .Z(n10414) );
  NAND U10698 ( .A(n10415), .B(n10414), .Z(n10553) );
  XNOR U10699 ( .A(n10554), .B(n10553), .Z(n10556) );
  NAND U10700 ( .A(b[0]), .B(a[85]), .Z(n10416) );
  XNOR U10701 ( .A(b[1]), .B(n10416), .Z(n10418) );
  NANDN U10702 ( .A(b[0]), .B(a[84]), .Z(n10417) );
  NAND U10703 ( .A(n10418), .B(n10417), .Z(n10502) );
  NANDN U10704 ( .A(n19394), .B(n10419), .Z(n10421) );
  XOR U10705 ( .A(b[29]), .B(a[57]), .Z(n10578) );
  NANDN U10706 ( .A(n19395), .B(n10578), .Z(n10420) );
  AND U10707 ( .A(n10421), .B(n10420), .Z(n10500) );
  AND U10708 ( .A(b[31]), .B(a[53]), .Z(n10499) );
  XNOR U10709 ( .A(n10500), .B(n10499), .Z(n10501) );
  XNOR U10710 ( .A(n10502), .B(n10501), .Z(n10542) );
  NANDN U10711 ( .A(n19005), .B(n10422), .Z(n10424) );
  XOR U10712 ( .A(b[23]), .B(a[63]), .Z(n10581) );
  NANDN U10713 ( .A(n19055), .B(n10581), .Z(n10423) );
  AND U10714 ( .A(n10424), .B(n10423), .Z(n10571) );
  NANDN U10715 ( .A(n17362), .B(n10425), .Z(n10427) );
  XOR U10716 ( .A(b[7]), .B(a[79]), .Z(n10584) );
  NANDN U10717 ( .A(n17522), .B(n10584), .Z(n10426) );
  AND U10718 ( .A(n10427), .B(n10426), .Z(n10570) );
  NANDN U10719 ( .A(n19116), .B(n10428), .Z(n10430) );
  XOR U10720 ( .A(b[25]), .B(a[61]), .Z(n10587) );
  NANDN U10721 ( .A(n19179), .B(n10587), .Z(n10429) );
  NAND U10722 ( .A(n10430), .B(n10429), .Z(n10569) );
  XOR U10723 ( .A(n10570), .B(n10569), .Z(n10572) );
  XOR U10724 ( .A(n10571), .B(n10572), .Z(n10541) );
  XOR U10725 ( .A(n10542), .B(n10541), .Z(n10544) );
  NANDN U10726 ( .A(n18113), .B(n10431), .Z(n10433) );
  XOR U10727 ( .A(b[13]), .B(a[73]), .Z(n10590) );
  NANDN U10728 ( .A(n18229), .B(n10590), .Z(n10432) );
  AND U10729 ( .A(n10433), .B(n10432), .Z(n10536) );
  NANDN U10730 ( .A(n17888), .B(n10434), .Z(n10436) );
  XOR U10731 ( .A(b[11]), .B(a[75]), .Z(n10593) );
  NANDN U10732 ( .A(n18025), .B(n10593), .Z(n10435) );
  NAND U10733 ( .A(n10436), .B(n10435), .Z(n10535) );
  XNOR U10734 ( .A(n10536), .B(n10535), .Z(n10538) );
  NANDN U10735 ( .A(n18487), .B(n10437), .Z(n10439) );
  XOR U10736 ( .A(b[15]), .B(a[71]), .Z(n10596) );
  NANDN U10737 ( .A(n18311), .B(n10596), .Z(n10438) );
  AND U10738 ( .A(n10439), .B(n10438), .Z(n10532) );
  NANDN U10739 ( .A(n18853), .B(n10440), .Z(n10442) );
  XOR U10740 ( .A(b[21]), .B(a[65]), .Z(n10599) );
  NANDN U10741 ( .A(n18926), .B(n10599), .Z(n10441) );
  AND U10742 ( .A(n10442), .B(n10441), .Z(n10530) );
  NANDN U10743 ( .A(n17613), .B(n10443), .Z(n10445) );
  XOR U10744 ( .A(b[9]), .B(a[77]), .Z(n10602) );
  NANDN U10745 ( .A(n17739), .B(n10602), .Z(n10444) );
  NAND U10746 ( .A(n10445), .B(n10444), .Z(n10529) );
  XNOR U10747 ( .A(n10530), .B(n10529), .Z(n10531) );
  XNOR U10748 ( .A(n10532), .B(n10531), .Z(n10537) );
  XOR U10749 ( .A(n10538), .B(n10537), .Z(n10543) );
  XOR U10750 ( .A(n10544), .B(n10543), .Z(n10555) );
  XOR U10751 ( .A(n10556), .B(n10555), .Z(n10487) );
  XNOR U10752 ( .A(n10488), .B(n10487), .Z(n10489) );
  XOR U10753 ( .A(n10490), .B(n10489), .Z(n10606) );
  XOR U10754 ( .A(n10605), .B(n10606), .Z(n10608) );
  XOR U10755 ( .A(n10607), .B(n10608), .Z(n10484) );
  NANDN U10756 ( .A(n10447), .B(n10446), .Z(n10451) );
  NAND U10757 ( .A(n10449), .B(n10448), .Z(n10450) );
  AND U10758 ( .A(n10451), .B(n10450), .Z(n10482) );
  NANDN U10759 ( .A(n10453), .B(n10452), .Z(n10457) );
  NANDN U10760 ( .A(n10455), .B(n10454), .Z(n10456) );
  AND U10761 ( .A(n10457), .B(n10456), .Z(n10481) );
  XNOR U10762 ( .A(n10482), .B(n10481), .Z(n10483) );
  XNOR U10763 ( .A(n10484), .B(n10483), .Z(n10475) );
  NANDN U10764 ( .A(n10459), .B(n10458), .Z(n10463) );
  OR U10765 ( .A(n10461), .B(n10460), .Z(n10462) );
  NAND U10766 ( .A(n10463), .B(n10462), .Z(n10476) );
  XNOR U10767 ( .A(n10475), .B(n10476), .Z(n10477) );
  XNOR U10768 ( .A(n10478), .B(n10477), .Z(n10469) );
  XNOR U10769 ( .A(n10470), .B(n10469), .Z(n10471) );
  XNOR U10770 ( .A(n10472), .B(n10471), .Z(n10611) );
  XNOR U10771 ( .A(sreg[181]), .B(n10611), .Z(n10613) );
  NANDN U10772 ( .A(sreg[180]), .B(n10464), .Z(n10468) );
  NAND U10773 ( .A(n10466), .B(n10465), .Z(n10467) );
  NAND U10774 ( .A(n10468), .B(n10467), .Z(n10612) );
  XNOR U10775 ( .A(n10613), .B(n10612), .Z(c[181]) );
  NANDN U10776 ( .A(n10470), .B(n10469), .Z(n10474) );
  NANDN U10777 ( .A(n10472), .B(n10471), .Z(n10473) );
  AND U10778 ( .A(n10474), .B(n10473), .Z(n10619) );
  NANDN U10779 ( .A(n10476), .B(n10475), .Z(n10480) );
  NANDN U10780 ( .A(n10478), .B(n10477), .Z(n10479) );
  AND U10781 ( .A(n10480), .B(n10479), .Z(n10617) );
  NANDN U10782 ( .A(n10482), .B(n10481), .Z(n10486) );
  NANDN U10783 ( .A(n10484), .B(n10483), .Z(n10485) );
  AND U10784 ( .A(n10486), .B(n10485), .Z(n10625) );
  NANDN U10785 ( .A(n10488), .B(n10487), .Z(n10492) );
  NANDN U10786 ( .A(n10490), .B(n10489), .Z(n10491) );
  AND U10787 ( .A(n10492), .B(n10491), .Z(n10629) );
  NANDN U10788 ( .A(n10494), .B(n10493), .Z(n10498) );
  NAND U10789 ( .A(n10496), .B(n10495), .Z(n10497) );
  AND U10790 ( .A(n10498), .B(n10497), .Z(n10628) );
  XNOR U10791 ( .A(n10629), .B(n10628), .Z(n10631) );
  NANDN U10792 ( .A(n10500), .B(n10499), .Z(n10504) );
  NANDN U10793 ( .A(n10502), .B(n10501), .Z(n10503) );
  AND U10794 ( .A(n10504), .B(n10503), .Z(n10696) );
  NANDN U10795 ( .A(n19237), .B(n10505), .Z(n10507) );
  XOR U10796 ( .A(b[27]), .B(a[60]), .Z(n10640) );
  NANDN U10797 ( .A(n19277), .B(n10640), .Z(n10506) );
  AND U10798 ( .A(n10507), .B(n10506), .Z(n10703) );
  NANDN U10799 ( .A(n17072), .B(n10508), .Z(n10510) );
  XOR U10800 ( .A(b[5]), .B(a[82]), .Z(n10643) );
  NANDN U10801 ( .A(n17223), .B(n10643), .Z(n10509) );
  AND U10802 ( .A(n10510), .B(n10509), .Z(n10701) );
  NANDN U10803 ( .A(n18673), .B(n10511), .Z(n10513) );
  XOR U10804 ( .A(b[19]), .B(a[68]), .Z(n10646) );
  NANDN U10805 ( .A(n18758), .B(n10646), .Z(n10512) );
  NAND U10806 ( .A(n10513), .B(n10512), .Z(n10700) );
  XNOR U10807 ( .A(n10701), .B(n10700), .Z(n10702) );
  XNOR U10808 ( .A(n10703), .B(n10702), .Z(n10694) );
  NANDN U10809 ( .A(n19425), .B(n10514), .Z(n10516) );
  XOR U10810 ( .A(b[31]), .B(a[56]), .Z(n10649) );
  NANDN U10811 ( .A(n19426), .B(n10649), .Z(n10515) );
  AND U10812 ( .A(n10516), .B(n10515), .Z(n10661) );
  NANDN U10813 ( .A(n17067), .B(n10517), .Z(n10519) );
  XOR U10814 ( .A(b[3]), .B(a[84]), .Z(n10652) );
  NANDN U10815 ( .A(n17068), .B(n10652), .Z(n10518) );
  AND U10816 ( .A(n10519), .B(n10518), .Z(n10659) );
  NANDN U10817 ( .A(n18514), .B(n10520), .Z(n10522) );
  XOR U10818 ( .A(b[17]), .B(a[70]), .Z(n10655) );
  NANDN U10819 ( .A(n18585), .B(n10655), .Z(n10521) );
  NAND U10820 ( .A(n10522), .B(n10521), .Z(n10658) );
  XNOR U10821 ( .A(n10659), .B(n10658), .Z(n10660) );
  XOR U10822 ( .A(n10661), .B(n10660), .Z(n10695) );
  XOR U10823 ( .A(n10694), .B(n10695), .Z(n10697) );
  XOR U10824 ( .A(n10696), .B(n10697), .Z(n10743) );
  NANDN U10825 ( .A(n10524), .B(n10523), .Z(n10528) );
  NANDN U10826 ( .A(n10526), .B(n10525), .Z(n10527) );
  AND U10827 ( .A(n10528), .B(n10527), .Z(n10682) );
  NANDN U10828 ( .A(n10530), .B(n10529), .Z(n10534) );
  NANDN U10829 ( .A(n10532), .B(n10531), .Z(n10533) );
  NAND U10830 ( .A(n10534), .B(n10533), .Z(n10683) );
  XNOR U10831 ( .A(n10682), .B(n10683), .Z(n10684) );
  NANDN U10832 ( .A(n10536), .B(n10535), .Z(n10540) );
  NAND U10833 ( .A(n10538), .B(n10537), .Z(n10539) );
  NAND U10834 ( .A(n10540), .B(n10539), .Z(n10685) );
  XNOR U10835 ( .A(n10684), .B(n10685), .Z(n10742) );
  XNOR U10836 ( .A(n10743), .B(n10742), .Z(n10745) );
  NAND U10837 ( .A(n10542), .B(n10541), .Z(n10546) );
  NAND U10838 ( .A(n10544), .B(n10543), .Z(n10545) );
  AND U10839 ( .A(n10546), .B(n10545), .Z(n10744) );
  XOR U10840 ( .A(n10745), .B(n10744), .Z(n10757) );
  NANDN U10841 ( .A(n10548), .B(n10547), .Z(n10552) );
  NANDN U10842 ( .A(n10550), .B(n10549), .Z(n10551) );
  AND U10843 ( .A(n10552), .B(n10551), .Z(n10754) );
  NANDN U10844 ( .A(n10558), .B(n10557), .Z(n10562) );
  OR U10845 ( .A(n10560), .B(n10559), .Z(n10561) );
  AND U10846 ( .A(n10562), .B(n10561), .Z(n10749) );
  NANDN U10847 ( .A(n10564), .B(n10563), .Z(n10568) );
  NANDN U10848 ( .A(n10566), .B(n10565), .Z(n10567) );
  AND U10849 ( .A(n10568), .B(n10567), .Z(n10689) );
  NANDN U10850 ( .A(n10570), .B(n10569), .Z(n10574) );
  OR U10851 ( .A(n10572), .B(n10571), .Z(n10573) );
  NAND U10852 ( .A(n10574), .B(n10573), .Z(n10688) );
  XNOR U10853 ( .A(n10689), .B(n10688), .Z(n10690) );
  NAND U10854 ( .A(b[0]), .B(a[86]), .Z(n10575) );
  XNOR U10855 ( .A(b[1]), .B(n10575), .Z(n10577) );
  NANDN U10856 ( .A(b[0]), .B(a[85]), .Z(n10576) );
  NAND U10857 ( .A(n10577), .B(n10576), .Z(n10637) );
  NANDN U10858 ( .A(n19394), .B(n10578), .Z(n10580) );
  XOR U10859 ( .A(b[29]), .B(a[58]), .Z(n10715) );
  NANDN U10860 ( .A(n19395), .B(n10715), .Z(n10579) );
  AND U10861 ( .A(n10580), .B(n10579), .Z(n10635) );
  AND U10862 ( .A(b[31]), .B(a[54]), .Z(n10634) );
  XNOR U10863 ( .A(n10635), .B(n10634), .Z(n10636) );
  XNOR U10864 ( .A(n10637), .B(n10636), .Z(n10676) );
  NANDN U10865 ( .A(n19005), .B(n10581), .Z(n10583) );
  XOR U10866 ( .A(b[23]), .B(a[64]), .Z(n10718) );
  NANDN U10867 ( .A(n19055), .B(n10718), .Z(n10582) );
  AND U10868 ( .A(n10583), .B(n10582), .Z(n10709) );
  NANDN U10869 ( .A(n17362), .B(n10584), .Z(n10586) );
  XOR U10870 ( .A(b[7]), .B(a[80]), .Z(n10721) );
  NANDN U10871 ( .A(n17522), .B(n10721), .Z(n10585) );
  AND U10872 ( .A(n10586), .B(n10585), .Z(n10707) );
  NANDN U10873 ( .A(n19116), .B(n10587), .Z(n10589) );
  XOR U10874 ( .A(b[25]), .B(a[62]), .Z(n10724) );
  NANDN U10875 ( .A(n19179), .B(n10724), .Z(n10588) );
  NAND U10876 ( .A(n10589), .B(n10588), .Z(n10706) );
  XNOR U10877 ( .A(n10707), .B(n10706), .Z(n10708) );
  XOR U10878 ( .A(n10709), .B(n10708), .Z(n10677) );
  XNOR U10879 ( .A(n10676), .B(n10677), .Z(n10678) );
  NANDN U10880 ( .A(n18113), .B(n10590), .Z(n10592) );
  XOR U10881 ( .A(b[13]), .B(a[74]), .Z(n10727) );
  NANDN U10882 ( .A(n18229), .B(n10727), .Z(n10591) );
  AND U10883 ( .A(n10592), .B(n10591), .Z(n10671) );
  NANDN U10884 ( .A(n17888), .B(n10593), .Z(n10595) );
  XOR U10885 ( .A(b[11]), .B(a[76]), .Z(n10730) );
  NANDN U10886 ( .A(n18025), .B(n10730), .Z(n10594) );
  NAND U10887 ( .A(n10595), .B(n10594), .Z(n10670) );
  XNOR U10888 ( .A(n10671), .B(n10670), .Z(n10672) );
  NANDN U10889 ( .A(n18487), .B(n10596), .Z(n10598) );
  XOR U10890 ( .A(b[15]), .B(a[72]), .Z(n10733) );
  NANDN U10891 ( .A(n18311), .B(n10733), .Z(n10597) );
  AND U10892 ( .A(n10598), .B(n10597), .Z(n10667) );
  NANDN U10893 ( .A(n18853), .B(n10599), .Z(n10601) );
  XOR U10894 ( .A(b[21]), .B(a[66]), .Z(n10736) );
  NANDN U10895 ( .A(n18926), .B(n10736), .Z(n10600) );
  AND U10896 ( .A(n10601), .B(n10600), .Z(n10665) );
  NANDN U10897 ( .A(n17613), .B(n10602), .Z(n10604) );
  XOR U10898 ( .A(b[9]), .B(a[78]), .Z(n10739) );
  NANDN U10899 ( .A(n17739), .B(n10739), .Z(n10603) );
  NAND U10900 ( .A(n10604), .B(n10603), .Z(n10664) );
  XNOR U10901 ( .A(n10665), .B(n10664), .Z(n10666) );
  XOR U10902 ( .A(n10667), .B(n10666), .Z(n10673) );
  XOR U10903 ( .A(n10672), .B(n10673), .Z(n10679) );
  XOR U10904 ( .A(n10678), .B(n10679), .Z(n10691) );
  XNOR U10905 ( .A(n10690), .B(n10691), .Z(n10748) );
  XNOR U10906 ( .A(n10749), .B(n10748), .Z(n10750) );
  XOR U10907 ( .A(n10751), .B(n10750), .Z(n10755) );
  XNOR U10908 ( .A(n10754), .B(n10755), .Z(n10756) );
  XNOR U10909 ( .A(n10757), .B(n10756), .Z(n10630) );
  XOR U10910 ( .A(n10631), .B(n10630), .Z(n10623) );
  NANDN U10911 ( .A(n10606), .B(n10605), .Z(n10610) );
  OR U10912 ( .A(n10608), .B(n10607), .Z(n10609) );
  AND U10913 ( .A(n10610), .B(n10609), .Z(n10622) );
  XNOR U10914 ( .A(n10623), .B(n10622), .Z(n10624) );
  XNOR U10915 ( .A(n10625), .B(n10624), .Z(n10616) );
  XNOR U10916 ( .A(n10617), .B(n10616), .Z(n10618) );
  XNOR U10917 ( .A(n10619), .B(n10618), .Z(n10760) );
  XNOR U10918 ( .A(sreg[182]), .B(n10760), .Z(n10762) );
  NANDN U10919 ( .A(sreg[181]), .B(n10611), .Z(n10615) );
  NAND U10920 ( .A(n10613), .B(n10612), .Z(n10614) );
  NAND U10921 ( .A(n10615), .B(n10614), .Z(n10761) );
  XNOR U10922 ( .A(n10762), .B(n10761), .Z(c[182]) );
  NANDN U10923 ( .A(n10617), .B(n10616), .Z(n10621) );
  NANDN U10924 ( .A(n10619), .B(n10618), .Z(n10620) );
  AND U10925 ( .A(n10621), .B(n10620), .Z(n10768) );
  NANDN U10926 ( .A(n10623), .B(n10622), .Z(n10627) );
  NANDN U10927 ( .A(n10625), .B(n10624), .Z(n10626) );
  AND U10928 ( .A(n10627), .B(n10626), .Z(n10766) );
  NANDN U10929 ( .A(n10629), .B(n10628), .Z(n10633) );
  NAND U10930 ( .A(n10631), .B(n10630), .Z(n10632) );
  AND U10931 ( .A(n10633), .B(n10632), .Z(n10773) );
  NANDN U10932 ( .A(n10635), .B(n10634), .Z(n10639) );
  NANDN U10933 ( .A(n10637), .B(n10636), .Z(n10638) );
  AND U10934 ( .A(n10639), .B(n10638), .Z(n10857) );
  NANDN U10935 ( .A(n19237), .B(n10640), .Z(n10642) );
  XOR U10936 ( .A(b[27]), .B(a[61]), .Z(n10801) );
  NANDN U10937 ( .A(n19277), .B(n10801), .Z(n10641) );
  AND U10938 ( .A(n10642), .B(n10641), .Z(n10864) );
  NANDN U10939 ( .A(n17072), .B(n10643), .Z(n10645) );
  XOR U10940 ( .A(b[5]), .B(a[83]), .Z(n10804) );
  NANDN U10941 ( .A(n17223), .B(n10804), .Z(n10644) );
  AND U10942 ( .A(n10645), .B(n10644), .Z(n10862) );
  NANDN U10943 ( .A(n18673), .B(n10646), .Z(n10648) );
  XOR U10944 ( .A(b[19]), .B(a[69]), .Z(n10807) );
  NANDN U10945 ( .A(n18758), .B(n10807), .Z(n10647) );
  NAND U10946 ( .A(n10648), .B(n10647), .Z(n10861) );
  XNOR U10947 ( .A(n10862), .B(n10861), .Z(n10863) );
  XNOR U10948 ( .A(n10864), .B(n10863), .Z(n10855) );
  NANDN U10949 ( .A(n19425), .B(n10649), .Z(n10651) );
  XOR U10950 ( .A(b[31]), .B(a[57]), .Z(n10810) );
  NANDN U10951 ( .A(n19426), .B(n10810), .Z(n10650) );
  AND U10952 ( .A(n10651), .B(n10650), .Z(n10822) );
  NANDN U10953 ( .A(n17067), .B(n10652), .Z(n10654) );
  XOR U10954 ( .A(b[3]), .B(a[85]), .Z(n10813) );
  NANDN U10955 ( .A(n17068), .B(n10813), .Z(n10653) );
  AND U10956 ( .A(n10654), .B(n10653), .Z(n10820) );
  NANDN U10957 ( .A(n18514), .B(n10655), .Z(n10657) );
  XOR U10958 ( .A(b[17]), .B(a[71]), .Z(n10816) );
  NANDN U10959 ( .A(n18585), .B(n10816), .Z(n10656) );
  NAND U10960 ( .A(n10657), .B(n10656), .Z(n10819) );
  XNOR U10961 ( .A(n10820), .B(n10819), .Z(n10821) );
  XOR U10962 ( .A(n10822), .B(n10821), .Z(n10856) );
  XOR U10963 ( .A(n10855), .B(n10856), .Z(n10858) );
  XOR U10964 ( .A(n10857), .B(n10858), .Z(n10790) );
  NANDN U10965 ( .A(n10659), .B(n10658), .Z(n10663) );
  NANDN U10966 ( .A(n10661), .B(n10660), .Z(n10662) );
  AND U10967 ( .A(n10663), .B(n10662), .Z(n10843) );
  NANDN U10968 ( .A(n10665), .B(n10664), .Z(n10669) );
  NANDN U10969 ( .A(n10667), .B(n10666), .Z(n10668) );
  NAND U10970 ( .A(n10669), .B(n10668), .Z(n10844) );
  XNOR U10971 ( .A(n10843), .B(n10844), .Z(n10845) );
  NANDN U10972 ( .A(n10671), .B(n10670), .Z(n10675) );
  NANDN U10973 ( .A(n10673), .B(n10672), .Z(n10674) );
  NAND U10974 ( .A(n10675), .B(n10674), .Z(n10846) );
  XNOR U10975 ( .A(n10845), .B(n10846), .Z(n10789) );
  XNOR U10976 ( .A(n10790), .B(n10789), .Z(n10792) );
  NANDN U10977 ( .A(n10677), .B(n10676), .Z(n10681) );
  NANDN U10978 ( .A(n10679), .B(n10678), .Z(n10680) );
  AND U10979 ( .A(n10681), .B(n10680), .Z(n10791) );
  XOR U10980 ( .A(n10792), .B(n10791), .Z(n10905) );
  NANDN U10981 ( .A(n10683), .B(n10682), .Z(n10687) );
  NANDN U10982 ( .A(n10685), .B(n10684), .Z(n10686) );
  AND U10983 ( .A(n10687), .B(n10686), .Z(n10903) );
  NANDN U10984 ( .A(n10689), .B(n10688), .Z(n10693) );
  NANDN U10985 ( .A(n10691), .B(n10690), .Z(n10692) );
  AND U10986 ( .A(n10693), .B(n10692), .Z(n10786) );
  NANDN U10987 ( .A(n10695), .B(n10694), .Z(n10699) );
  OR U10988 ( .A(n10697), .B(n10696), .Z(n10698) );
  AND U10989 ( .A(n10699), .B(n10698), .Z(n10784) );
  NANDN U10990 ( .A(n10701), .B(n10700), .Z(n10705) );
  NANDN U10991 ( .A(n10703), .B(n10702), .Z(n10704) );
  AND U10992 ( .A(n10705), .B(n10704), .Z(n10850) );
  NANDN U10993 ( .A(n10707), .B(n10706), .Z(n10711) );
  NANDN U10994 ( .A(n10709), .B(n10708), .Z(n10710) );
  NAND U10995 ( .A(n10711), .B(n10710), .Z(n10849) );
  XNOR U10996 ( .A(n10850), .B(n10849), .Z(n10851) );
  NAND U10997 ( .A(b[0]), .B(a[87]), .Z(n10712) );
  XNOR U10998 ( .A(b[1]), .B(n10712), .Z(n10714) );
  NANDN U10999 ( .A(b[0]), .B(a[86]), .Z(n10713) );
  NAND U11000 ( .A(n10714), .B(n10713), .Z(n10798) );
  NANDN U11001 ( .A(n19394), .B(n10715), .Z(n10717) );
  XOR U11002 ( .A(b[29]), .B(a[59]), .Z(n10876) );
  NANDN U11003 ( .A(n19395), .B(n10876), .Z(n10716) );
  AND U11004 ( .A(n10717), .B(n10716), .Z(n10796) );
  AND U11005 ( .A(b[31]), .B(a[55]), .Z(n10795) );
  XNOR U11006 ( .A(n10796), .B(n10795), .Z(n10797) );
  XNOR U11007 ( .A(n10798), .B(n10797), .Z(n10837) );
  NANDN U11008 ( .A(n19005), .B(n10718), .Z(n10720) );
  XOR U11009 ( .A(b[23]), .B(a[65]), .Z(n10879) );
  NANDN U11010 ( .A(n19055), .B(n10879), .Z(n10719) );
  AND U11011 ( .A(n10720), .B(n10719), .Z(n10870) );
  NANDN U11012 ( .A(n17362), .B(n10721), .Z(n10723) );
  XOR U11013 ( .A(b[7]), .B(a[81]), .Z(n10882) );
  NANDN U11014 ( .A(n17522), .B(n10882), .Z(n10722) );
  AND U11015 ( .A(n10723), .B(n10722), .Z(n10868) );
  NANDN U11016 ( .A(n19116), .B(n10724), .Z(n10726) );
  XOR U11017 ( .A(b[25]), .B(a[63]), .Z(n10885) );
  NANDN U11018 ( .A(n19179), .B(n10885), .Z(n10725) );
  NAND U11019 ( .A(n10726), .B(n10725), .Z(n10867) );
  XNOR U11020 ( .A(n10868), .B(n10867), .Z(n10869) );
  XOR U11021 ( .A(n10870), .B(n10869), .Z(n10838) );
  XNOR U11022 ( .A(n10837), .B(n10838), .Z(n10839) );
  NANDN U11023 ( .A(n18113), .B(n10727), .Z(n10729) );
  XOR U11024 ( .A(b[13]), .B(a[75]), .Z(n10888) );
  NANDN U11025 ( .A(n18229), .B(n10888), .Z(n10728) );
  AND U11026 ( .A(n10729), .B(n10728), .Z(n10832) );
  NANDN U11027 ( .A(n17888), .B(n10730), .Z(n10732) );
  XOR U11028 ( .A(b[11]), .B(a[77]), .Z(n10891) );
  NANDN U11029 ( .A(n18025), .B(n10891), .Z(n10731) );
  NAND U11030 ( .A(n10732), .B(n10731), .Z(n10831) );
  XNOR U11031 ( .A(n10832), .B(n10831), .Z(n10833) );
  NANDN U11032 ( .A(n18487), .B(n10733), .Z(n10735) );
  XOR U11033 ( .A(b[15]), .B(a[73]), .Z(n10894) );
  NANDN U11034 ( .A(n18311), .B(n10894), .Z(n10734) );
  AND U11035 ( .A(n10735), .B(n10734), .Z(n10828) );
  NANDN U11036 ( .A(n18853), .B(n10736), .Z(n10738) );
  XOR U11037 ( .A(b[21]), .B(a[67]), .Z(n10897) );
  NANDN U11038 ( .A(n18926), .B(n10897), .Z(n10737) );
  AND U11039 ( .A(n10738), .B(n10737), .Z(n10826) );
  NANDN U11040 ( .A(n17613), .B(n10739), .Z(n10741) );
  XOR U11041 ( .A(b[9]), .B(a[79]), .Z(n10900) );
  NANDN U11042 ( .A(n17739), .B(n10900), .Z(n10740) );
  NAND U11043 ( .A(n10741), .B(n10740), .Z(n10825) );
  XNOR U11044 ( .A(n10826), .B(n10825), .Z(n10827) );
  XOR U11045 ( .A(n10828), .B(n10827), .Z(n10834) );
  XOR U11046 ( .A(n10833), .B(n10834), .Z(n10840) );
  XOR U11047 ( .A(n10839), .B(n10840), .Z(n10852) );
  XNOR U11048 ( .A(n10851), .B(n10852), .Z(n10783) );
  XNOR U11049 ( .A(n10784), .B(n10783), .Z(n10785) );
  XOR U11050 ( .A(n10786), .B(n10785), .Z(n10904) );
  XOR U11051 ( .A(n10903), .B(n10904), .Z(n10906) );
  XOR U11052 ( .A(n10905), .B(n10906), .Z(n10780) );
  NANDN U11053 ( .A(n10743), .B(n10742), .Z(n10747) );
  NAND U11054 ( .A(n10745), .B(n10744), .Z(n10746) );
  AND U11055 ( .A(n10747), .B(n10746), .Z(n10778) );
  NANDN U11056 ( .A(n10749), .B(n10748), .Z(n10753) );
  NANDN U11057 ( .A(n10751), .B(n10750), .Z(n10752) );
  AND U11058 ( .A(n10753), .B(n10752), .Z(n10777) );
  XNOR U11059 ( .A(n10778), .B(n10777), .Z(n10779) );
  XNOR U11060 ( .A(n10780), .B(n10779), .Z(n10771) );
  NANDN U11061 ( .A(n10755), .B(n10754), .Z(n10759) );
  NANDN U11062 ( .A(n10757), .B(n10756), .Z(n10758) );
  NAND U11063 ( .A(n10759), .B(n10758), .Z(n10772) );
  XOR U11064 ( .A(n10771), .B(n10772), .Z(n10774) );
  XNOR U11065 ( .A(n10773), .B(n10774), .Z(n10765) );
  XNOR U11066 ( .A(n10766), .B(n10765), .Z(n10767) );
  XNOR U11067 ( .A(n10768), .B(n10767), .Z(n10909) );
  XNOR U11068 ( .A(sreg[183]), .B(n10909), .Z(n10911) );
  NANDN U11069 ( .A(sreg[182]), .B(n10760), .Z(n10764) );
  NAND U11070 ( .A(n10762), .B(n10761), .Z(n10763) );
  NAND U11071 ( .A(n10764), .B(n10763), .Z(n10910) );
  XNOR U11072 ( .A(n10911), .B(n10910), .Z(c[183]) );
  NANDN U11073 ( .A(n10766), .B(n10765), .Z(n10770) );
  NANDN U11074 ( .A(n10768), .B(n10767), .Z(n10769) );
  AND U11075 ( .A(n10770), .B(n10769), .Z(n10917) );
  NANDN U11076 ( .A(n10772), .B(n10771), .Z(n10776) );
  NANDN U11077 ( .A(n10774), .B(n10773), .Z(n10775) );
  AND U11078 ( .A(n10776), .B(n10775), .Z(n10915) );
  NANDN U11079 ( .A(n10778), .B(n10777), .Z(n10782) );
  NANDN U11080 ( .A(n10780), .B(n10779), .Z(n10781) );
  AND U11081 ( .A(n10782), .B(n10781), .Z(n10923) );
  NANDN U11082 ( .A(n10784), .B(n10783), .Z(n10788) );
  NANDN U11083 ( .A(n10786), .B(n10785), .Z(n10787) );
  AND U11084 ( .A(n10788), .B(n10787), .Z(n10927) );
  NANDN U11085 ( .A(n10790), .B(n10789), .Z(n10794) );
  NAND U11086 ( .A(n10792), .B(n10791), .Z(n10793) );
  AND U11087 ( .A(n10794), .B(n10793), .Z(n10926) );
  XNOR U11088 ( .A(n10927), .B(n10926), .Z(n10929) );
  NANDN U11089 ( .A(n10796), .B(n10795), .Z(n10800) );
  NANDN U11090 ( .A(n10798), .B(n10797), .Z(n10799) );
  AND U11091 ( .A(n10800), .B(n10799), .Z(n11006) );
  NANDN U11092 ( .A(n19237), .B(n10801), .Z(n10803) );
  XOR U11093 ( .A(b[27]), .B(a[62]), .Z(n10950) );
  NANDN U11094 ( .A(n19277), .B(n10950), .Z(n10802) );
  AND U11095 ( .A(n10803), .B(n10802), .Z(n11013) );
  NANDN U11096 ( .A(n17072), .B(n10804), .Z(n10806) );
  XOR U11097 ( .A(b[5]), .B(a[84]), .Z(n10953) );
  NANDN U11098 ( .A(n17223), .B(n10953), .Z(n10805) );
  AND U11099 ( .A(n10806), .B(n10805), .Z(n11011) );
  NANDN U11100 ( .A(n18673), .B(n10807), .Z(n10809) );
  XOR U11101 ( .A(b[19]), .B(a[70]), .Z(n10956) );
  NANDN U11102 ( .A(n18758), .B(n10956), .Z(n10808) );
  NAND U11103 ( .A(n10809), .B(n10808), .Z(n11010) );
  XNOR U11104 ( .A(n11011), .B(n11010), .Z(n11012) );
  XNOR U11105 ( .A(n11013), .B(n11012), .Z(n11004) );
  NANDN U11106 ( .A(n19425), .B(n10810), .Z(n10812) );
  XOR U11107 ( .A(b[31]), .B(a[58]), .Z(n10959) );
  NANDN U11108 ( .A(n19426), .B(n10959), .Z(n10811) );
  AND U11109 ( .A(n10812), .B(n10811), .Z(n10971) );
  NANDN U11110 ( .A(n17067), .B(n10813), .Z(n10815) );
  XOR U11111 ( .A(b[3]), .B(a[86]), .Z(n10962) );
  NANDN U11112 ( .A(n17068), .B(n10962), .Z(n10814) );
  AND U11113 ( .A(n10815), .B(n10814), .Z(n10969) );
  NANDN U11114 ( .A(n18514), .B(n10816), .Z(n10818) );
  XOR U11115 ( .A(b[17]), .B(a[72]), .Z(n10965) );
  NANDN U11116 ( .A(n18585), .B(n10965), .Z(n10817) );
  NAND U11117 ( .A(n10818), .B(n10817), .Z(n10968) );
  XNOR U11118 ( .A(n10969), .B(n10968), .Z(n10970) );
  XOR U11119 ( .A(n10971), .B(n10970), .Z(n11005) );
  XOR U11120 ( .A(n11004), .B(n11005), .Z(n11007) );
  XOR U11121 ( .A(n11006), .B(n11007), .Z(n10939) );
  NANDN U11122 ( .A(n10820), .B(n10819), .Z(n10824) );
  NANDN U11123 ( .A(n10822), .B(n10821), .Z(n10823) );
  AND U11124 ( .A(n10824), .B(n10823), .Z(n10992) );
  NANDN U11125 ( .A(n10826), .B(n10825), .Z(n10830) );
  NANDN U11126 ( .A(n10828), .B(n10827), .Z(n10829) );
  NAND U11127 ( .A(n10830), .B(n10829), .Z(n10993) );
  XNOR U11128 ( .A(n10992), .B(n10993), .Z(n10994) );
  NANDN U11129 ( .A(n10832), .B(n10831), .Z(n10836) );
  NANDN U11130 ( .A(n10834), .B(n10833), .Z(n10835) );
  NAND U11131 ( .A(n10836), .B(n10835), .Z(n10995) );
  XNOR U11132 ( .A(n10994), .B(n10995), .Z(n10938) );
  XNOR U11133 ( .A(n10939), .B(n10938), .Z(n10941) );
  NANDN U11134 ( .A(n10838), .B(n10837), .Z(n10842) );
  NANDN U11135 ( .A(n10840), .B(n10839), .Z(n10841) );
  AND U11136 ( .A(n10842), .B(n10841), .Z(n10940) );
  XOR U11137 ( .A(n10941), .B(n10940), .Z(n11055) );
  NANDN U11138 ( .A(n10844), .B(n10843), .Z(n10848) );
  NANDN U11139 ( .A(n10846), .B(n10845), .Z(n10847) );
  AND U11140 ( .A(n10848), .B(n10847), .Z(n11052) );
  NANDN U11141 ( .A(n10850), .B(n10849), .Z(n10854) );
  NANDN U11142 ( .A(n10852), .B(n10851), .Z(n10853) );
  AND U11143 ( .A(n10854), .B(n10853), .Z(n10935) );
  NANDN U11144 ( .A(n10856), .B(n10855), .Z(n10860) );
  OR U11145 ( .A(n10858), .B(n10857), .Z(n10859) );
  AND U11146 ( .A(n10860), .B(n10859), .Z(n10933) );
  NANDN U11147 ( .A(n10862), .B(n10861), .Z(n10866) );
  NANDN U11148 ( .A(n10864), .B(n10863), .Z(n10865) );
  AND U11149 ( .A(n10866), .B(n10865), .Z(n10999) );
  NANDN U11150 ( .A(n10868), .B(n10867), .Z(n10872) );
  NANDN U11151 ( .A(n10870), .B(n10869), .Z(n10871) );
  NAND U11152 ( .A(n10872), .B(n10871), .Z(n10998) );
  XNOR U11153 ( .A(n10999), .B(n10998), .Z(n11000) );
  NAND U11154 ( .A(b[0]), .B(a[88]), .Z(n10873) );
  XNOR U11155 ( .A(b[1]), .B(n10873), .Z(n10875) );
  NANDN U11156 ( .A(b[0]), .B(a[87]), .Z(n10874) );
  NAND U11157 ( .A(n10875), .B(n10874), .Z(n10947) );
  NANDN U11158 ( .A(n19394), .B(n10876), .Z(n10878) );
  XOR U11159 ( .A(b[29]), .B(a[60]), .Z(n11025) );
  NANDN U11160 ( .A(n19395), .B(n11025), .Z(n10877) );
  AND U11161 ( .A(n10878), .B(n10877), .Z(n10945) );
  AND U11162 ( .A(b[31]), .B(a[56]), .Z(n10944) );
  XNOR U11163 ( .A(n10945), .B(n10944), .Z(n10946) );
  XNOR U11164 ( .A(n10947), .B(n10946), .Z(n10986) );
  NANDN U11165 ( .A(n19005), .B(n10879), .Z(n10881) );
  XOR U11166 ( .A(b[23]), .B(a[66]), .Z(n11028) );
  NANDN U11167 ( .A(n19055), .B(n11028), .Z(n10880) );
  AND U11168 ( .A(n10881), .B(n10880), .Z(n11019) );
  NANDN U11169 ( .A(n17362), .B(n10882), .Z(n10884) );
  XOR U11170 ( .A(b[7]), .B(a[82]), .Z(n11031) );
  NANDN U11171 ( .A(n17522), .B(n11031), .Z(n10883) );
  AND U11172 ( .A(n10884), .B(n10883), .Z(n11017) );
  NANDN U11173 ( .A(n19116), .B(n10885), .Z(n10887) );
  XOR U11174 ( .A(b[25]), .B(a[64]), .Z(n11034) );
  NANDN U11175 ( .A(n19179), .B(n11034), .Z(n10886) );
  NAND U11176 ( .A(n10887), .B(n10886), .Z(n11016) );
  XNOR U11177 ( .A(n11017), .B(n11016), .Z(n11018) );
  XOR U11178 ( .A(n11019), .B(n11018), .Z(n10987) );
  XNOR U11179 ( .A(n10986), .B(n10987), .Z(n10988) );
  NANDN U11180 ( .A(n18113), .B(n10888), .Z(n10890) );
  XOR U11181 ( .A(b[13]), .B(a[76]), .Z(n11037) );
  NANDN U11182 ( .A(n18229), .B(n11037), .Z(n10889) );
  AND U11183 ( .A(n10890), .B(n10889), .Z(n10981) );
  NANDN U11184 ( .A(n17888), .B(n10891), .Z(n10893) );
  XOR U11185 ( .A(b[11]), .B(a[78]), .Z(n11040) );
  NANDN U11186 ( .A(n18025), .B(n11040), .Z(n10892) );
  NAND U11187 ( .A(n10893), .B(n10892), .Z(n10980) );
  XNOR U11188 ( .A(n10981), .B(n10980), .Z(n10982) );
  NANDN U11189 ( .A(n18487), .B(n10894), .Z(n10896) );
  XOR U11190 ( .A(b[15]), .B(a[74]), .Z(n11043) );
  NANDN U11191 ( .A(n18311), .B(n11043), .Z(n10895) );
  AND U11192 ( .A(n10896), .B(n10895), .Z(n10977) );
  NANDN U11193 ( .A(n18853), .B(n10897), .Z(n10899) );
  XOR U11194 ( .A(b[21]), .B(a[68]), .Z(n11046) );
  NANDN U11195 ( .A(n18926), .B(n11046), .Z(n10898) );
  AND U11196 ( .A(n10899), .B(n10898), .Z(n10975) );
  NANDN U11197 ( .A(n17613), .B(n10900), .Z(n10902) );
  XOR U11198 ( .A(b[9]), .B(a[80]), .Z(n11049) );
  NANDN U11199 ( .A(n17739), .B(n11049), .Z(n10901) );
  NAND U11200 ( .A(n10902), .B(n10901), .Z(n10974) );
  XNOR U11201 ( .A(n10975), .B(n10974), .Z(n10976) );
  XOR U11202 ( .A(n10977), .B(n10976), .Z(n10983) );
  XOR U11203 ( .A(n10982), .B(n10983), .Z(n10989) );
  XOR U11204 ( .A(n10988), .B(n10989), .Z(n11001) );
  XNOR U11205 ( .A(n11000), .B(n11001), .Z(n10932) );
  XNOR U11206 ( .A(n10933), .B(n10932), .Z(n10934) );
  XOR U11207 ( .A(n10935), .B(n10934), .Z(n11053) );
  XNOR U11208 ( .A(n11052), .B(n11053), .Z(n11054) );
  XNOR U11209 ( .A(n11055), .B(n11054), .Z(n10928) );
  XOR U11210 ( .A(n10929), .B(n10928), .Z(n10921) );
  NANDN U11211 ( .A(n10904), .B(n10903), .Z(n10908) );
  OR U11212 ( .A(n10906), .B(n10905), .Z(n10907) );
  AND U11213 ( .A(n10908), .B(n10907), .Z(n10920) );
  XNOR U11214 ( .A(n10921), .B(n10920), .Z(n10922) );
  XNOR U11215 ( .A(n10923), .B(n10922), .Z(n10914) );
  XNOR U11216 ( .A(n10915), .B(n10914), .Z(n10916) );
  XNOR U11217 ( .A(n10917), .B(n10916), .Z(n11058) );
  XNOR U11218 ( .A(sreg[184]), .B(n11058), .Z(n11060) );
  NANDN U11219 ( .A(sreg[183]), .B(n10909), .Z(n10913) );
  NAND U11220 ( .A(n10911), .B(n10910), .Z(n10912) );
  NAND U11221 ( .A(n10913), .B(n10912), .Z(n11059) );
  XNOR U11222 ( .A(n11060), .B(n11059), .Z(c[184]) );
  NANDN U11223 ( .A(n10915), .B(n10914), .Z(n10919) );
  NANDN U11224 ( .A(n10917), .B(n10916), .Z(n10918) );
  AND U11225 ( .A(n10919), .B(n10918), .Z(n11066) );
  NANDN U11226 ( .A(n10921), .B(n10920), .Z(n10925) );
  NANDN U11227 ( .A(n10923), .B(n10922), .Z(n10924) );
  AND U11228 ( .A(n10925), .B(n10924), .Z(n11064) );
  NANDN U11229 ( .A(n10927), .B(n10926), .Z(n10931) );
  NAND U11230 ( .A(n10929), .B(n10928), .Z(n10930) );
  AND U11231 ( .A(n10931), .B(n10930), .Z(n11071) );
  NANDN U11232 ( .A(n10933), .B(n10932), .Z(n10937) );
  NANDN U11233 ( .A(n10935), .B(n10934), .Z(n10936) );
  AND U11234 ( .A(n10937), .B(n10936), .Z(n11076) );
  NANDN U11235 ( .A(n10939), .B(n10938), .Z(n10943) );
  NAND U11236 ( .A(n10941), .B(n10940), .Z(n10942) );
  AND U11237 ( .A(n10943), .B(n10942), .Z(n11075) );
  XNOR U11238 ( .A(n11076), .B(n11075), .Z(n11078) );
  NANDN U11239 ( .A(n10945), .B(n10944), .Z(n10949) );
  NANDN U11240 ( .A(n10947), .B(n10946), .Z(n10948) );
  AND U11241 ( .A(n10949), .B(n10948), .Z(n11155) );
  NANDN U11242 ( .A(n19237), .B(n10950), .Z(n10952) );
  XOR U11243 ( .A(b[27]), .B(a[63]), .Z(n11099) );
  NANDN U11244 ( .A(n19277), .B(n11099), .Z(n10951) );
  AND U11245 ( .A(n10952), .B(n10951), .Z(n11162) );
  NANDN U11246 ( .A(n17072), .B(n10953), .Z(n10955) );
  XOR U11247 ( .A(b[5]), .B(a[85]), .Z(n11102) );
  NANDN U11248 ( .A(n17223), .B(n11102), .Z(n10954) );
  AND U11249 ( .A(n10955), .B(n10954), .Z(n11160) );
  NANDN U11250 ( .A(n18673), .B(n10956), .Z(n10958) );
  XOR U11251 ( .A(b[19]), .B(a[71]), .Z(n11105) );
  NANDN U11252 ( .A(n18758), .B(n11105), .Z(n10957) );
  NAND U11253 ( .A(n10958), .B(n10957), .Z(n11159) );
  XNOR U11254 ( .A(n11160), .B(n11159), .Z(n11161) );
  XNOR U11255 ( .A(n11162), .B(n11161), .Z(n11153) );
  NANDN U11256 ( .A(n19425), .B(n10959), .Z(n10961) );
  XOR U11257 ( .A(b[31]), .B(a[59]), .Z(n11108) );
  NANDN U11258 ( .A(n19426), .B(n11108), .Z(n10960) );
  AND U11259 ( .A(n10961), .B(n10960), .Z(n11120) );
  NANDN U11260 ( .A(n17067), .B(n10962), .Z(n10964) );
  XOR U11261 ( .A(b[3]), .B(a[87]), .Z(n11111) );
  NANDN U11262 ( .A(n17068), .B(n11111), .Z(n10963) );
  AND U11263 ( .A(n10964), .B(n10963), .Z(n11118) );
  NANDN U11264 ( .A(n18514), .B(n10965), .Z(n10967) );
  XOR U11265 ( .A(b[17]), .B(a[73]), .Z(n11114) );
  NANDN U11266 ( .A(n18585), .B(n11114), .Z(n10966) );
  NAND U11267 ( .A(n10967), .B(n10966), .Z(n11117) );
  XNOR U11268 ( .A(n11118), .B(n11117), .Z(n11119) );
  XOR U11269 ( .A(n11120), .B(n11119), .Z(n11154) );
  XOR U11270 ( .A(n11153), .B(n11154), .Z(n11156) );
  XOR U11271 ( .A(n11155), .B(n11156), .Z(n11088) );
  NANDN U11272 ( .A(n10969), .B(n10968), .Z(n10973) );
  NANDN U11273 ( .A(n10971), .B(n10970), .Z(n10972) );
  AND U11274 ( .A(n10973), .B(n10972), .Z(n11141) );
  NANDN U11275 ( .A(n10975), .B(n10974), .Z(n10979) );
  NANDN U11276 ( .A(n10977), .B(n10976), .Z(n10978) );
  NAND U11277 ( .A(n10979), .B(n10978), .Z(n11142) );
  XNOR U11278 ( .A(n11141), .B(n11142), .Z(n11143) );
  NANDN U11279 ( .A(n10981), .B(n10980), .Z(n10985) );
  NANDN U11280 ( .A(n10983), .B(n10982), .Z(n10984) );
  NAND U11281 ( .A(n10985), .B(n10984), .Z(n11144) );
  XNOR U11282 ( .A(n11143), .B(n11144), .Z(n11087) );
  XNOR U11283 ( .A(n11088), .B(n11087), .Z(n11090) );
  NANDN U11284 ( .A(n10987), .B(n10986), .Z(n10991) );
  NANDN U11285 ( .A(n10989), .B(n10988), .Z(n10990) );
  AND U11286 ( .A(n10991), .B(n10990), .Z(n11089) );
  XOR U11287 ( .A(n11090), .B(n11089), .Z(n11204) );
  NANDN U11288 ( .A(n10993), .B(n10992), .Z(n10997) );
  NANDN U11289 ( .A(n10995), .B(n10994), .Z(n10996) );
  AND U11290 ( .A(n10997), .B(n10996), .Z(n11201) );
  NANDN U11291 ( .A(n10999), .B(n10998), .Z(n11003) );
  NANDN U11292 ( .A(n11001), .B(n11000), .Z(n11002) );
  AND U11293 ( .A(n11003), .B(n11002), .Z(n11084) );
  NANDN U11294 ( .A(n11005), .B(n11004), .Z(n11009) );
  OR U11295 ( .A(n11007), .B(n11006), .Z(n11008) );
  AND U11296 ( .A(n11009), .B(n11008), .Z(n11082) );
  NANDN U11297 ( .A(n11011), .B(n11010), .Z(n11015) );
  NANDN U11298 ( .A(n11013), .B(n11012), .Z(n11014) );
  AND U11299 ( .A(n11015), .B(n11014), .Z(n11148) );
  NANDN U11300 ( .A(n11017), .B(n11016), .Z(n11021) );
  NANDN U11301 ( .A(n11019), .B(n11018), .Z(n11020) );
  NAND U11302 ( .A(n11021), .B(n11020), .Z(n11147) );
  XNOR U11303 ( .A(n11148), .B(n11147), .Z(n11149) );
  NAND U11304 ( .A(b[0]), .B(a[89]), .Z(n11022) );
  XNOR U11305 ( .A(b[1]), .B(n11022), .Z(n11024) );
  NANDN U11306 ( .A(b[0]), .B(a[88]), .Z(n11023) );
  NAND U11307 ( .A(n11024), .B(n11023), .Z(n11096) );
  NANDN U11308 ( .A(n19394), .B(n11025), .Z(n11027) );
  XOR U11309 ( .A(b[29]), .B(a[61]), .Z(n11174) );
  NANDN U11310 ( .A(n19395), .B(n11174), .Z(n11026) );
  AND U11311 ( .A(n11027), .B(n11026), .Z(n11094) );
  AND U11312 ( .A(b[31]), .B(a[57]), .Z(n11093) );
  XNOR U11313 ( .A(n11094), .B(n11093), .Z(n11095) );
  XNOR U11314 ( .A(n11096), .B(n11095), .Z(n11135) );
  NANDN U11315 ( .A(n19005), .B(n11028), .Z(n11030) );
  XOR U11316 ( .A(b[23]), .B(a[67]), .Z(n11177) );
  NANDN U11317 ( .A(n19055), .B(n11177), .Z(n11029) );
  AND U11318 ( .A(n11030), .B(n11029), .Z(n11168) );
  NANDN U11319 ( .A(n17362), .B(n11031), .Z(n11033) );
  XOR U11320 ( .A(b[7]), .B(a[83]), .Z(n11180) );
  NANDN U11321 ( .A(n17522), .B(n11180), .Z(n11032) );
  AND U11322 ( .A(n11033), .B(n11032), .Z(n11166) );
  NANDN U11323 ( .A(n19116), .B(n11034), .Z(n11036) );
  XOR U11324 ( .A(b[25]), .B(a[65]), .Z(n11183) );
  NANDN U11325 ( .A(n19179), .B(n11183), .Z(n11035) );
  NAND U11326 ( .A(n11036), .B(n11035), .Z(n11165) );
  XNOR U11327 ( .A(n11166), .B(n11165), .Z(n11167) );
  XOR U11328 ( .A(n11168), .B(n11167), .Z(n11136) );
  XNOR U11329 ( .A(n11135), .B(n11136), .Z(n11137) );
  NANDN U11330 ( .A(n18113), .B(n11037), .Z(n11039) );
  XOR U11331 ( .A(b[13]), .B(a[77]), .Z(n11186) );
  NANDN U11332 ( .A(n18229), .B(n11186), .Z(n11038) );
  AND U11333 ( .A(n11039), .B(n11038), .Z(n11130) );
  NANDN U11334 ( .A(n17888), .B(n11040), .Z(n11042) );
  XOR U11335 ( .A(b[11]), .B(a[79]), .Z(n11189) );
  NANDN U11336 ( .A(n18025), .B(n11189), .Z(n11041) );
  NAND U11337 ( .A(n11042), .B(n11041), .Z(n11129) );
  XNOR U11338 ( .A(n11130), .B(n11129), .Z(n11131) );
  NANDN U11339 ( .A(n18487), .B(n11043), .Z(n11045) );
  XOR U11340 ( .A(b[15]), .B(a[75]), .Z(n11192) );
  NANDN U11341 ( .A(n18311), .B(n11192), .Z(n11044) );
  AND U11342 ( .A(n11045), .B(n11044), .Z(n11126) );
  NANDN U11343 ( .A(n18853), .B(n11046), .Z(n11048) );
  XOR U11344 ( .A(b[21]), .B(a[69]), .Z(n11195) );
  NANDN U11345 ( .A(n18926), .B(n11195), .Z(n11047) );
  AND U11346 ( .A(n11048), .B(n11047), .Z(n11124) );
  NANDN U11347 ( .A(n17613), .B(n11049), .Z(n11051) );
  XOR U11348 ( .A(b[9]), .B(a[81]), .Z(n11198) );
  NANDN U11349 ( .A(n17739), .B(n11198), .Z(n11050) );
  NAND U11350 ( .A(n11051), .B(n11050), .Z(n11123) );
  XNOR U11351 ( .A(n11124), .B(n11123), .Z(n11125) );
  XOR U11352 ( .A(n11126), .B(n11125), .Z(n11132) );
  XOR U11353 ( .A(n11131), .B(n11132), .Z(n11138) );
  XOR U11354 ( .A(n11137), .B(n11138), .Z(n11150) );
  XNOR U11355 ( .A(n11149), .B(n11150), .Z(n11081) );
  XNOR U11356 ( .A(n11082), .B(n11081), .Z(n11083) );
  XOR U11357 ( .A(n11084), .B(n11083), .Z(n11202) );
  XNOR U11358 ( .A(n11201), .B(n11202), .Z(n11203) );
  XNOR U11359 ( .A(n11204), .B(n11203), .Z(n11077) );
  XOR U11360 ( .A(n11078), .B(n11077), .Z(n11070) );
  NANDN U11361 ( .A(n11053), .B(n11052), .Z(n11057) );
  NANDN U11362 ( .A(n11055), .B(n11054), .Z(n11056) );
  AND U11363 ( .A(n11057), .B(n11056), .Z(n11069) );
  XOR U11364 ( .A(n11070), .B(n11069), .Z(n11072) );
  XNOR U11365 ( .A(n11071), .B(n11072), .Z(n11063) );
  XNOR U11366 ( .A(n11064), .B(n11063), .Z(n11065) );
  XNOR U11367 ( .A(n11066), .B(n11065), .Z(n11207) );
  XNOR U11368 ( .A(sreg[185]), .B(n11207), .Z(n11209) );
  NANDN U11369 ( .A(sreg[184]), .B(n11058), .Z(n11062) );
  NAND U11370 ( .A(n11060), .B(n11059), .Z(n11061) );
  NAND U11371 ( .A(n11062), .B(n11061), .Z(n11208) );
  XNOR U11372 ( .A(n11209), .B(n11208), .Z(c[185]) );
  NANDN U11373 ( .A(n11064), .B(n11063), .Z(n11068) );
  NANDN U11374 ( .A(n11066), .B(n11065), .Z(n11067) );
  AND U11375 ( .A(n11068), .B(n11067), .Z(n11215) );
  NANDN U11376 ( .A(n11070), .B(n11069), .Z(n11074) );
  NANDN U11377 ( .A(n11072), .B(n11071), .Z(n11073) );
  AND U11378 ( .A(n11074), .B(n11073), .Z(n11213) );
  NANDN U11379 ( .A(n11076), .B(n11075), .Z(n11080) );
  NAND U11380 ( .A(n11078), .B(n11077), .Z(n11079) );
  AND U11381 ( .A(n11080), .B(n11079), .Z(n11220) );
  NANDN U11382 ( .A(n11082), .B(n11081), .Z(n11086) );
  NANDN U11383 ( .A(n11084), .B(n11083), .Z(n11085) );
  AND U11384 ( .A(n11086), .B(n11085), .Z(n11225) );
  NANDN U11385 ( .A(n11088), .B(n11087), .Z(n11092) );
  NAND U11386 ( .A(n11090), .B(n11089), .Z(n11091) );
  AND U11387 ( .A(n11092), .B(n11091), .Z(n11224) );
  XNOR U11388 ( .A(n11225), .B(n11224), .Z(n11227) );
  NANDN U11389 ( .A(n11094), .B(n11093), .Z(n11098) );
  NANDN U11390 ( .A(n11096), .B(n11095), .Z(n11097) );
  AND U11391 ( .A(n11098), .B(n11097), .Z(n11304) );
  NANDN U11392 ( .A(n19237), .B(n11099), .Z(n11101) );
  XOR U11393 ( .A(b[27]), .B(a[64]), .Z(n11248) );
  NANDN U11394 ( .A(n19277), .B(n11248), .Z(n11100) );
  AND U11395 ( .A(n11101), .B(n11100), .Z(n11311) );
  NANDN U11396 ( .A(n17072), .B(n11102), .Z(n11104) );
  XOR U11397 ( .A(b[5]), .B(a[86]), .Z(n11251) );
  NANDN U11398 ( .A(n17223), .B(n11251), .Z(n11103) );
  AND U11399 ( .A(n11104), .B(n11103), .Z(n11309) );
  NANDN U11400 ( .A(n18673), .B(n11105), .Z(n11107) );
  XOR U11401 ( .A(b[19]), .B(a[72]), .Z(n11254) );
  NANDN U11402 ( .A(n18758), .B(n11254), .Z(n11106) );
  NAND U11403 ( .A(n11107), .B(n11106), .Z(n11308) );
  XNOR U11404 ( .A(n11309), .B(n11308), .Z(n11310) );
  XNOR U11405 ( .A(n11311), .B(n11310), .Z(n11302) );
  NANDN U11406 ( .A(n19425), .B(n11108), .Z(n11110) );
  XOR U11407 ( .A(b[31]), .B(a[60]), .Z(n11257) );
  NANDN U11408 ( .A(n19426), .B(n11257), .Z(n11109) );
  AND U11409 ( .A(n11110), .B(n11109), .Z(n11269) );
  NANDN U11410 ( .A(n17067), .B(n11111), .Z(n11113) );
  XOR U11411 ( .A(b[3]), .B(a[88]), .Z(n11260) );
  NANDN U11412 ( .A(n17068), .B(n11260), .Z(n11112) );
  AND U11413 ( .A(n11113), .B(n11112), .Z(n11267) );
  NANDN U11414 ( .A(n18514), .B(n11114), .Z(n11116) );
  XOR U11415 ( .A(b[17]), .B(a[74]), .Z(n11263) );
  NANDN U11416 ( .A(n18585), .B(n11263), .Z(n11115) );
  NAND U11417 ( .A(n11116), .B(n11115), .Z(n11266) );
  XNOR U11418 ( .A(n11267), .B(n11266), .Z(n11268) );
  XOR U11419 ( .A(n11269), .B(n11268), .Z(n11303) );
  XOR U11420 ( .A(n11302), .B(n11303), .Z(n11305) );
  XOR U11421 ( .A(n11304), .B(n11305), .Z(n11237) );
  NANDN U11422 ( .A(n11118), .B(n11117), .Z(n11122) );
  NANDN U11423 ( .A(n11120), .B(n11119), .Z(n11121) );
  AND U11424 ( .A(n11122), .B(n11121), .Z(n11290) );
  NANDN U11425 ( .A(n11124), .B(n11123), .Z(n11128) );
  NANDN U11426 ( .A(n11126), .B(n11125), .Z(n11127) );
  NAND U11427 ( .A(n11128), .B(n11127), .Z(n11291) );
  XNOR U11428 ( .A(n11290), .B(n11291), .Z(n11292) );
  NANDN U11429 ( .A(n11130), .B(n11129), .Z(n11134) );
  NANDN U11430 ( .A(n11132), .B(n11131), .Z(n11133) );
  NAND U11431 ( .A(n11134), .B(n11133), .Z(n11293) );
  XNOR U11432 ( .A(n11292), .B(n11293), .Z(n11236) );
  XNOR U11433 ( .A(n11237), .B(n11236), .Z(n11239) );
  NANDN U11434 ( .A(n11136), .B(n11135), .Z(n11140) );
  NANDN U11435 ( .A(n11138), .B(n11137), .Z(n11139) );
  AND U11436 ( .A(n11140), .B(n11139), .Z(n11238) );
  XOR U11437 ( .A(n11239), .B(n11238), .Z(n11353) );
  NANDN U11438 ( .A(n11142), .B(n11141), .Z(n11146) );
  NANDN U11439 ( .A(n11144), .B(n11143), .Z(n11145) );
  AND U11440 ( .A(n11146), .B(n11145), .Z(n11350) );
  NANDN U11441 ( .A(n11148), .B(n11147), .Z(n11152) );
  NANDN U11442 ( .A(n11150), .B(n11149), .Z(n11151) );
  AND U11443 ( .A(n11152), .B(n11151), .Z(n11233) );
  NANDN U11444 ( .A(n11154), .B(n11153), .Z(n11158) );
  OR U11445 ( .A(n11156), .B(n11155), .Z(n11157) );
  AND U11446 ( .A(n11158), .B(n11157), .Z(n11231) );
  NANDN U11447 ( .A(n11160), .B(n11159), .Z(n11164) );
  NANDN U11448 ( .A(n11162), .B(n11161), .Z(n11163) );
  AND U11449 ( .A(n11164), .B(n11163), .Z(n11297) );
  NANDN U11450 ( .A(n11166), .B(n11165), .Z(n11170) );
  NANDN U11451 ( .A(n11168), .B(n11167), .Z(n11169) );
  NAND U11452 ( .A(n11170), .B(n11169), .Z(n11296) );
  XNOR U11453 ( .A(n11297), .B(n11296), .Z(n11298) );
  NAND U11454 ( .A(b[0]), .B(a[90]), .Z(n11171) );
  XNOR U11455 ( .A(b[1]), .B(n11171), .Z(n11173) );
  NANDN U11456 ( .A(b[0]), .B(a[89]), .Z(n11172) );
  NAND U11457 ( .A(n11173), .B(n11172), .Z(n11245) );
  NANDN U11458 ( .A(n19394), .B(n11174), .Z(n11176) );
  XOR U11459 ( .A(b[29]), .B(a[62]), .Z(n11323) );
  NANDN U11460 ( .A(n19395), .B(n11323), .Z(n11175) );
  AND U11461 ( .A(n11176), .B(n11175), .Z(n11243) );
  AND U11462 ( .A(b[31]), .B(a[58]), .Z(n11242) );
  XNOR U11463 ( .A(n11243), .B(n11242), .Z(n11244) );
  XNOR U11464 ( .A(n11245), .B(n11244), .Z(n11284) );
  NANDN U11465 ( .A(n19005), .B(n11177), .Z(n11179) );
  XOR U11466 ( .A(b[23]), .B(a[68]), .Z(n11326) );
  NANDN U11467 ( .A(n19055), .B(n11326), .Z(n11178) );
  AND U11468 ( .A(n11179), .B(n11178), .Z(n11317) );
  NANDN U11469 ( .A(n17362), .B(n11180), .Z(n11182) );
  XOR U11470 ( .A(b[7]), .B(a[84]), .Z(n11329) );
  NANDN U11471 ( .A(n17522), .B(n11329), .Z(n11181) );
  AND U11472 ( .A(n11182), .B(n11181), .Z(n11315) );
  NANDN U11473 ( .A(n19116), .B(n11183), .Z(n11185) );
  XOR U11474 ( .A(b[25]), .B(a[66]), .Z(n11332) );
  NANDN U11475 ( .A(n19179), .B(n11332), .Z(n11184) );
  NAND U11476 ( .A(n11185), .B(n11184), .Z(n11314) );
  XNOR U11477 ( .A(n11315), .B(n11314), .Z(n11316) );
  XOR U11478 ( .A(n11317), .B(n11316), .Z(n11285) );
  XNOR U11479 ( .A(n11284), .B(n11285), .Z(n11286) );
  NANDN U11480 ( .A(n18113), .B(n11186), .Z(n11188) );
  XOR U11481 ( .A(b[13]), .B(a[78]), .Z(n11335) );
  NANDN U11482 ( .A(n18229), .B(n11335), .Z(n11187) );
  AND U11483 ( .A(n11188), .B(n11187), .Z(n11279) );
  NANDN U11484 ( .A(n17888), .B(n11189), .Z(n11191) );
  XOR U11485 ( .A(b[11]), .B(a[80]), .Z(n11338) );
  NANDN U11486 ( .A(n18025), .B(n11338), .Z(n11190) );
  NAND U11487 ( .A(n11191), .B(n11190), .Z(n11278) );
  XNOR U11488 ( .A(n11279), .B(n11278), .Z(n11280) );
  NANDN U11489 ( .A(n18487), .B(n11192), .Z(n11194) );
  XOR U11490 ( .A(b[15]), .B(a[76]), .Z(n11341) );
  NANDN U11491 ( .A(n18311), .B(n11341), .Z(n11193) );
  AND U11492 ( .A(n11194), .B(n11193), .Z(n11275) );
  NANDN U11493 ( .A(n18853), .B(n11195), .Z(n11197) );
  XOR U11494 ( .A(b[21]), .B(a[70]), .Z(n11344) );
  NANDN U11495 ( .A(n18926), .B(n11344), .Z(n11196) );
  AND U11496 ( .A(n11197), .B(n11196), .Z(n11273) );
  NANDN U11497 ( .A(n17613), .B(n11198), .Z(n11200) );
  XOR U11498 ( .A(b[9]), .B(a[82]), .Z(n11347) );
  NANDN U11499 ( .A(n17739), .B(n11347), .Z(n11199) );
  NAND U11500 ( .A(n11200), .B(n11199), .Z(n11272) );
  XNOR U11501 ( .A(n11273), .B(n11272), .Z(n11274) );
  XOR U11502 ( .A(n11275), .B(n11274), .Z(n11281) );
  XOR U11503 ( .A(n11280), .B(n11281), .Z(n11287) );
  XOR U11504 ( .A(n11286), .B(n11287), .Z(n11299) );
  XNOR U11505 ( .A(n11298), .B(n11299), .Z(n11230) );
  XNOR U11506 ( .A(n11231), .B(n11230), .Z(n11232) );
  XOR U11507 ( .A(n11233), .B(n11232), .Z(n11351) );
  XNOR U11508 ( .A(n11350), .B(n11351), .Z(n11352) );
  XNOR U11509 ( .A(n11353), .B(n11352), .Z(n11226) );
  XOR U11510 ( .A(n11227), .B(n11226), .Z(n11219) );
  NANDN U11511 ( .A(n11202), .B(n11201), .Z(n11206) );
  NANDN U11512 ( .A(n11204), .B(n11203), .Z(n11205) );
  AND U11513 ( .A(n11206), .B(n11205), .Z(n11218) );
  XOR U11514 ( .A(n11219), .B(n11218), .Z(n11221) );
  XNOR U11515 ( .A(n11220), .B(n11221), .Z(n11212) );
  XNOR U11516 ( .A(n11213), .B(n11212), .Z(n11214) );
  XNOR U11517 ( .A(n11215), .B(n11214), .Z(n11356) );
  XNOR U11518 ( .A(sreg[186]), .B(n11356), .Z(n11358) );
  NANDN U11519 ( .A(sreg[185]), .B(n11207), .Z(n11211) );
  NAND U11520 ( .A(n11209), .B(n11208), .Z(n11210) );
  NAND U11521 ( .A(n11211), .B(n11210), .Z(n11357) );
  XNOR U11522 ( .A(n11358), .B(n11357), .Z(c[186]) );
  NANDN U11523 ( .A(n11213), .B(n11212), .Z(n11217) );
  NANDN U11524 ( .A(n11215), .B(n11214), .Z(n11216) );
  AND U11525 ( .A(n11217), .B(n11216), .Z(n11364) );
  NANDN U11526 ( .A(n11219), .B(n11218), .Z(n11223) );
  NANDN U11527 ( .A(n11221), .B(n11220), .Z(n11222) );
  AND U11528 ( .A(n11223), .B(n11222), .Z(n11362) );
  NANDN U11529 ( .A(n11225), .B(n11224), .Z(n11229) );
  NAND U11530 ( .A(n11227), .B(n11226), .Z(n11228) );
  AND U11531 ( .A(n11229), .B(n11228), .Z(n11369) );
  NANDN U11532 ( .A(n11231), .B(n11230), .Z(n11235) );
  NANDN U11533 ( .A(n11233), .B(n11232), .Z(n11234) );
  AND U11534 ( .A(n11235), .B(n11234), .Z(n11374) );
  NANDN U11535 ( .A(n11237), .B(n11236), .Z(n11241) );
  NAND U11536 ( .A(n11239), .B(n11238), .Z(n11240) );
  AND U11537 ( .A(n11241), .B(n11240), .Z(n11373) );
  XNOR U11538 ( .A(n11374), .B(n11373), .Z(n11376) );
  NANDN U11539 ( .A(n11243), .B(n11242), .Z(n11247) );
  NANDN U11540 ( .A(n11245), .B(n11244), .Z(n11246) );
  AND U11541 ( .A(n11247), .B(n11246), .Z(n11453) );
  NANDN U11542 ( .A(n19237), .B(n11248), .Z(n11250) );
  XOR U11543 ( .A(b[27]), .B(a[65]), .Z(n11397) );
  NANDN U11544 ( .A(n19277), .B(n11397), .Z(n11249) );
  AND U11545 ( .A(n11250), .B(n11249), .Z(n11460) );
  NANDN U11546 ( .A(n17072), .B(n11251), .Z(n11253) );
  XOR U11547 ( .A(b[5]), .B(a[87]), .Z(n11400) );
  NANDN U11548 ( .A(n17223), .B(n11400), .Z(n11252) );
  AND U11549 ( .A(n11253), .B(n11252), .Z(n11458) );
  NANDN U11550 ( .A(n18673), .B(n11254), .Z(n11256) );
  XOR U11551 ( .A(b[19]), .B(a[73]), .Z(n11403) );
  NANDN U11552 ( .A(n18758), .B(n11403), .Z(n11255) );
  NAND U11553 ( .A(n11256), .B(n11255), .Z(n11457) );
  XNOR U11554 ( .A(n11458), .B(n11457), .Z(n11459) );
  XNOR U11555 ( .A(n11460), .B(n11459), .Z(n11451) );
  NANDN U11556 ( .A(n19425), .B(n11257), .Z(n11259) );
  XOR U11557 ( .A(b[31]), .B(a[61]), .Z(n11406) );
  NANDN U11558 ( .A(n19426), .B(n11406), .Z(n11258) );
  AND U11559 ( .A(n11259), .B(n11258), .Z(n11418) );
  NANDN U11560 ( .A(n17067), .B(n11260), .Z(n11262) );
  XOR U11561 ( .A(b[3]), .B(a[89]), .Z(n11409) );
  NANDN U11562 ( .A(n17068), .B(n11409), .Z(n11261) );
  AND U11563 ( .A(n11262), .B(n11261), .Z(n11416) );
  NANDN U11564 ( .A(n18514), .B(n11263), .Z(n11265) );
  XOR U11565 ( .A(b[17]), .B(a[75]), .Z(n11412) );
  NANDN U11566 ( .A(n18585), .B(n11412), .Z(n11264) );
  NAND U11567 ( .A(n11265), .B(n11264), .Z(n11415) );
  XNOR U11568 ( .A(n11416), .B(n11415), .Z(n11417) );
  XOR U11569 ( .A(n11418), .B(n11417), .Z(n11452) );
  XOR U11570 ( .A(n11451), .B(n11452), .Z(n11454) );
  XOR U11571 ( .A(n11453), .B(n11454), .Z(n11386) );
  NANDN U11572 ( .A(n11267), .B(n11266), .Z(n11271) );
  NANDN U11573 ( .A(n11269), .B(n11268), .Z(n11270) );
  AND U11574 ( .A(n11271), .B(n11270), .Z(n11439) );
  NANDN U11575 ( .A(n11273), .B(n11272), .Z(n11277) );
  NANDN U11576 ( .A(n11275), .B(n11274), .Z(n11276) );
  NAND U11577 ( .A(n11277), .B(n11276), .Z(n11440) );
  XNOR U11578 ( .A(n11439), .B(n11440), .Z(n11441) );
  NANDN U11579 ( .A(n11279), .B(n11278), .Z(n11283) );
  NANDN U11580 ( .A(n11281), .B(n11280), .Z(n11282) );
  NAND U11581 ( .A(n11283), .B(n11282), .Z(n11442) );
  XNOR U11582 ( .A(n11441), .B(n11442), .Z(n11385) );
  XNOR U11583 ( .A(n11386), .B(n11385), .Z(n11388) );
  NANDN U11584 ( .A(n11285), .B(n11284), .Z(n11289) );
  NANDN U11585 ( .A(n11287), .B(n11286), .Z(n11288) );
  AND U11586 ( .A(n11289), .B(n11288), .Z(n11387) );
  XOR U11587 ( .A(n11388), .B(n11387), .Z(n11502) );
  NANDN U11588 ( .A(n11291), .B(n11290), .Z(n11295) );
  NANDN U11589 ( .A(n11293), .B(n11292), .Z(n11294) );
  AND U11590 ( .A(n11295), .B(n11294), .Z(n11499) );
  NANDN U11591 ( .A(n11297), .B(n11296), .Z(n11301) );
  NANDN U11592 ( .A(n11299), .B(n11298), .Z(n11300) );
  AND U11593 ( .A(n11301), .B(n11300), .Z(n11382) );
  NANDN U11594 ( .A(n11303), .B(n11302), .Z(n11307) );
  OR U11595 ( .A(n11305), .B(n11304), .Z(n11306) );
  AND U11596 ( .A(n11307), .B(n11306), .Z(n11380) );
  NANDN U11597 ( .A(n11309), .B(n11308), .Z(n11313) );
  NANDN U11598 ( .A(n11311), .B(n11310), .Z(n11312) );
  AND U11599 ( .A(n11313), .B(n11312), .Z(n11446) );
  NANDN U11600 ( .A(n11315), .B(n11314), .Z(n11319) );
  NANDN U11601 ( .A(n11317), .B(n11316), .Z(n11318) );
  NAND U11602 ( .A(n11319), .B(n11318), .Z(n11445) );
  XNOR U11603 ( .A(n11446), .B(n11445), .Z(n11447) );
  NAND U11604 ( .A(b[0]), .B(a[91]), .Z(n11320) );
  XNOR U11605 ( .A(b[1]), .B(n11320), .Z(n11322) );
  NANDN U11606 ( .A(b[0]), .B(a[90]), .Z(n11321) );
  NAND U11607 ( .A(n11322), .B(n11321), .Z(n11394) );
  NANDN U11608 ( .A(n19394), .B(n11323), .Z(n11325) );
  XOR U11609 ( .A(b[29]), .B(a[63]), .Z(n11472) );
  NANDN U11610 ( .A(n19395), .B(n11472), .Z(n11324) );
  AND U11611 ( .A(n11325), .B(n11324), .Z(n11392) );
  AND U11612 ( .A(b[31]), .B(a[59]), .Z(n11391) );
  XNOR U11613 ( .A(n11392), .B(n11391), .Z(n11393) );
  XNOR U11614 ( .A(n11394), .B(n11393), .Z(n11433) );
  NANDN U11615 ( .A(n19005), .B(n11326), .Z(n11328) );
  XOR U11616 ( .A(b[23]), .B(a[69]), .Z(n11475) );
  NANDN U11617 ( .A(n19055), .B(n11475), .Z(n11327) );
  AND U11618 ( .A(n11328), .B(n11327), .Z(n11466) );
  NANDN U11619 ( .A(n17362), .B(n11329), .Z(n11331) );
  XOR U11620 ( .A(b[7]), .B(a[85]), .Z(n11478) );
  NANDN U11621 ( .A(n17522), .B(n11478), .Z(n11330) );
  AND U11622 ( .A(n11331), .B(n11330), .Z(n11464) );
  NANDN U11623 ( .A(n19116), .B(n11332), .Z(n11334) );
  XOR U11624 ( .A(b[25]), .B(a[67]), .Z(n11481) );
  NANDN U11625 ( .A(n19179), .B(n11481), .Z(n11333) );
  NAND U11626 ( .A(n11334), .B(n11333), .Z(n11463) );
  XNOR U11627 ( .A(n11464), .B(n11463), .Z(n11465) );
  XOR U11628 ( .A(n11466), .B(n11465), .Z(n11434) );
  XNOR U11629 ( .A(n11433), .B(n11434), .Z(n11435) );
  NANDN U11630 ( .A(n18113), .B(n11335), .Z(n11337) );
  XOR U11631 ( .A(b[13]), .B(a[79]), .Z(n11484) );
  NANDN U11632 ( .A(n18229), .B(n11484), .Z(n11336) );
  AND U11633 ( .A(n11337), .B(n11336), .Z(n11428) );
  NANDN U11634 ( .A(n17888), .B(n11338), .Z(n11340) );
  XOR U11635 ( .A(b[11]), .B(a[81]), .Z(n11487) );
  NANDN U11636 ( .A(n18025), .B(n11487), .Z(n11339) );
  NAND U11637 ( .A(n11340), .B(n11339), .Z(n11427) );
  XNOR U11638 ( .A(n11428), .B(n11427), .Z(n11429) );
  NANDN U11639 ( .A(n18487), .B(n11341), .Z(n11343) );
  XOR U11640 ( .A(b[15]), .B(a[77]), .Z(n11490) );
  NANDN U11641 ( .A(n18311), .B(n11490), .Z(n11342) );
  AND U11642 ( .A(n11343), .B(n11342), .Z(n11424) );
  NANDN U11643 ( .A(n18853), .B(n11344), .Z(n11346) );
  XOR U11644 ( .A(b[21]), .B(a[71]), .Z(n11493) );
  NANDN U11645 ( .A(n18926), .B(n11493), .Z(n11345) );
  AND U11646 ( .A(n11346), .B(n11345), .Z(n11422) );
  NANDN U11647 ( .A(n17613), .B(n11347), .Z(n11349) );
  XOR U11648 ( .A(b[9]), .B(a[83]), .Z(n11496) );
  NANDN U11649 ( .A(n17739), .B(n11496), .Z(n11348) );
  NAND U11650 ( .A(n11349), .B(n11348), .Z(n11421) );
  XNOR U11651 ( .A(n11422), .B(n11421), .Z(n11423) );
  XOR U11652 ( .A(n11424), .B(n11423), .Z(n11430) );
  XOR U11653 ( .A(n11429), .B(n11430), .Z(n11436) );
  XOR U11654 ( .A(n11435), .B(n11436), .Z(n11448) );
  XNOR U11655 ( .A(n11447), .B(n11448), .Z(n11379) );
  XNOR U11656 ( .A(n11380), .B(n11379), .Z(n11381) );
  XOR U11657 ( .A(n11382), .B(n11381), .Z(n11500) );
  XNOR U11658 ( .A(n11499), .B(n11500), .Z(n11501) );
  XNOR U11659 ( .A(n11502), .B(n11501), .Z(n11375) );
  XOR U11660 ( .A(n11376), .B(n11375), .Z(n11368) );
  NANDN U11661 ( .A(n11351), .B(n11350), .Z(n11355) );
  NANDN U11662 ( .A(n11353), .B(n11352), .Z(n11354) );
  AND U11663 ( .A(n11355), .B(n11354), .Z(n11367) );
  XOR U11664 ( .A(n11368), .B(n11367), .Z(n11370) );
  XNOR U11665 ( .A(n11369), .B(n11370), .Z(n11361) );
  XNOR U11666 ( .A(n11362), .B(n11361), .Z(n11363) );
  XNOR U11667 ( .A(n11364), .B(n11363), .Z(n11505) );
  XNOR U11668 ( .A(sreg[187]), .B(n11505), .Z(n11507) );
  NANDN U11669 ( .A(sreg[186]), .B(n11356), .Z(n11360) );
  NAND U11670 ( .A(n11358), .B(n11357), .Z(n11359) );
  NAND U11671 ( .A(n11360), .B(n11359), .Z(n11506) );
  XNOR U11672 ( .A(n11507), .B(n11506), .Z(c[187]) );
  NANDN U11673 ( .A(n11362), .B(n11361), .Z(n11366) );
  NANDN U11674 ( .A(n11364), .B(n11363), .Z(n11365) );
  AND U11675 ( .A(n11366), .B(n11365), .Z(n11513) );
  NANDN U11676 ( .A(n11368), .B(n11367), .Z(n11372) );
  NANDN U11677 ( .A(n11370), .B(n11369), .Z(n11371) );
  AND U11678 ( .A(n11372), .B(n11371), .Z(n11511) );
  NANDN U11679 ( .A(n11374), .B(n11373), .Z(n11378) );
  NAND U11680 ( .A(n11376), .B(n11375), .Z(n11377) );
  AND U11681 ( .A(n11378), .B(n11377), .Z(n11518) );
  NANDN U11682 ( .A(n11380), .B(n11379), .Z(n11384) );
  NANDN U11683 ( .A(n11382), .B(n11381), .Z(n11383) );
  AND U11684 ( .A(n11384), .B(n11383), .Z(n11523) );
  NANDN U11685 ( .A(n11386), .B(n11385), .Z(n11390) );
  NAND U11686 ( .A(n11388), .B(n11387), .Z(n11389) );
  AND U11687 ( .A(n11390), .B(n11389), .Z(n11522) );
  XNOR U11688 ( .A(n11523), .B(n11522), .Z(n11525) );
  NANDN U11689 ( .A(n11392), .B(n11391), .Z(n11396) );
  NANDN U11690 ( .A(n11394), .B(n11393), .Z(n11395) );
  AND U11691 ( .A(n11396), .B(n11395), .Z(n11602) );
  NANDN U11692 ( .A(n19237), .B(n11397), .Z(n11399) );
  XOR U11693 ( .A(b[27]), .B(a[66]), .Z(n11546) );
  NANDN U11694 ( .A(n19277), .B(n11546), .Z(n11398) );
  AND U11695 ( .A(n11399), .B(n11398), .Z(n11609) );
  NANDN U11696 ( .A(n17072), .B(n11400), .Z(n11402) );
  XOR U11697 ( .A(b[5]), .B(a[88]), .Z(n11549) );
  NANDN U11698 ( .A(n17223), .B(n11549), .Z(n11401) );
  AND U11699 ( .A(n11402), .B(n11401), .Z(n11607) );
  NANDN U11700 ( .A(n18673), .B(n11403), .Z(n11405) );
  XOR U11701 ( .A(b[19]), .B(a[74]), .Z(n11552) );
  NANDN U11702 ( .A(n18758), .B(n11552), .Z(n11404) );
  NAND U11703 ( .A(n11405), .B(n11404), .Z(n11606) );
  XNOR U11704 ( .A(n11607), .B(n11606), .Z(n11608) );
  XNOR U11705 ( .A(n11609), .B(n11608), .Z(n11600) );
  NANDN U11706 ( .A(n19425), .B(n11406), .Z(n11408) );
  XOR U11707 ( .A(b[31]), .B(a[62]), .Z(n11555) );
  NANDN U11708 ( .A(n19426), .B(n11555), .Z(n11407) );
  AND U11709 ( .A(n11408), .B(n11407), .Z(n11567) );
  NANDN U11710 ( .A(n17067), .B(n11409), .Z(n11411) );
  XOR U11711 ( .A(b[3]), .B(a[90]), .Z(n11558) );
  NANDN U11712 ( .A(n17068), .B(n11558), .Z(n11410) );
  AND U11713 ( .A(n11411), .B(n11410), .Z(n11565) );
  NANDN U11714 ( .A(n18514), .B(n11412), .Z(n11414) );
  XOR U11715 ( .A(b[17]), .B(a[76]), .Z(n11561) );
  NANDN U11716 ( .A(n18585), .B(n11561), .Z(n11413) );
  NAND U11717 ( .A(n11414), .B(n11413), .Z(n11564) );
  XNOR U11718 ( .A(n11565), .B(n11564), .Z(n11566) );
  XOR U11719 ( .A(n11567), .B(n11566), .Z(n11601) );
  XOR U11720 ( .A(n11600), .B(n11601), .Z(n11603) );
  XOR U11721 ( .A(n11602), .B(n11603), .Z(n11535) );
  NANDN U11722 ( .A(n11416), .B(n11415), .Z(n11420) );
  NANDN U11723 ( .A(n11418), .B(n11417), .Z(n11419) );
  AND U11724 ( .A(n11420), .B(n11419), .Z(n11588) );
  NANDN U11725 ( .A(n11422), .B(n11421), .Z(n11426) );
  NANDN U11726 ( .A(n11424), .B(n11423), .Z(n11425) );
  NAND U11727 ( .A(n11426), .B(n11425), .Z(n11589) );
  XNOR U11728 ( .A(n11588), .B(n11589), .Z(n11590) );
  NANDN U11729 ( .A(n11428), .B(n11427), .Z(n11432) );
  NANDN U11730 ( .A(n11430), .B(n11429), .Z(n11431) );
  NAND U11731 ( .A(n11432), .B(n11431), .Z(n11591) );
  XNOR U11732 ( .A(n11590), .B(n11591), .Z(n11534) );
  XNOR U11733 ( .A(n11535), .B(n11534), .Z(n11537) );
  NANDN U11734 ( .A(n11434), .B(n11433), .Z(n11438) );
  NANDN U11735 ( .A(n11436), .B(n11435), .Z(n11437) );
  AND U11736 ( .A(n11438), .B(n11437), .Z(n11536) );
  XOR U11737 ( .A(n11537), .B(n11536), .Z(n11651) );
  NANDN U11738 ( .A(n11440), .B(n11439), .Z(n11444) );
  NANDN U11739 ( .A(n11442), .B(n11441), .Z(n11443) );
  AND U11740 ( .A(n11444), .B(n11443), .Z(n11648) );
  NANDN U11741 ( .A(n11446), .B(n11445), .Z(n11450) );
  NANDN U11742 ( .A(n11448), .B(n11447), .Z(n11449) );
  AND U11743 ( .A(n11450), .B(n11449), .Z(n11531) );
  NANDN U11744 ( .A(n11452), .B(n11451), .Z(n11456) );
  OR U11745 ( .A(n11454), .B(n11453), .Z(n11455) );
  AND U11746 ( .A(n11456), .B(n11455), .Z(n11529) );
  NANDN U11747 ( .A(n11458), .B(n11457), .Z(n11462) );
  NANDN U11748 ( .A(n11460), .B(n11459), .Z(n11461) );
  AND U11749 ( .A(n11462), .B(n11461), .Z(n11595) );
  NANDN U11750 ( .A(n11464), .B(n11463), .Z(n11468) );
  NANDN U11751 ( .A(n11466), .B(n11465), .Z(n11467) );
  NAND U11752 ( .A(n11468), .B(n11467), .Z(n11594) );
  XNOR U11753 ( .A(n11595), .B(n11594), .Z(n11596) );
  NAND U11754 ( .A(b[0]), .B(a[92]), .Z(n11469) );
  XNOR U11755 ( .A(b[1]), .B(n11469), .Z(n11471) );
  NANDN U11756 ( .A(b[0]), .B(a[91]), .Z(n11470) );
  NAND U11757 ( .A(n11471), .B(n11470), .Z(n11543) );
  NANDN U11758 ( .A(n19394), .B(n11472), .Z(n11474) );
  XOR U11759 ( .A(b[29]), .B(a[64]), .Z(n11621) );
  NANDN U11760 ( .A(n19395), .B(n11621), .Z(n11473) );
  AND U11761 ( .A(n11474), .B(n11473), .Z(n11541) );
  AND U11762 ( .A(b[31]), .B(a[60]), .Z(n11540) );
  XNOR U11763 ( .A(n11541), .B(n11540), .Z(n11542) );
  XNOR U11764 ( .A(n11543), .B(n11542), .Z(n11582) );
  NANDN U11765 ( .A(n19005), .B(n11475), .Z(n11477) );
  XOR U11766 ( .A(b[23]), .B(a[70]), .Z(n11624) );
  NANDN U11767 ( .A(n19055), .B(n11624), .Z(n11476) );
  AND U11768 ( .A(n11477), .B(n11476), .Z(n11615) );
  NANDN U11769 ( .A(n17362), .B(n11478), .Z(n11480) );
  XOR U11770 ( .A(b[7]), .B(a[86]), .Z(n11627) );
  NANDN U11771 ( .A(n17522), .B(n11627), .Z(n11479) );
  AND U11772 ( .A(n11480), .B(n11479), .Z(n11613) );
  NANDN U11773 ( .A(n19116), .B(n11481), .Z(n11483) );
  XOR U11774 ( .A(b[25]), .B(a[68]), .Z(n11630) );
  NANDN U11775 ( .A(n19179), .B(n11630), .Z(n11482) );
  NAND U11776 ( .A(n11483), .B(n11482), .Z(n11612) );
  XNOR U11777 ( .A(n11613), .B(n11612), .Z(n11614) );
  XOR U11778 ( .A(n11615), .B(n11614), .Z(n11583) );
  XNOR U11779 ( .A(n11582), .B(n11583), .Z(n11584) );
  NANDN U11780 ( .A(n18113), .B(n11484), .Z(n11486) );
  XOR U11781 ( .A(b[13]), .B(a[80]), .Z(n11633) );
  NANDN U11782 ( .A(n18229), .B(n11633), .Z(n11485) );
  AND U11783 ( .A(n11486), .B(n11485), .Z(n11577) );
  NANDN U11784 ( .A(n17888), .B(n11487), .Z(n11489) );
  XOR U11785 ( .A(b[11]), .B(a[82]), .Z(n11636) );
  NANDN U11786 ( .A(n18025), .B(n11636), .Z(n11488) );
  NAND U11787 ( .A(n11489), .B(n11488), .Z(n11576) );
  XNOR U11788 ( .A(n11577), .B(n11576), .Z(n11578) );
  NANDN U11789 ( .A(n18487), .B(n11490), .Z(n11492) );
  XOR U11790 ( .A(b[15]), .B(a[78]), .Z(n11639) );
  NANDN U11791 ( .A(n18311), .B(n11639), .Z(n11491) );
  AND U11792 ( .A(n11492), .B(n11491), .Z(n11573) );
  NANDN U11793 ( .A(n18853), .B(n11493), .Z(n11495) );
  XOR U11794 ( .A(b[21]), .B(a[72]), .Z(n11642) );
  NANDN U11795 ( .A(n18926), .B(n11642), .Z(n11494) );
  AND U11796 ( .A(n11495), .B(n11494), .Z(n11571) );
  NANDN U11797 ( .A(n17613), .B(n11496), .Z(n11498) );
  XOR U11798 ( .A(b[9]), .B(a[84]), .Z(n11645) );
  NANDN U11799 ( .A(n17739), .B(n11645), .Z(n11497) );
  NAND U11800 ( .A(n11498), .B(n11497), .Z(n11570) );
  XNOR U11801 ( .A(n11571), .B(n11570), .Z(n11572) );
  XOR U11802 ( .A(n11573), .B(n11572), .Z(n11579) );
  XOR U11803 ( .A(n11578), .B(n11579), .Z(n11585) );
  XOR U11804 ( .A(n11584), .B(n11585), .Z(n11597) );
  XNOR U11805 ( .A(n11596), .B(n11597), .Z(n11528) );
  XNOR U11806 ( .A(n11529), .B(n11528), .Z(n11530) );
  XOR U11807 ( .A(n11531), .B(n11530), .Z(n11649) );
  XNOR U11808 ( .A(n11648), .B(n11649), .Z(n11650) );
  XNOR U11809 ( .A(n11651), .B(n11650), .Z(n11524) );
  XOR U11810 ( .A(n11525), .B(n11524), .Z(n11517) );
  NANDN U11811 ( .A(n11500), .B(n11499), .Z(n11504) );
  NANDN U11812 ( .A(n11502), .B(n11501), .Z(n11503) );
  AND U11813 ( .A(n11504), .B(n11503), .Z(n11516) );
  XOR U11814 ( .A(n11517), .B(n11516), .Z(n11519) );
  XNOR U11815 ( .A(n11518), .B(n11519), .Z(n11510) );
  XNOR U11816 ( .A(n11511), .B(n11510), .Z(n11512) );
  XNOR U11817 ( .A(n11513), .B(n11512), .Z(n11654) );
  XNOR U11818 ( .A(sreg[188]), .B(n11654), .Z(n11656) );
  NANDN U11819 ( .A(sreg[187]), .B(n11505), .Z(n11509) );
  NAND U11820 ( .A(n11507), .B(n11506), .Z(n11508) );
  NAND U11821 ( .A(n11509), .B(n11508), .Z(n11655) );
  XNOR U11822 ( .A(n11656), .B(n11655), .Z(c[188]) );
  NANDN U11823 ( .A(n11511), .B(n11510), .Z(n11515) );
  NANDN U11824 ( .A(n11513), .B(n11512), .Z(n11514) );
  AND U11825 ( .A(n11515), .B(n11514), .Z(n11662) );
  NANDN U11826 ( .A(n11517), .B(n11516), .Z(n11521) );
  NANDN U11827 ( .A(n11519), .B(n11518), .Z(n11520) );
  AND U11828 ( .A(n11521), .B(n11520), .Z(n11660) );
  NANDN U11829 ( .A(n11523), .B(n11522), .Z(n11527) );
  NAND U11830 ( .A(n11525), .B(n11524), .Z(n11526) );
  AND U11831 ( .A(n11527), .B(n11526), .Z(n11667) );
  NANDN U11832 ( .A(n11529), .B(n11528), .Z(n11533) );
  NANDN U11833 ( .A(n11531), .B(n11530), .Z(n11532) );
  AND U11834 ( .A(n11533), .B(n11532), .Z(n11672) );
  NANDN U11835 ( .A(n11535), .B(n11534), .Z(n11539) );
  NAND U11836 ( .A(n11537), .B(n11536), .Z(n11538) );
  AND U11837 ( .A(n11539), .B(n11538), .Z(n11671) );
  XNOR U11838 ( .A(n11672), .B(n11671), .Z(n11674) );
  NANDN U11839 ( .A(n11541), .B(n11540), .Z(n11545) );
  NANDN U11840 ( .A(n11543), .B(n11542), .Z(n11544) );
  AND U11841 ( .A(n11545), .B(n11544), .Z(n11751) );
  NANDN U11842 ( .A(n19237), .B(n11546), .Z(n11548) );
  XOR U11843 ( .A(b[27]), .B(a[67]), .Z(n11695) );
  NANDN U11844 ( .A(n19277), .B(n11695), .Z(n11547) );
  AND U11845 ( .A(n11548), .B(n11547), .Z(n11758) );
  NANDN U11846 ( .A(n17072), .B(n11549), .Z(n11551) );
  XOR U11847 ( .A(b[5]), .B(a[89]), .Z(n11698) );
  NANDN U11848 ( .A(n17223), .B(n11698), .Z(n11550) );
  AND U11849 ( .A(n11551), .B(n11550), .Z(n11756) );
  NANDN U11850 ( .A(n18673), .B(n11552), .Z(n11554) );
  XOR U11851 ( .A(b[19]), .B(a[75]), .Z(n11701) );
  NANDN U11852 ( .A(n18758), .B(n11701), .Z(n11553) );
  NAND U11853 ( .A(n11554), .B(n11553), .Z(n11755) );
  XNOR U11854 ( .A(n11756), .B(n11755), .Z(n11757) );
  XNOR U11855 ( .A(n11758), .B(n11757), .Z(n11749) );
  NANDN U11856 ( .A(n19425), .B(n11555), .Z(n11557) );
  XOR U11857 ( .A(b[31]), .B(a[63]), .Z(n11704) );
  NANDN U11858 ( .A(n19426), .B(n11704), .Z(n11556) );
  AND U11859 ( .A(n11557), .B(n11556), .Z(n11716) );
  NANDN U11860 ( .A(n17067), .B(n11558), .Z(n11560) );
  XOR U11861 ( .A(b[3]), .B(a[91]), .Z(n11707) );
  NANDN U11862 ( .A(n17068), .B(n11707), .Z(n11559) );
  AND U11863 ( .A(n11560), .B(n11559), .Z(n11714) );
  NANDN U11864 ( .A(n18514), .B(n11561), .Z(n11563) );
  XOR U11865 ( .A(b[17]), .B(a[77]), .Z(n11710) );
  NANDN U11866 ( .A(n18585), .B(n11710), .Z(n11562) );
  NAND U11867 ( .A(n11563), .B(n11562), .Z(n11713) );
  XNOR U11868 ( .A(n11714), .B(n11713), .Z(n11715) );
  XOR U11869 ( .A(n11716), .B(n11715), .Z(n11750) );
  XOR U11870 ( .A(n11749), .B(n11750), .Z(n11752) );
  XOR U11871 ( .A(n11751), .B(n11752), .Z(n11684) );
  NANDN U11872 ( .A(n11565), .B(n11564), .Z(n11569) );
  NANDN U11873 ( .A(n11567), .B(n11566), .Z(n11568) );
  AND U11874 ( .A(n11569), .B(n11568), .Z(n11737) );
  NANDN U11875 ( .A(n11571), .B(n11570), .Z(n11575) );
  NANDN U11876 ( .A(n11573), .B(n11572), .Z(n11574) );
  NAND U11877 ( .A(n11575), .B(n11574), .Z(n11738) );
  XNOR U11878 ( .A(n11737), .B(n11738), .Z(n11739) );
  NANDN U11879 ( .A(n11577), .B(n11576), .Z(n11581) );
  NANDN U11880 ( .A(n11579), .B(n11578), .Z(n11580) );
  NAND U11881 ( .A(n11581), .B(n11580), .Z(n11740) );
  XNOR U11882 ( .A(n11739), .B(n11740), .Z(n11683) );
  XNOR U11883 ( .A(n11684), .B(n11683), .Z(n11686) );
  NANDN U11884 ( .A(n11583), .B(n11582), .Z(n11587) );
  NANDN U11885 ( .A(n11585), .B(n11584), .Z(n11586) );
  AND U11886 ( .A(n11587), .B(n11586), .Z(n11685) );
  XOR U11887 ( .A(n11686), .B(n11685), .Z(n11800) );
  NANDN U11888 ( .A(n11589), .B(n11588), .Z(n11593) );
  NANDN U11889 ( .A(n11591), .B(n11590), .Z(n11592) );
  AND U11890 ( .A(n11593), .B(n11592), .Z(n11797) );
  NANDN U11891 ( .A(n11595), .B(n11594), .Z(n11599) );
  NANDN U11892 ( .A(n11597), .B(n11596), .Z(n11598) );
  AND U11893 ( .A(n11599), .B(n11598), .Z(n11680) );
  NANDN U11894 ( .A(n11601), .B(n11600), .Z(n11605) );
  OR U11895 ( .A(n11603), .B(n11602), .Z(n11604) );
  AND U11896 ( .A(n11605), .B(n11604), .Z(n11678) );
  NANDN U11897 ( .A(n11607), .B(n11606), .Z(n11611) );
  NANDN U11898 ( .A(n11609), .B(n11608), .Z(n11610) );
  AND U11899 ( .A(n11611), .B(n11610), .Z(n11744) );
  NANDN U11900 ( .A(n11613), .B(n11612), .Z(n11617) );
  NANDN U11901 ( .A(n11615), .B(n11614), .Z(n11616) );
  NAND U11902 ( .A(n11617), .B(n11616), .Z(n11743) );
  XNOR U11903 ( .A(n11744), .B(n11743), .Z(n11745) );
  NAND U11904 ( .A(b[0]), .B(a[93]), .Z(n11618) );
  XNOR U11905 ( .A(b[1]), .B(n11618), .Z(n11620) );
  NANDN U11906 ( .A(b[0]), .B(a[92]), .Z(n11619) );
  NAND U11907 ( .A(n11620), .B(n11619), .Z(n11692) );
  NANDN U11908 ( .A(n19394), .B(n11621), .Z(n11623) );
  XOR U11909 ( .A(b[29]), .B(a[65]), .Z(n11770) );
  NANDN U11910 ( .A(n19395), .B(n11770), .Z(n11622) );
  AND U11911 ( .A(n11623), .B(n11622), .Z(n11690) );
  AND U11912 ( .A(b[31]), .B(a[61]), .Z(n11689) );
  XNOR U11913 ( .A(n11690), .B(n11689), .Z(n11691) );
  XNOR U11914 ( .A(n11692), .B(n11691), .Z(n11731) );
  NANDN U11915 ( .A(n19005), .B(n11624), .Z(n11626) );
  XOR U11916 ( .A(b[23]), .B(a[71]), .Z(n11773) );
  NANDN U11917 ( .A(n19055), .B(n11773), .Z(n11625) );
  AND U11918 ( .A(n11626), .B(n11625), .Z(n11764) );
  NANDN U11919 ( .A(n17362), .B(n11627), .Z(n11629) );
  XOR U11920 ( .A(b[7]), .B(a[87]), .Z(n11776) );
  NANDN U11921 ( .A(n17522), .B(n11776), .Z(n11628) );
  AND U11922 ( .A(n11629), .B(n11628), .Z(n11762) );
  NANDN U11923 ( .A(n19116), .B(n11630), .Z(n11632) );
  XOR U11924 ( .A(b[25]), .B(a[69]), .Z(n11779) );
  NANDN U11925 ( .A(n19179), .B(n11779), .Z(n11631) );
  NAND U11926 ( .A(n11632), .B(n11631), .Z(n11761) );
  XNOR U11927 ( .A(n11762), .B(n11761), .Z(n11763) );
  XOR U11928 ( .A(n11764), .B(n11763), .Z(n11732) );
  XNOR U11929 ( .A(n11731), .B(n11732), .Z(n11733) );
  NANDN U11930 ( .A(n18113), .B(n11633), .Z(n11635) );
  XOR U11931 ( .A(b[13]), .B(a[81]), .Z(n11782) );
  NANDN U11932 ( .A(n18229), .B(n11782), .Z(n11634) );
  AND U11933 ( .A(n11635), .B(n11634), .Z(n11726) );
  NANDN U11934 ( .A(n17888), .B(n11636), .Z(n11638) );
  XOR U11935 ( .A(b[11]), .B(a[83]), .Z(n11785) );
  NANDN U11936 ( .A(n18025), .B(n11785), .Z(n11637) );
  NAND U11937 ( .A(n11638), .B(n11637), .Z(n11725) );
  XNOR U11938 ( .A(n11726), .B(n11725), .Z(n11727) );
  NANDN U11939 ( .A(n18487), .B(n11639), .Z(n11641) );
  XOR U11940 ( .A(b[15]), .B(a[79]), .Z(n11788) );
  NANDN U11941 ( .A(n18311), .B(n11788), .Z(n11640) );
  AND U11942 ( .A(n11641), .B(n11640), .Z(n11722) );
  NANDN U11943 ( .A(n18853), .B(n11642), .Z(n11644) );
  XOR U11944 ( .A(b[21]), .B(a[73]), .Z(n11791) );
  NANDN U11945 ( .A(n18926), .B(n11791), .Z(n11643) );
  AND U11946 ( .A(n11644), .B(n11643), .Z(n11720) );
  NANDN U11947 ( .A(n17613), .B(n11645), .Z(n11647) );
  XOR U11948 ( .A(b[9]), .B(a[85]), .Z(n11794) );
  NANDN U11949 ( .A(n17739), .B(n11794), .Z(n11646) );
  NAND U11950 ( .A(n11647), .B(n11646), .Z(n11719) );
  XNOR U11951 ( .A(n11720), .B(n11719), .Z(n11721) );
  XOR U11952 ( .A(n11722), .B(n11721), .Z(n11728) );
  XOR U11953 ( .A(n11727), .B(n11728), .Z(n11734) );
  XOR U11954 ( .A(n11733), .B(n11734), .Z(n11746) );
  XNOR U11955 ( .A(n11745), .B(n11746), .Z(n11677) );
  XNOR U11956 ( .A(n11678), .B(n11677), .Z(n11679) );
  XOR U11957 ( .A(n11680), .B(n11679), .Z(n11798) );
  XNOR U11958 ( .A(n11797), .B(n11798), .Z(n11799) );
  XNOR U11959 ( .A(n11800), .B(n11799), .Z(n11673) );
  XOR U11960 ( .A(n11674), .B(n11673), .Z(n11666) );
  NANDN U11961 ( .A(n11649), .B(n11648), .Z(n11653) );
  NANDN U11962 ( .A(n11651), .B(n11650), .Z(n11652) );
  AND U11963 ( .A(n11653), .B(n11652), .Z(n11665) );
  XOR U11964 ( .A(n11666), .B(n11665), .Z(n11668) );
  XNOR U11965 ( .A(n11667), .B(n11668), .Z(n11659) );
  XNOR U11966 ( .A(n11660), .B(n11659), .Z(n11661) );
  XNOR U11967 ( .A(n11662), .B(n11661), .Z(n11803) );
  XNOR U11968 ( .A(sreg[189]), .B(n11803), .Z(n11805) );
  NANDN U11969 ( .A(sreg[188]), .B(n11654), .Z(n11658) );
  NAND U11970 ( .A(n11656), .B(n11655), .Z(n11657) );
  NAND U11971 ( .A(n11658), .B(n11657), .Z(n11804) );
  XNOR U11972 ( .A(n11805), .B(n11804), .Z(c[189]) );
  NANDN U11973 ( .A(n11660), .B(n11659), .Z(n11664) );
  NANDN U11974 ( .A(n11662), .B(n11661), .Z(n11663) );
  AND U11975 ( .A(n11664), .B(n11663), .Z(n11811) );
  NANDN U11976 ( .A(n11666), .B(n11665), .Z(n11670) );
  NANDN U11977 ( .A(n11668), .B(n11667), .Z(n11669) );
  AND U11978 ( .A(n11670), .B(n11669), .Z(n11809) );
  NANDN U11979 ( .A(n11672), .B(n11671), .Z(n11676) );
  NAND U11980 ( .A(n11674), .B(n11673), .Z(n11675) );
  AND U11981 ( .A(n11676), .B(n11675), .Z(n11816) );
  NANDN U11982 ( .A(n11678), .B(n11677), .Z(n11682) );
  NANDN U11983 ( .A(n11680), .B(n11679), .Z(n11681) );
  AND U11984 ( .A(n11682), .B(n11681), .Z(n11821) );
  NANDN U11985 ( .A(n11684), .B(n11683), .Z(n11688) );
  NAND U11986 ( .A(n11686), .B(n11685), .Z(n11687) );
  AND U11987 ( .A(n11688), .B(n11687), .Z(n11820) );
  XNOR U11988 ( .A(n11821), .B(n11820), .Z(n11823) );
  NANDN U11989 ( .A(n11690), .B(n11689), .Z(n11694) );
  NANDN U11990 ( .A(n11692), .B(n11691), .Z(n11693) );
  AND U11991 ( .A(n11694), .B(n11693), .Z(n11900) );
  NANDN U11992 ( .A(n19237), .B(n11695), .Z(n11697) );
  XOR U11993 ( .A(b[27]), .B(a[68]), .Z(n11844) );
  NANDN U11994 ( .A(n19277), .B(n11844), .Z(n11696) );
  AND U11995 ( .A(n11697), .B(n11696), .Z(n11907) );
  NANDN U11996 ( .A(n17072), .B(n11698), .Z(n11700) );
  XOR U11997 ( .A(b[5]), .B(a[90]), .Z(n11847) );
  NANDN U11998 ( .A(n17223), .B(n11847), .Z(n11699) );
  AND U11999 ( .A(n11700), .B(n11699), .Z(n11905) );
  NANDN U12000 ( .A(n18673), .B(n11701), .Z(n11703) );
  XOR U12001 ( .A(b[19]), .B(a[76]), .Z(n11850) );
  NANDN U12002 ( .A(n18758), .B(n11850), .Z(n11702) );
  NAND U12003 ( .A(n11703), .B(n11702), .Z(n11904) );
  XNOR U12004 ( .A(n11905), .B(n11904), .Z(n11906) );
  XNOR U12005 ( .A(n11907), .B(n11906), .Z(n11898) );
  NANDN U12006 ( .A(n19425), .B(n11704), .Z(n11706) );
  XOR U12007 ( .A(b[31]), .B(a[64]), .Z(n11853) );
  NANDN U12008 ( .A(n19426), .B(n11853), .Z(n11705) );
  AND U12009 ( .A(n11706), .B(n11705), .Z(n11865) );
  NANDN U12010 ( .A(n17067), .B(n11707), .Z(n11709) );
  XOR U12011 ( .A(b[3]), .B(a[92]), .Z(n11856) );
  NANDN U12012 ( .A(n17068), .B(n11856), .Z(n11708) );
  AND U12013 ( .A(n11709), .B(n11708), .Z(n11863) );
  NANDN U12014 ( .A(n18514), .B(n11710), .Z(n11712) );
  XOR U12015 ( .A(b[17]), .B(a[78]), .Z(n11859) );
  NANDN U12016 ( .A(n18585), .B(n11859), .Z(n11711) );
  NAND U12017 ( .A(n11712), .B(n11711), .Z(n11862) );
  XNOR U12018 ( .A(n11863), .B(n11862), .Z(n11864) );
  XOR U12019 ( .A(n11865), .B(n11864), .Z(n11899) );
  XOR U12020 ( .A(n11898), .B(n11899), .Z(n11901) );
  XOR U12021 ( .A(n11900), .B(n11901), .Z(n11833) );
  NANDN U12022 ( .A(n11714), .B(n11713), .Z(n11718) );
  NANDN U12023 ( .A(n11716), .B(n11715), .Z(n11717) );
  AND U12024 ( .A(n11718), .B(n11717), .Z(n11886) );
  NANDN U12025 ( .A(n11720), .B(n11719), .Z(n11724) );
  NANDN U12026 ( .A(n11722), .B(n11721), .Z(n11723) );
  NAND U12027 ( .A(n11724), .B(n11723), .Z(n11887) );
  XNOR U12028 ( .A(n11886), .B(n11887), .Z(n11888) );
  NANDN U12029 ( .A(n11726), .B(n11725), .Z(n11730) );
  NANDN U12030 ( .A(n11728), .B(n11727), .Z(n11729) );
  NAND U12031 ( .A(n11730), .B(n11729), .Z(n11889) );
  XNOR U12032 ( .A(n11888), .B(n11889), .Z(n11832) );
  XNOR U12033 ( .A(n11833), .B(n11832), .Z(n11835) );
  NANDN U12034 ( .A(n11732), .B(n11731), .Z(n11736) );
  NANDN U12035 ( .A(n11734), .B(n11733), .Z(n11735) );
  AND U12036 ( .A(n11736), .B(n11735), .Z(n11834) );
  XOR U12037 ( .A(n11835), .B(n11834), .Z(n11949) );
  NANDN U12038 ( .A(n11738), .B(n11737), .Z(n11742) );
  NANDN U12039 ( .A(n11740), .B(n11739), .Z(n11741) );
  AND U12040 ( .A(n11742), .B(n11741), .Z(n11946) );
  NANDN U12041 ( .A(n11744), .B(n11743), .Z(n11748) );
  NANDN U12042 ( .A(n11746), .B(n11745), .Z(n11747) );
  AND U12043 ( .A(n11748), .B(n11747), .Z(n11829) );
  NANDN U12044 ( .A(n11750), .B(n11749), .Z(n11754) );
  OR U12045 ( .A(n11752), .B(n11751), .Z(n11753) );
  AND U12046 ( .A(n11754), .B(n11753), .Z(n11827) );
  NANDN U12047 ( .A(n11756), .B(n11755), .Z(n11760) );
  NANDN U12048 ( .A(n11758), .B(n11757), .Z(n11759) );
  AND U12049 ( .A(n11760), .B(n11759), .Z(n11893) );
  NANDN U12050 ( .A(n11762), .B(n11761), .Z(n11766) );
  NANDN U12051 ( .A(n11764), .B(n11763), .Z(n11765) );
  NAND U12052 ( .A(n11766), .B(n11765), .Z(n11892) );
  XNOR U12053 ( .A(n11893), .B(n11892), .Z(n11894) );
  NAND U12054 ( .A(b[0]), .B(a[94]), .Z(n11767) );
  XNOR U12055 ( .A(b[1]), .B(n11767), .Z(n11769) );
  NANDN U12056 ( .A(b[0]), .B(a[93]), .Z(n11768) );
  NAND U12057 ( .A(n11769), .B(n11768), .Z(n11841) );
  NANDN U12058 ( .A(n19394), .B(n11770), .Z(n11772) );
  XOR U12059 ( .A(b[29]), .B(a[66]), .Z(n11919) );
  NANDN U12060 ( .A(n19395), .B(n11919), .Z(n11771) );
  AND U12061 ( .A(n11772), .B(n11771), .Z(n11839) );
  AND U12062 ( .A(b[31]), .B(a[62]), .Z(n11838) );
  XNOR U12063 ( .A(n11839), .B(n11838), .Z(n11840) );
  XNOR U12064 ( .A(n11841), .B(n11840), .Z(n11880) );
  NANDN U12065 ( .A(n19005), .B(n11773), .Z(n11775) );
  XOR U12066 ( .A(b[23]), .B(a[72]), .Z(n11922) );
  NANDN U12067 ( .A(n19055), .B(n11922), .Z(n11774) );
  AND U12068 ( .A(n11775), .B(n11774), .Z(n11913) );
  NANDN U12069 ( .A(n17362), .B(n11776), .Z(n11778) );
  XOR U12070 ( .A(b[7]), .B(a[88]), .Z(n11925) );
  NANDN U12071 ( .A(n17522), .B(n11925), .Z(n11777) );
  AND U12072 ( .A(n11778), .B(n11777), .Z(n11911) );
  NANDN U12073 ( .A(n19116), .B(n11779), .Z(n11781) );
  XOR U12074 ( .A(b[25]), .B(a[70]), .Z(n11928) );
  NANDN U12075 ( .A(n19179), .B(n11928), .Z(n11780) );
  NAND U12076 ( .A(n11781), .B(n11780), .Z(n11910) );
  XNOR U12077 ( .A(n11911), .B(n11910), .Z(n11912) );
  XOR U12078 ( .A(n11913), .B(n11912), .Z(n11881) );
  XNOR U12079 ( .A(n11880), .B(n11881), .Z(n11882) );
  NANDN U12080 ( .A(n18113), .B(n11782), .Z(n11784) );
  XOR U12081 ( .A(b[13]), .B(a[82]), .Z(n11931) );
  NANDN U12082 ( .A(n18229), .B(n11931), .Z(n11783) );
  AND U12083 ( .A(n11784), .B(n11783), .Z(n11875) );
  NANDN U12084 ( .A(n17888), .B(n11785), .Z(n11787) );
  XOR U12085 ( .A(b[11]), .B(a[84]), .Z(n11934) );
  NANDN U12086 ( .A(n18025), .B(n11934), .Z(n11786) );
  NAND U12087 ( .A(n11787), .B(n11786), .Z(n11874) );
  XNOR U12088 ( .A(n11875), .B(n11874), .Z(n11876) );
  NANDN U12089 ( .A(n18487), .B(n11788), .Z(n11790) );
  XOR U12090 ( .A(b[15]), .B(a[80]), .Z(n11937) );
  NANDN U12091 ( .A(n18311), .B(n11937), .Z(n11789) );
  AND U12092 ( .A(n11790), .B(n11789), .Z(n11871) );
  NANDN U12093 ( .A(n18853), .B(n11791), .Z(n11793) );
  XOR U12094 ( .A(b[21]), .B(a[74]), .Z(n11940) );
  NANDN U12095 ( .A(n18926), .B(n11940), .Z(n11792) );
  AND U12096 ( .A(n11793), .B(n11792), .Z(n11869) );
  NANDN U12097 ( .A(n17613), .B(n11794), .Z(n11796) );
  XOR U12098 ( .A(b[9]), .B(a[86]), .Z(n11943) );
  NANDN U12099 ( .A(n17739), .B(n11943), .Z(n11795) );
  NAND U12100 ( .A(n11796), .B(n11795), .Z(n11868) );
  XNOR U12101 ( .A(n11869), .B(n11868), .Z(n11870) );
  XOR U12102 ( .A(n11871), .B(n11870), .Z(n11877) );
  XOR U12103 ( .A(n11876), .B(n11877), .Z(n11883) );
  XOR U12104 ( .A(n11882), .B(n11883), .Z(n11895) );
  XNOR U12105 ( .A(n11894), .B(n11895), .Z(n11826) );
  XNOR U12106 ( .A(n11827), .B(n11826), .Z(n11828) );
  XOR U12107 ( .A(n11829), .B(n11828), .Z(n11947) );
  XNOR U12108 ( .A(n11946), .B(n11947), .Z(n11948) );
  XNOR U12109 ( .A(n11949), .B(n11948), .Z(n11822) );
  XOR U12110 ( .A(n11823), .B(n11822), .Z(n11815) );
  NANDN U12111 ( .A(n11798), .B(n11797), .Z(n11802) );
  NANDN U12112 ( .A(n11800), .B(n11799), .Z(n11801) );
  AND U12113 ( .A(n11802), .B(n11801), .Z(n11814) );
  XOR U12114 ( .A(n11815), .B(n11814), .Z(n11817) );
  XNOR U12115 ( .A(n11816), .B(n11817), .Z(n11808) );
  XNOR U12116 ( .A(n11809), .B(n11808), .Z(n11810) );
  XNOR U12117 ( .A(n11811), .B(n11810), .Z(n11952) );
  XNOR U12118 ( .A(sreg[190]), .B(n11952), .Z(n11954) );
  NANDN U12119 ( .A(sreg[189]), .B(n11803), .Z(n11807) );
  NAND U12120 ( .A(n11805), .B(n11804), .Z(n11806) );
  NAND U12121 ( .A(n11807), .B(n11806), .Z(n11953) );
  XNOR U12122 ( .A(n11954), .B(n11953), .Z(c[190]) );
  NANDN U12123 ( .A(n11809), .B(n11808), .Z(n11813) );
  NANDN U12124 ( .A(n11811), .B(n11810), .Z(n11812) );
  AND U12125 ( .A(n11813), .B(n11812), .Z(n11960) );
  NANDN U12126 ( .A(n11815), .B(n11814), .Z(n11819) );
  NANDN U12127 ( .A(n11817), .B(n11816), .Z(n11818) );
  AND U12128 ( .A(n11819), .B(n11818), .Z(n11958) );
  NANDN U12129 ( .A(n11821), .B(n11820), .Z(n11825) );
  NAND U12130 ( .A(n11823), .B(n11822), .Z(n11824) );
  AND U12131 ( .A(n11825), .B(n11824), .Z(n11965) );
  NANDN U12132 ( .A(n11827), .B(n11826), .Z(n11831) );
  NANDN U12133 ( .A(n11829), .B(n11828), .Z(n11830) );
  AND U12134 ( .A(n11831), .B(n11830), .Z(n11970) );
  NANDN U12135 ( .A(n11833), .B(n11832), .Z(n11837) );
  NAND U12136 ( .A(n11835), .B(n11834), .Z(n11836) );
  AND U12137 ( .A(n11837), .B(n11836), .Z(n11969) );
  XNOR U12138 ( .A(n11970), .B(n11969), .Z(n11972) );
  NANDN U12139 ( .A(n11839), .B(n11838), .Z(n11843) );
  NANDN U12140 ( .A(n11841), .B(n11840), .Z(n11842) );
  AND U12141 ( .A(n11843), .B(n11842), .Z(n12049) );
  NANDN U12142 ( .A(n19237), .B(n11844), .Z(n11846) );
  XOR U12143 ( .A(b[27]), .B(a[69]), .Z(n11993) );
  NANDN U12144 ( .A(n19277), .B(n11993), .Z(n11845) );
  AND U12145 ( .A(n11846), .B(n11845), .Z(n12056) );
  NANDN U12146 ( .A(n17072), .B(n11847), .Z(n11849) );
  XOR U12147 ( .A(b[5]), .B(a[91]), .Z(n11996) );
  NANDN U12148 ( .A(n17223), .B(n11996), .Z(n11848) );
  AND U12149 ( .A(n11849), .B(n11848), .Z(n12054) );
  NANDN U12150 ( .A(n18673), .B(n11850), .Z(n11852) );
  XOR U12151 ( .A(b[19]), .B(a[77]), .Z(n11999) );
  NANDN U12152 ( .A(n18758), .B(n11999), .Z(n11851) );
  NAND U12153 ( .A(n11852), .B(n11851), .Z(n12053) );
  XNOR U12154 ( .A(n12054), .B(n12053), .Z(n12055) );
  XNOR U12155 ( .A(n12056), .B(n12055), .Z(n12047) );
  NANDN U12156 ( .A(n19425), .B(n11853), .Z(n11855) );
  XOR U12157 ( .A(b[31]), .B(a[65]), .Z(n12002) );
  NANDN U12158 ( .A(n19426), .B(n12002), .Z(n11854) );
  AND U12159 ( .A(n11855), .B(n11854), .Z(n12014) );
  NANDN U12160 ( .A(n17067), .B(n11856), .Z(n11858) );
  XOR U12161 ( .A(b[3]), .B(a[93]), .Z(n12005) );
  NANDN U12162 ( .A(n17068), .B(n12005), .Z(n11857) );
  AND U12163 ( .A(n11858), .B(n11857), .Z(n12012) );
  NANDN U12164 ( .A(n18514), .B(n11859), .Z(n11861) );
  XOR U12165 ( .A(b[17]), .B(a[79]), .Z(n12008) );
  NANDN U12166 ( .A(n18585), .B(n12008), .Z(n11860) );
  NAND U12167 ( .A(n11861), .B(n11860), .Z(n12011) );
  XNOR U12168 ( .A(n12012), .B(n12011), .Z(n12013) );
  XOR U12169 ( .A(n12014), .B(n12013), .Z(n12048) );
  XOR U12170 ( .A(n12047), .B(n12048), .Z(n12050) );
  XOR U12171 ( .A(n12049), .B(n12050), .Z(n11982) );
  NANDN U12172 ( .A(n11863), .B(n11862), .Z(n11867) );
  NANDN U12173 ( .A(n11865), .B(n11864), .Z(n11866) );
  AND U12174 ( .A(n11867), .B(n11866), .Z(n12035) );
  NANDN U12175 ( .A(n11869), .B(n11868), .Z(n11873) );
  NANDN U12176 ( .A(n11871), .B(n11870), .Z(n11872) );
  NAND U12177 ( .A(n11873), .B(n11872), .Z(n12036) );
  XNOR U12178 ( .A(n12035), .B(n12036), .Z(n12037) );
  NANDN U12179 ( .A(n11875), .B(n11874), .Z(n11879) );
  NANDN U12180 ( .A(n11877), .B(n11876), .Z(n11878) );
  NAND U12181 ( .A(n11879), .B(n11878), .Z(n12038) );
  XNOR U12182 ( .A(n12037), .B(n12038), .Z(n11981) );
  XNOR U12183 ( .A(n11982), .B(n11981), .Z(n11984) );
  NANDN U12184 ( .A(n11881), .B(n11880), .Z(n11885) );
  NANDN U12185 ( .A(n11883), .B(n11882), .Z(n11884) );
  AND U12186 ( .A(n11885), .B(n11884), .Z(n11983) );
  XOR U12187 ( .A(n11984), .B(n11983), .Z(n12098) );
  NANDN U12188 ( .A(n11887), .B(n11886), .Z(n11891) );
  NANDN U12189 ( .A(n11889), .B(n11888), .Z(n11890) );
  AND U12190 ( .A(n11891), .B(n11890), .Z(n12095) );
  NANDN U12191 ( .A(n11893), .B(n11892), .Z(n11897) );
  NANDN U12192 ( .A(n11895), .B(n11894), .Z(n11896) );
  AND U12193 ( .A(n11897), .B(n11896), .Z(n11978) );
  NANDN U12194 ( .A(n11899), .B(n11898), .Z(n11903) );
  OR U12195 ( .A(n11901), .B(n11900), .Z(n11902) );
  AND U12196 ( .A(n11903), .B(n11902), .Z(n11976) );
  NANDN U12197 ( .A(n11905), .B(n11904), .Z(n11909) );
  NANDN U12198 ( .A(n11907), .B(n11906), .Z(n11908) );
  AND U12199 ( .A(n11909), .B(n11908), .Z(n12042) );
  NANDN U12200 ( .A(n11911), .B(n11910), .Z(n11915) );
  NANDN U12201 ( .A(n11913), .B(n11912), .Z(n11914) );
  NAND U12202 ( .A(n11915), .B(n11914), .Z(n12041) );
  XNOR U12203 ( .A(n12042), .B(n12041), .Z(n12043) );
  NAND U12204 ( .A(b[0]), .B(a[95]), .Z(n11916) );
  XNOR U12205 ( .A(b[1]), .B(n11916), .Z(n11918) );
  NANDN U12206 ( .A(b[0]), .B(a[94]), .Z(n11917) );
  NAND U12207 ( .A(n11918), .B(n11917), .Z(n11990) );
  NANDN U12208 ( .A(n19394), .B(n11919), .Z(n11921) );
  XOR U12209 ( .A(b[29]), .B(a[67]), .Z(n12065) );
  NANDN U12210 ( .A(n19395), .B(n12065), .Z(n11920) );
  AND U12211 ( .A(n11921), .B(n11920), .Z(n11988) );
  AND U12212 ( .A(b[31]), .B(a[63]), .Z(n11987) );
  XNOR U12213 ( .A(n11988), .B(n11987), .Z(n11989) );
  XNOR U12214 ( .A(n11990), .B(n11989), .Z(n12029) );
  NANDN U12215 ( .A(n19005), .B(n11922), .Z(n11924) );
  XOR U12216 ( .A(b[23]), .B(a[73]), .Z(n12071) );
  NANDN U12217 ( .A(n19055), .B(n12071), .Z(n11923) );
  AND U12218 ( .A(n11924), .B(n11923), .Z(n12062) );
  NANDN U12219 ( .A(n17362), .B(n11925), .Z(n11927) );
  XOR U12220 ( .A(b[7]), .B(a[89]), .Z(n12074) );
  NANDN U12221 ( .A(n17522), .B(n12074), .Z(n11926) );
  AND U12222 ( .A(n11927), .B(n11926), .Z(n12060) );
  NANDN U12223 ( .A(n19116), .B(n11928), .Z(n11930) );
  XOR U12224 ( .A(b[25]), .B(a[71]), .Z(n12077) );
  NANDN U12225 ( .A(n19179), .B(n12077), .Z(n11929) );
  NAND U12226 ( .A(n11930), .B(n11929), .Z(n12059) );
  XNOR U12227 ( .A(n12060), .B(n12059), .Z(n12061) );
  XOR U12228 ( .A(n12062), .B(n12061), .Z(n12030) );
  XNOR U12229 ( .A(n12029), .B(n12030), .Z(n12031) );
  NANDN U12230 ( .A(n18113), .B(n11931), .Z(n11933) );
  XOR U12231 ( .A(b[13]), .B(a[83]), .Z(n12080) );
  NANDN U12232 ( .A(n18229), .B(n12080), .Z(n11932) );
  AND U12233 ( .A(n11933), .B(n11932), .Z(n12024) );
  NANDN U12234 ( .A(n17888), .B(n11934), .Z(n11936) );
  XOR U12235 ( .A(b[11]), .B(a[85]), .Z(n12083) );
  NANDN U12236 ( .A(n18025), .B(n12083), .Z(n11935) );
  NAND U12237 ( .A(n11936), .B(n11935), .Z(n12023) );
  XNOR U12238 ( .A(n12024), .B(n12023), .Z(n12025) );
  NANDN U12239 ( .A(n18487), .B(n11937), .Z(n11939) );
  XOR U12240 ( .A(b[15]), .B(a[81]), .Z(n12086) );
  NANDN U12241 ( .A(n18311), .B(n12086), .Z(n11938) );
  AND U12242 ( .A(n11939), .B(n11938), .Z(n12020) );
  NANDN U12243 ( .A(n18853), .B(n11940), .Z(n11942) );
  XOR U12244 ( .A(b[21]), .B(a[75]), .Z(n12089) );
  NANDN U12245 ( .A(n18926), .B(n12089), .Z(n11941) );
  AND U12246 ( .A(n11942), .B(n11941), .Z(n12018) );
  NANDN U12247 ( .A(n17613), .B(n11943), .Z(n11945) );
  XOR U12248 ( .A(b[9]), .B(a[87]), .Z(n12092) );
  NANDN U12249 ( .A(n17739), .B(n12092), .Z(n11944) );
  NAND U12250 ( .A(n11945), .B(n11944), .Z(n12017) );
  XNOR U12251 ( .A(n12018), .B(n12017), .Z(n12019) );
  XOR U12252 ( .A(n12020), .B(n12019), .Z(n12026) );
  XOR U12253 ( .A(n12025), .B(n12026), .Z(n12032) );
  XOR U12254 ( .A(n12031), .B(n12032), .Z(n12044) );
  XNOR U12255 ( .A(n12043), .B(n12044), .Z(n11975) );
  XNOR U12256 ( .A(n11976), .B(n11975), .Z(n11977) );
  XOR U12257 ( .A(n11978), .B(n11977), .Z(n12096) );
  XNOR U12258 ( .A(n12095), .B(n12096), .Z(n12097) );
  XNOR U12259 ( .A(n12098), .B(n12097), .Z(n11971) );
  XOR U12260 ( .A(n11972), .B(n11971), .Z(n11964) );
  NANDN U12261 ( .A(n11947), .B(n11946), .Z(n11951) );
  NANDN U12262 ( .A(n11949), .B(n11948), .Z(n11950) );
  AND U12263 ( .A(n11951), .B(n11950), .Z(n11963) );
  XOR U12264 ( .A(n11964), .B(n11963), .Z(n11966) );
  XNOR U12265 ( .A(n11965), .B(n11966), .Z(n11957) );
  XNOR U12266 ( .A(n11958), .B(n11957), .Z(n11959) );
  XNOR U12267 ( .A(n11960), .B(n11959), .Z(n12101) );
  XNOR U12268 ( .A(sreg[191]), .B(n12101), .Z(n12103) );
  NANDN U12269 ( .A(sreg[190]), .B(n11952), .Z(n11956) );
  NAND U12270 ( .A(n11954), .B(n11953), .Z(n11955) );
  NAND U12271 ( .A(n11956), .B(n11955), .Z(n12102) );
  XNOR U12272 ( .A(n12103), .B(n12102), .Z(c[191]) );
  NANDN U12273 ( .A(n11958), .B(n11957), .Z(n11962) );
  NANDN U12274 ( .A(n11960), .B(n11959), .Z(n11961) );
  AND U12275 ( .A(n11962), .B(n11961), .Z(n12109) );
  NANDN U12276 ( .A(n11964), .B(n11963), .Z(n11968) );
  NANDN U12277 ( .A(n11966), .B(n11965), .Z(n11967) );
  AND U12278 ( .A(n11968), .B(n11967), .Z(n12107) );
  NANDN U12279 ( .A(n11970), .B(n11969), .Z(n11974) );
  NAND U12280 ( .A(n11972), .B(n11971), .Z(n11973) );
  AND U12281 ( .A(n11974), .B(n11973), .Z(n12114) );
  NANDN U12282 ( .A(n11976), .B(n11975), .Z(n11980) );
  NANDN U12283 ( .A(n11978), .B(n11977), .Z(n11979) );
  AND U12284 ( .A(n11980), .B(n11979), .Z(n12243) );
  NANDN U12285 ( .A(n11982), .B(n11981), .Z(n11986) );
  NAND U12286 ( .A(n11984), .B(n11983), .Z(n11985) );
  AND U12287 ( .A(n11986), .B(n11985), .Z(n12242) );
  XNOR U12288 ( .A(n12243), .B(n12242), .Z(n12245) );
  NANDN U12289 ( .A(n11988), .B(n11987), .Z(n11992) );
  NANDN U12290 ( .A(n11990), .B(n11989), .Z(n11991) );
  AND U12291 ( .A(n11992), .B(n11991), .Z(n12190) );
  NANDN U12292 ( .A(n19237), .B(n11993), .Z(n11995) );
  XOR U12293 ( .A(b[27]), .B(a[70]), .Z(n12136) );
  NANDN U12294 ( .A(n19277), .B(n12136), .Z(n11994) );
  AND U12295 ( .A(n11995), .B(n11994), .Z(n12197) );
  NANDN U12296 ( .A(n17072), .B(n11996), .Z(n11998) );
  XOR U12297 ( .A(b[5]), .B(a[92]), .Z(n12139) );
  NANDN U12298 ( .A(n17223), .B(n12139), .Z(n11997) );
  AND U12299 ( .A(n11998), .B(n11997), .Z(n12195) );
  NANDN U12300 ( .A(n18673), .B(n11999), .Z(n12001) );
  XOR U12301 ( .A(b[19]), .B(a[78]), .Z(n12142) );
  NANDN U12302 ( .A(n18758), .B(n12142), .Z(n12000) );
  NAND U12303 ( .A(n12001), .B(n12000), .Z(n12194) );
  XNOR U12304 ( .A(n12195), .B(n12194), .Z(n12196) );
  XNOR U12305 ( .A(n12197), .B(n12196), .Z(n12188) );
  NANDN U12306 ( .A(n19425), .B(n12002), .Z(n12004) );
  XOR U12307 ( .A(b[31]), .B(a[66]), .Z(n12145) );
  NANDN U12308 ( .A(n19426), .B(n12145), .Z(n12003) );
  AND U12309 ( .A(n12004), .B(n12003), .Z(n12157) );
  NANDN U12310 ( .A(n17067), .B(n12005), .Z(n12007) );
  XOR U12311 ( .A(b[3]), .B(a[94]), .Z(n12148) );
  NANDN U12312 ( .A(n17068), .B(n12148), .Z(n12006) );
  AND U12313 ( .A(n12007), .B(n12006), .Z(n12155) );
  NANDN U12314 ( .A(n18514), .B(n12008), .Z(n12010) );
  XOR U12315 ( .A(b[17]), .B(a[80]), .Z(n12151) );
  NANDN U12316 ( .A(n18585), .B(n12151), .Z(n12009) );
  NAND U12317 ( .A(n12010), .B(n12009), .Z(n12154) );
  XNOR U12318 ( .A(n12155), .B(n12154), .Z(n12156) );
  XOR U12319 ( .A(n12157), .B(n12156), .Z(n12189) );
  XOR U12320 ( .A(n12188), .B(n12189), .Z(n12191) );
  XOR U12321 ( .A(n12190), .B(n12191), .Z(n12125) );
  NANDN U12322 ( .A(n12012), .B(n12011), .Z(n12016) );
  NANDN U12323 ( .A(n12014), .B(n12013), .Z(n12015) );
  AND U12324 ( .A(n12016), .B(n12015), .Z(n12178) );
  NANDN U12325 ( .A(n12018), .B(n12017), .Z(n12022) );
  NANDN U12326 ( .A(n12020), .B(n12019), .Z(n12021) );
  NAND U12327 ( .A(n12022), .B(n12021), .Z(n12179) );
  XNOR U12328 ( .A(n12178), .B(n12179), .Z(n12180) );
  NANDN U12329 ( .A(n12024), .B(n12023), .Z(n12028) );
  NANDN U12330 ( .A(n12026), .B(n12025), .Z(n12027) );
  NAND U12331 ( .A(n12028), .B(n12027), .Z(n12181) );
  XNOR U12332 ( .A(n12180), .B(n12181), .Z(n12124) );
  XNOR U12333 ( .A(n12125), .B(n12124), .Z(n12127) );
  NANDN U12334 ( .A(n12030), .B(n12029), .Z(n12034) );
  NANDN U12335 ( .A(n12032), .B(n12031), .Z(n12033) );
  AND U12336 ( .A(n12034), .B(n12033), .Z(n12126) );
  XOR U12337 ( .A(n12127), .B(n12126), .Z(n12239) );
  NANDN U12338 ( .A(n12036), .B(n12035), .Z(n12040) );
  NANDN U12339 ( .A(n12038), .B(n12037), .Z(n12039) );
  AND U12340 ( .A(n12040), .B(n12039), .Z(n12236) );
  NANDN U12341 ( .A(n12042), .B(n12041), .Z(n12046) );
  NANDN U12342 ( .A(n12044), .B(n12043), .Z(n12045) );
  AND U12343 ( .A(n12046), .B(n12045), .Z(n12121) );
  NANDN U12344 ( .A(n12048), .B(n12047), .Z(n12052) );
  OR U12345 ( .A(n12050), .B(n12049), .Z(n12051) );
  AND U12346 ( .A(n12052), .B(n12051), .Z(n12119) );
  NANDN U12347 ( .A(n12054), .B(n12053), .Z(n12058) );
  NANDN U12348 ( .A(n12056), .B(n12055), .Z(n12057) );
  AND U12349 ( .A(n12058), .B(n12057), .Z(n12185) );
  NANDN U12350 ( .A(n12060), .B(n12059), .Z(n12064) );
  NANDN U12351 ( .A(n12062), .B(n12061), .Z(n12063) );
  NAND U12352 ( .A(n12064), .B(n12063), .Z(n12184) );
  XNOR U12353 ( .A(n12185), .B(n12184), .Z(n12187) );
  NANDN U12354 ( .A(n19394), .B(n12065), .Z(n12067) );
  XOR U12355 ( .A(b[29]), .B(a[68]), .Z(n12209) );
  NANDN U12356 ( .A(n19395), .B(n12209), .Z(n12066) );
  AND U12357 ( .A(n12067), .B(n12066), .Z(n12131) );
  AND U12358 ( .A(b[31]), .B(a[64]), .Z(n12130) );
  XNOR U12359 ( .A(n12131), .B(n12130), .Z(n12132) );
  NAND U12360 ( .A(b[0]), .B(a[96]), .Z(n12068) );
  XNOR U12361 ( .A(b[1]), .B(n12068), .Z(n12070) );
  NANDN U12362 ( .A(b[0]), .B(a[95]), .Z(n12069) );
  NAND U12363 ( .A(n12070), .B(n12069), .Z(n12133) );
  XNOR U12364 ( .A(n12132), .B(n12133), .Z(n12173) );
  NANDN U12365 ( .A(n19005), .B(n12071), .Z(n12073) );
  XOR U12366 ( .A(b[23]), .B(a[74]), .Z(n12212) );
  NANDN U12367 ( .A(n19055), .B(n12212), .Z(n12072) );
  AND U12368 ( .A(n12073), .B(n12072), .Z(n12202) );
  NANDN U12369 ( .A(n17362), .B(n12074), .Z(n12076) );
  XOR U12370 ( .A(b[7]), .B(a[90]), .Z(n12215) );
  NANDN U12371 ( .A(n17522), .B(n12215), .Z(n12075) );
  AND U12372 ( .A(n12076), .B(n12075), .Z(n12201) );
  NANDN U12373 ( .A(n19116), .B(n12077), .Z(n12079) );
  XOR U12374 ( .A(b[25]), .B(a[72]), .Z(n12218) );
  NANDN U12375 ( .A(n19179), .B(n12218), .Z(n12078) );
  NAND U12376 ( .A(n12079), .B(n12078), .Z(n12200) );
  XOR U12377 ( .A(n12201), .B(n12200), .Z(n12203) );
  XOR U12378 ( .A(n12202), .B(n12203), .Z(n12172) );
  XOR U12379 ( .A(n12173), .B(n12172), .Z(n12175) );
  NANDN U12380 ( .A(n18113), .B(n12080), .Z(n12082) );
  XOR U12381 ( .A(b[13]), .B(a[84]), .Z(n12221) );
  NANDN U12382 ( .A(n18229), .B(n12221), .Z(n12081) );
  AND U12383 ( .A(n12082), .B(n12081), .Z(n12167) );
  NANDN U12384 ( .A(n17888), .B(n12083), .Z(n12085) );
  XOR U12385 ( .A(b[11]), .B(a[86]), .Z(n12224) );
  NANDN U12386 ( .A(n18025), .B(n12224), .Z(n12084) );
  NAND U12387 ( .A(n12085), .B(n12084), .Z(n12166) );
  XNOR U12388 ( .A(n12167), .B(n12166), .Z(n12169) );
  NANDN U12389 ( .A(n18487), .B(n12086), .Z(n12088) );
  XOR U12390 ( .A(b[15]), .B(a[82]), .Z(n12227) );
  NANDN U12391 ( .A(n18311), .B(n12227), .Z(n12087) );
  AND U12392 ( .A(n12088), .B(n12087), .Z(n12163) );
  NANDN U12393 ( .A(n18853), .B(n12089), .Z(n12091) );
  XOR U12394 ( .A(b[21]), .B(a[76]), .Z(n12230) );
  NANDN U12395 ( .A(n18926), .B(n12230), .Z(n12090) );
  AND U12396 ( .A(n12091), .B(n12090), .Z(n12161) );
  NANDN U12397 ( .A(n17613), .B(n12092), .Z(n12094) );
  XOR U12398 ( .A(b[9]), .B(a[88]), .Z(n12233) );
  NANDN U12399 ( .A(n17739), .B(n12233), .Z(n12093) );
  NAND U12400 ( .A(n12094), .B(n12093), .Z(n12160) );
  XNOR U12401 ( .A(n12161), .B(n12160), .Z(n12162) );
  XNOR U12402 ( .A(n12163), .B(n12162), .Z(n12168) );
  XOR U12403 ( .A(n12169), .B(n12168), .Z(n12174) );
  XOR U12404 ( .A(n12175), .B(n12174), .Z(n12186) );
  XOR U12405 ( .A(n12187), .B(n12186), .Z(n12118) );
  XNOR U12406 ( .A(n12119), .B(n12118), .Z(n12120) );
  XOR U12407 ( .A(n12121), .B(n12120), .Z(n12237) );
  XNOR U12408 ( .A(n12236), .B(n12237), .Z(n12238) );
  XNOR U12409 ( .A(n12239), .B(n12238), .Z(n12244) );
  XOR U12410 ( .A(n12245), .B(n12244), .Z(n12113) );
  NANDN U12411 ( .A(n12096), .B(n12095), .Z(n12100) );
  NANDN U12412 ( .A(n12098), .B(n12097), .Z(n12099) );
  AND U12413 ( .A(n12100), .B(n12099), .Z(n12112) );
  XOR U12414 ( .A(n12113), .B(n12112), .Z(n12115) );
  XNOR U12415 ( .A(n12114), .B(n12115), .Z(n12106) );
  XNOR U12416 ( .A(n12107), .B(n12106), .Z(n12108) );
  XNOR U12417 ( .A(n12109), .B(n12108), .Z(n12248) );
  XNOR U12418 ( .A(sreg[192]), .B(n12248), .Z(n12250) );
  NANDN U12419 ( .A(sreg[191]), .B(n12101), .Z(n12105) );
  NAND U12420 ( .A(n12103), .B(n12102), .Z(n12104) );
  NAND U12421 ( .A(n12105), .B(n12104), .Z(n12249) );
  XNOR U12422 ( .A(n12250), .B(n12249), .Z(c[192]) );
  NANDN U12423 ( .A(n12107), .B(n12106), .Z(n12111) );
  NANDN U12424 ( .A(n12109), .B(n12108), .Z(n12110) );
  AND U12425 ( .A(n12111), .B(n12110), .Z(n12256) );
  NANDN U12426 ( .A(n12113), .B(n12112), .Z(n12117) );
  NANDN U12427 ( .A(n12115), .B(n12114), .Z(n12116) );
  AND U12428 ( .A(n12117), .B(n12116), .Z(n12254) );
  NANDN U12429 ( .A(n12119), .B(n12118), .Z(n12123) );
  NANDN U12430 ( .A(n12121), .B(n12120), .Z(n12122) );
  AND U12431 ( .A(n12123), .B(n12122), .Z(n12390) );
  NANDN U12432 ( .A(n12125), .B(n12124), .Z(n12129) );
  NAND U12433 ( .A(n12127), .B(n12126), .Z(n12128) );
  AND U12434 ( .A(n12129), .B(n12128), .Z(n12389) );
  XNOR U12435 ( .A(n12390), .B(n12389), .Z(n12392) );
  NANDN U12436 ( .A(n12131), .B(n12130), .Z(n12135) );
  NANDN U12437 ( .A(n12133), .B(n12132), .Z(n12134) );
  AND U12438 ( .A(n12135), .B(n12134), .Z(n12325) );
  NANDN U12439 ( .A(n19237), .B(n12136), .Z(n12138) );
  XOR U12440 ( .A(b[27]), .B(a[71]), .Z(n12271) );
  NANDN U12441 ( .A(n19277), .B(n12271), .Z(n12137) );
  AND U12442 ( .A(n12138), .B(n12137), .Z(n12332) );
  NANDN U12443 ( .A(n17072), .B(n12139), .Z(n12141) );
  XOR U12444 ( .A(b[5]), .B(a[93]), .Z(n12274) );
  NANDN U12445 ( .A(n17223), .B(n12274), .Z(n12140) );
  AND U12446 ( .A(n12141), .B(n12140), .Z(n12330) );
  NANDN U12447 ( .A(n18673), .B(n12142), .Z(n12144) );
  XOR U12448 ( .A(b[19]), .B(a[79]), .Z(n12277) );
  NANDN U12449 ( .A(n18758), .B(n12277), .Z(n12143) );
  NAND U12450 ( .A(n12144), .B(n12143), .Z(n12329) );
  XNOR U12451 ( .A(n12330), .B(n12329), .Z(n12331) );
  XNOR U12452 ( .A(n12332), .B(n12331), .Z(n12323) );
  NANDN U12453 ( .A(n19425), .B(n12145), .Z(n12147) );
  XOR U12454 ( .A(b[31]), .B(a[67]), .Z(n12280) );
  NANDN U12455 ( .A(n19426), .B(n12280), .Z(n12146) );
  AND U12456 ( .A(n12147), .B(n12146), .Z(n12292) );
  NANDN U12457 ( .A(n17067), .B(n12148), .Z(n12150) );
  XOR U12458 ( .A(b[3]), .B(a[95]), .Z(n12283) );
  NANDN U12459 ( .A(n17068), .B(n12283), .Z(n12149) );
  AND U12460 ( .A(n12150), .B(n12149), .Z(n12290) );
  NANDN U12461 ( .A(n18514), .B(n12151), .Z(n12153) );
  XOR U12462 ( .A(b[17]), .B(a[81]), .Z(n12286) );
  NANDN U12463 ( .A(n18585), .B(n12286), .Z(n12152) );
  NAND U12464 ( .A(n12153), .B(n12152), .Z(n12289) );
  XNOR U12465 ( .A(n12290), .B(n12289), .Z(n12291) );
  XOR U12466 ( .A(n12292), .B(n12291), .Z(n12324) );
  XOR U12467 ( .A(n12323), .B(n12324), .Z(n12326) );
  XOR U12468 ( .A(n12325), .B(n12326), .Z(n12372) );
  NANDN U12469 ( .A(n12155), .B(n12154), .Z(n12159) );
  NANDN U12470 ( .A(n12157), .B(n12156), .Z(n12158) );
  AND U12471 ( .A(n12159), .B(n12158), .Z(n12313) );
  NANDN U12472 ( .A(n12161), .B(n12160), .Z(n12165) );
  NANDN U12473 ( .A(n12163), .B(n12162), .Z(n12164) );
  NAND U12474 ( .A(n12165), .B(n12164), .Z(n12314) );
  XNOR U12475 ( .A(n12313), .B(n12314), .Z(n12315) );
  NANDN U12476 ( .A(n12167), .B(n12166), .Z(n12171) );
  NAND U12477 ( .A(n12169), .B(n12168), .Z(n12170) );
  NAND U12478 ( .A(n12171), .B(n12170), .Z(n12316) );
  XNOR U12479 ( .A(n12315), .B(n12316), .Z(n12371) );
  XNOR U12480 ( .A(n12372), .B(n12371), .Z(n12374) );
  NAND U12481 ( .A(n12173), .B(n12172), .Z(n12177) );
  NAND U12482 ( .A(n12175), .B(n12174), .Z(n12176) );
  AND U12483 ( .A(n12177), .B(n12176), .Z(n12373) );
  XOR U12484 ( .A(n12374), .B(n12373), .Z(n12386) );
  NANDN U12485 ( .A(n12179), .B(n12178), .Z(n12183) );
  NANDN U12486 ( .A(n12181), .B(n12180), .Z(n12182) );
  AND U12487 ( .A(n12183), .B(n12182), .Z(n12383) );
  NANDN U12488 ( .A(n12189), .B(n12188), .Z(n12193) );
  OR U12489 ( .A(n12191), .B(n12190), .Z(n12192) );
  AND U12490 ( .A(n12193), .B(n12192), .Z(n12378) );
  NANDN U12491 ( .A(n12195), .B(n12194), .Z(n12199) );
  NANDN U12492 ( .A(n12197), .B(n12196), .Z(n12198) );
  AND U12493 ( .A(n12199), .B(n12198), .Z(n12320) );
  NANDN U12494 ( .A(n12201), .B(n12200), .Z(n12205) );
  OR U12495 ( .A(n12203), .B(n12202), .Z(n12204) );
  NAND U12496 ( .A(n12205), .B(n12204), .Z(n12319) );
  XNOR U12497 ( .A(n12320), .B(n12319), .Z(n12322) );
  NAND U12498 ( .A(b[0]), .B(a[97]), .Z(n12206) );
  XNOR U12499 ( .A(b[1]), .B(n12206), .Z(n12208) );
  NANDN U12500 ( .A(b[0]), .B(a[96]), .Z(n12207) );
  NAND U12501 ( .A(n12208), .B(n12207), .Z(n12268) );
  NANDN U12502 ( .A(n19394), .B(n12209), .Z(n12211) );
  XOR U12503 ( .A(b[29]), .B(a[69]), .Z(n12344) );
  NANDN U12504 ( .A(n19395), .B(n12344), .Z(n12210) );
  AND U12505 ( .A(n12211), .B(n12210), .Z(n12266) );
  AND U12506 ( .A(b[31]), .B(a[65]), .Z(n12265) );
  XNOR U12507 ( .A(n12266), .B(n12265), .Z(n12267) );
  XNOR U12508 ( .A(n12268), .B(n12267), .Z(n12308) );
  NANDN U12509 ( .A(n19005), .B(n12212), .Z(n12214) );
  XOR U12510 ( .A(b[23]), .B(a[75]), .Z(n12347) );
  NANDN U12511 ( .A(n19055), .B(n12347), .Z(n12213) );
  AND U12512 ( .A(n12214), .B(n12213), .Z(n12337) );
  NANDN U12513 ( .A(n17362), .B(n12215), .Z(n12217) );
  XOR U12514 ( .A(b[7]), .B(a[91]), .Z(n12350) );
  NANDN U12515 ( .A(n17522), .B(n12350), .Z(n12216) );
  AND U12516 ( .A(n12217), .B(n12216), .Z(n12336) );
  NANDN U12517 ( .A(n19116), .B(n12218), .Z(n12220) );
  XOR U12518 ( .A(b[25]), .B(a[73]), .Z(n12353) );
  NANDN U12519 ( .A(n19179), .B(n12353), .Z(n12219) );
  NAND U12520 ( .A(n12220), .B(n12219), .Z(n12335) );
  XOR U12521 ( .A(n12336), .B(n12335), .Z(n12338) );
  XOR U12522 ( .A(n12337), .B(n12338), .Z(n12307) );
  XOR U12523 ( .A(n12308), .B(n12307), .Z(n12310) );
  NANDN U12524 ( .A(n18113), .B(n12221), .Z(n12223) );
  XOR U12525 ( .A(b[13]), .B(a[85]), .Z(n12356) );
  NANDN U12526 ( .A(n18229), .B(n12356), .Z(n12222) );
  AND U12527 ( .A(n12223), .B(n12222), .Z(n12302) );
  NANDN U12528 ( .A(n17888), .B(n12224), .Z(n12226) );
  XOR U12529 ( .A(b[11]), .B(a[87]), .Z(n12359) );
  NANDN U12530 ( .A(n18025), .B(n12359), .Z(n12225) );
  NAND U12531 ( .A(n12226), .B(n12225), .Z(n12301) );
  XNOR U12532 ( .A(n12302), .B(n12301), .Z(n12304) );
  NANDN U12533 ( .A(n18487), .B(n12227), .Z(n12229) );
  XOR U12534 ( .A(b[15]), .B(a[83]), .Z(n12362) );
  NANDN U12535 ( .A(n18311), .B(n12362), .Z(n12228) );
  AND U12536 ( .A(n12229), .B(n12228), .Z(n12298) );
  NANDN U12537 ( .A(n18853), .B(n12230), .Z(n12232) );
  XOR U12538 ( .A(b[21]), .B(a[77]), .Z(n12365) );
  NANDN U12539 ( .A(n18926), .B(n12365), .Z(n12231) );
  AND U12540 ( .A(n12232), .B(n12231), .Z(n12296) );
  NANDN U12541 ( .A(n17613), .B(n12233), .Z(n12235) );
  XOR U12542 ( .A(b[9]), .B(a[89]), .Z(n12368) );
  NANDN U12543 ( .A(n17739), .B(n12368), .Z(n12234) );
  NAND U12544 ( .A(n12235), .B(n12234), .Z(n12295) );
  XNOR U12545 ( .A(n12296), .B(n12295), .Z(n12297) );
  XNOR U12546 ( .A(n12298), .B(n12297), .Z(n12303) );
  XOR U12547 ( .A(n12304), .B(n12303), .Z(n12309) );
  XOR U12548 ( .A(n12310), .B(n12309), .Z(n12321) );
  XOR U12549 ( .A(n12322), .B(n12321), .Z(n12377) );
  XNOR U12550 ( .A(n12378), .B(n12377), .Z(n12379) );
  XOR U12551 ( .A(n12380), .B(n12379), .Z(n12384) );
  XNOR U12552 ( .A(n12383), .B(n12384), .Z(n12385) );
  XNOR U12553 ( .A(n12386), .B(n12385), .Z(n12391) );
  XOR U12554 ( .A(n12392), .B(n12391), .Z(n12260) );
  NANDN U12555 ( .A(n12237), .B(n12236), .Z(n12241) );
  NANDN U12556 ( .A(n12239), .B(n12238), .Z(n12240) );
  AND U12557 ( .A(n12241), .B(n12240), .Z(n12259) );
  XNOR U12558 ( .A(n12260), .B(n12259), .Z(n12261) );
  NANDN U12559 ( .A(n12243), .B(n12242), .Z(n12247) );
  NAND U12560 ( .A(n12245), .B(n12244), .Z(n12246) );
  NAND U12561 ( .A(n12247), .B(n12246), .Z(n12262) );
  XNOR U12562 ( .A(n12261), .B(n12262), .Z(n12253) );
  XNOR U12563 ( .A(n12254), .B(n12253), .Z(n12255) );
  XNOR U12564 ( .A(n12256), .B(n12255), .Z(n12395) );
  XNOR U12565 ( .A(sreg[193]), .B(n12395), .Z(n12397) );
  NANDN U12566 ( .A(sreg[192]), .B(n12248), .Z(n12252) );
  NAND U12567 ( .A(n12250), .B(n12249), .Z(n12251) );
  NAND U12568 ( .A(n12252), .B(n12251), .Z(n12396) );
  XNOR U12569 ( .A(n12397), .B(n12396), .Z(c[193]) );
  NANDN U12570 ( .A(n12254), .B(n12253), .Z(n12258) );
  NANDN U12571 ( .A(n12256), .B(n12255), .Z(n12257) );
  AND U12572 ( .A(n12258), .B(n12257), .Z(n12403) );
  NANDN U12573 ( .A(n12260), .B(n12259), .Z(n12264) );
  NANDN U12574 ( .A(n12262), .B(n12261), .Z(n12263) );
  AND U12575 ( .A(n12264), .B(n12263), .Z(n12401) );
  NANDN U12576 ( .A(n12266), .B(n12265), .Z(n12270) );
  NANDN U12577 ( .A(n12268), .B(n12267), .Z(n12269) );
  AND U12578 ( .A(n12270), .B(n12269), .Z(n12480) );
  NANDN U12579 ( .A(n19237), .B(n12271), .Z(n12273) );
  XOR U12580 ( .A(b[27]), .B(a[72]), .Z(n12424) );
  NANDN U12581 ( .A(n19277), .B(n12424), .Z(n12272) );
  AND U12582 ( .A(n12273), .B(n12272), .Z(n12487) );
  NANDN U12583 ( .A(n17072), .B(n12274), .Z(n12276) );
  XOR U12584 ( .A(b[5]), .B(a[94]), .Z(n12427) );
  NANDN U12585 ( .A(n17223), .B(n12427), .Z(n12275) );
  AND U12586 ( .A(n12276), .B(n12275), .Z(n12485) );
  NANDN U12587 ( .A(n18673), .B(n12277), .Z(n12279) );
  XOR U12588 ( .A(b[19]), .B(a[80]), .Z(n12430) );
  NANDN U12589 ( .A(n18758), .B(n12430), .Z(n12278) );
  NAND U12590 ( .A(n12279), .B(n12278), .Z(n12484) );
  XNOR U12591 ( .A(n12485), .B(n12484), .Z(n12486) );
  XNOR U12592 ( .A(n12487), .B(n12486), .Z(n12478) );
  NANDN U12593 ( .A(n19425), .B(n12280), .Z(n12282) );
  XOR U12594 ( .A(b[31]), .B(a[68]), .Z(n12433) );
  NANDN U12595 ( .A(n19426), .B(n12433), .Z(n12281) );
  AND U12596 ( .A(n12282), .B(n12281), .Z(n12445) );
  NANDN U12597 ( .A(n17067), .B(n12283), .Z(n12285) );
  XOR U12598 ( .A(b[3]), .B(a[96]), .Z(n12436) );
  NANDN U12599 ( .A(n17068), .B(n12436), .Z(n12284) );
  AND U12600 ( .A(n12285), .B(n12284), .Z(n12443) );
  NANDN U12601 ( .A(n18514), .B(n12286), .Z(n12288) );
  XOR U12602 ( .A(b[17]), .B(a[82]), .Z(n12439) );
  NANDN U12603 ( .A(n18585), .B(n12439), .Z(n12287) );
  NAND U12604 ( .A(n12288), .B(n12287), .Z(n12442) );
  XNOR U12605 ( .A(n12443), .B(n12442), .Z(n12444) );
  XOR U12606 ( .A(n12445), .B(n12444), .Z(n12479) );
  XOR U12607 ( .A(n12478), .B(n12479), .Z(n12481) );
  XOR U12608 ( .A(n12480), .B(n12481), .Z(n12527) );
  NANDN U12609 ( .A(n12290), .B(n12289), .Z(n12294) );
  NANDN U12610 ( .A(n12292), .B(n12291), .Z(n12293) );
  AND U12611 ( .A(n12294), .B(n12293), .Z(n12466) );
  NANDN U12612 ( .A(n12296), .B(n12295), .Z(n12300) );
  NANDN U12613 ( .A(n12298), .B(n12297), .Z(n12299) );
  NAND U12614 ( .A(n12300), .B(n12299), .Z(n12467) );
  XNOR U12615 ( .A(n12466), .B(n12467), .Z(n12468) );
  NANDN U12616 ( .A(n12302), .B(n12301), .Z(n12306) );
  NAND U12617 ( .A(n12304), .B(n12303), .Z(n12305) );
  NAND U12618 ( .A(n12306), .B(n12305), .Z(n12469) );
  XNOR U12619 ( .A(n12468), .B(n12469), .Z(n12526) );
  XNOR U12620 ( .A(n12527), .B(n12526), .Z(n12529) );
  NAND U12621 ( .A(n12308), .B(n12307), .Z(n12312) );
  NAND U12622 ( .A(n12310), .B(n12309), .Z(n12311) );
  AND U12623 ( .A(n12312), .B(n12311), .Z(n12528) );
  XOR U12624 ( .A(n12529), .B(n12528), .Z(n12540) );
  NANDN U12625 ( .A(n12314), .B(n12313), .Z(n12318) );
  NANDN U12626 ( .A(n12316), .B(n12315), .Z(n12317) );
  AND U12627 ( .A(n12318), .B(n12317), .Z(n12538) );
  NANDN U12628 ( .A(n12324), .B(n12323), .Z(n12328) );
  OR U12629 ( .A(n12326), .B(n12325), .Z(n12327) );
  AND U12630 ( .A(n12328), .B(n12327), .Z(n12533) );
  NANDN U12631 ( .A(n12330), .B(n12329), .Z(n12334) );
  NANDN U12632 ( .A(n12332), .B(n12331), .Z(n12333) );
  AND U12633 ( .A(n12334), .B(n12333), .Z(n12473) );
  NANDN U12634 ( .A(n12336), .B(n12335), .Z(n12340) );
  OR U12635 ( .A(n12338), .B(n12337), .Z(n12339) );
  NAND U12636 ( .A(n12340), .B(n12339), .Z(n12472) );
  XNOR U12637 ( .A(n12473), .B(n12472), .Z(n12474) );
  NAND U12638 ( .A(b[0]), .B(a[98]), .Z(n12341) );
  XNOR U12639 ( .A(b[1]), .B(n12341), .Z(n12343) );
  NANDN U12640 ( .A(b[0]), .B(a[97]), .Z(n12342) );
  NAND U12641 ( .A(n12343), .B(n12342), .Z(n12421) );
  NANDN U12642 ( .A(n19394), .B(n12344), .Z(n12346) );
  XOR U12643 ( .A(b[29]), .B(a[70]), .Z(n12496) );
  NANDN U12644 ( .A(n19395), .B(n12496), .Z(n12345) );
  AND U12645 ( .A(n12346), .B(n12345), .Z(n12419) );
  AND U12646 ( .A(b[31]), .B(a[66]), .Z(n12418) );
  XNOR U12647 ( .A(n12419), .B(n12418), .Z(n12420) );
  XNOR U12648 ( .A(n12421), .B(n12420), .Z(n12460) );
  NANDN U12649 ( .A(n19005), .B(n12347), .Z(n12349) );
  XOR U12650 ( .A(b[23]), .B(a[76]), .Z(n12502) );
  NANDN U12651 ( .A(n19055), .B(n12502), .Z(n12348) );
  AND U12652 ( .A(n12349), .B(n12348), .Z(n12493) );
  NANDN U12653 ( .A(n17362), .B(n12350), .Z(n12352) );
  XOR U12654 ( .A(b[7]), .B(a[92]), .Z(n12505) );
  NANDN U12655 ( .A(n17522), .B(n12505), .Z(n12351) );
  AND U12656 ( .A(n12352), .B(n12351), .Z(n12491) );
  NANDN U12657 ( .A(n19116), .B(n12353), .Z(n12355) );
  XOR U12658 ( .A(b[25]), .B(a[74]), .Z(n12508) );
  NANDN U12659 ( .A(n19179), .B(n12508), .Z(n12354) );
  NAND U12660 ( .A(n12355), .B(n12354), .Z(n12490) );
  XNOR U12661 ( .A(n12491), .B(n12490), .Z(n12492) );
  XOR U12662 ( .A(n12493), .B(n12492), .Z(n12461) );
  XNOR U12663 ( .A(n12460), .B(n12461), .Z(n12462) );
  NANDN U12664 ( .A(n18113), .B(n12356), .Z(n12358) );
  XOR U12665 ( .A(b[13]), .B(a[86]), .Z(n12511) );
  NANDN U12666 ( .A(n18229), .B(n12511), .Z(n12357) );
  AND U12667 ( .A(n12358), .B(n12357), .Z(n12455) );
  NANDN U12668 ( .A(n17888), .B(n12359), .Z(n12361) );
  XOR U12669 ( .A(b[11]), .B(a[88]), .Z(n12514) );
  NANDN U12670 ( .A(n18025), .B(n12514), .Z(n12360) );
  NAND U12671 ( .A(n12361), .B(n12360), .Z(n12454) );
  XNOR U12672 ( .A(n12455), .B(n12454), .Z(n12456) );
  NANDN U12673 ( .A(n18487), .B(n12362), .Z(n12364) );
  XOR U12674 ( .A(b[15]), .B(a[84]), .Z(n12517) );
  NANDN U12675 ( .A(n18311), .B(n12517), .Z(n12363) );
  AND U12676 ( .A(n12364), .B(n12363), .Z(n12451) );
  NANDN U12677 ( .A(n18853), .B(n12365), .Z(n12367) );
  XOR U12678 ( .A(b[21]), .B(a[78]), .Z(n12520) );
  NANDN U12679 ( .A(n18926), .B(n12520), .Z(n12366) );
  AND U12680 ( .A(n12367), .B(n12366), .Z(n12449) );
  NANDN U12681 ( .A(n17613), .B(n12368), .Z(n12370) );
  XOR U12682 ( .A(b[9]), .B(a[90]), .Z(n12523) );
  NANDN U12683 ( .A(n17739), .B(n12523), .Z(n12369) );
  NAND U12684 ( .A(n12370), .B(n12369), .Z(n12448) );
  XNOR U12685 ( .A(n12449), .B(n12448), .Z(n12450) );
  XOR U12686 ( .A(n12451), .B(n12450), .Z(n12457) );
  XOR U12687 ( .A(n12456), .B(n12457), .Z(n12463) );
  XOR U12688 ( .A(n12462), .B(n12463), .Z(n12475) );
  XNOR U12689 ( .A(n12474), .B(n12475), .Z(n12532) );
  XNOR U12690 ( .A(n12533), .B(n12532), .Z(n12534) );
  XOR U12691 ( .A(n12535), .B(n12534), .Z(n12539) );
  XOR U12692 ( .A(n12538), .B(n12539), .Z(n12541) );
  XOR U12693 ( .A(n12540), .B(n12541), .Z(n12415) );
  NANDN U12694 ( .A(n12372), .B(n12371), .Z(n12376) );
  NAND U12695 ( .A(n12374), .B(n12373), .Z(n12375) );
  AND U12696 ( .A(n12376), .B(n12375), .Z(n12413) );
  NANDN U12697 ( .A(n12378), .B(n12377), .Z(n12382) );
  NANDN U12698 ( .A(n12380), .B(n12379), .Z(n12381) );
  AND U12699 ( .A(n12382), .B(n12381), .Z(n12412) );
  XNOR U12700 ( .A(n12413), .B(n12412), .Z(n12414) );
  XNOR U12701 ( .A(n12415), .B(n12414), .Z(n12406) );
  NANDN U12702 ( .A(n12384), .B(n12383), .Z(n12388) );
  NANDN U12703 ( .A(n12386), .B(n12385), .Z(n12387) );
  NAND U12704 ( .A(n12388), .B(n12387), .Z(n12407) );
  XNOR U12705 ( .A(n12406), .B(n12407), .Z(n12408) );
  NANDN U12706 ( .A(n12390), .B(n12389), .Z(n12394) );
  NAND U12707 ( .A(n12392), .B(n12391), .Z(n12393) );
  NAND U12708 ( .A(n12394), .B(n12393), .Z(n12409) );
  XNOR U12709 ( .A(n12408), .B(n12409), .Z(n12400) );
  XNOR U12710 ( .A(n12401), .B(n12400), .Z(n12402) );
  XNOR U12711 ( .A(n12403), .B(n12402), .Z(n12544) );
  XNOR U12712 ( .A(sreg[194]), .B(n12544), .Z(n12546) );
  NANDN U12713 ( .A(sreg[193]), .B(n12395), .Z(n12399) );
  NAND U12714 ( .A(n12397), .B(n12396), .Z(n12398) );
  NAND U12715 ( .A(n12399), .B(n12398), .Z(n12545) );
  XNOR U12716 ( .A(n12546), .B(n12545), .Z(c[194]) );
  NANDN U12717 ( .A(n12401), .B(n12400), .Z(n12405) );
  NANDN U12718 ( .A(n12403), .B(n12402), .Z(n12404) );
  AND U12719 ( .A(n12405), .B(n12404), .Z(n12552) );
  NANDN U12720 ( .A(n12407), .B(n12406), .Z(n12411) );
  NANDN U12721 ( .A(n12409), .B(n12408), .Z(n12410) );
  AND U12722 ( .A(n12411), .B(n12410), .Z(n12550) );
  NANDN U12723 ( .A(n12413), .B(n12412), .Z(n12417) );
  NANDN U12724 ( .A(n12415), .B(n12414), .Z(n12416) );
  AND U12725 ( .A(n12417), .B(n12416), .Z(n12558) );
  NANDN U12726 ( .A(n12419), .B(n12418), .Z(n12423) );
  NANDN U12727 ( .A(n12421), .B(n12420), .Z(n12422) );
  AND U12728 ( .A(n12423), .B(n12422), .Z(n12641) );
  NANDN U12729 ( .A(n19237), .B(n12424), .Z(n12426) );
  XOR U12730 ( .A(b[27]), .B(a[73]), .Z(n12585) );
  NANDN U12731 ( .A(n19277), .B(n12585), .Z(n12425) );
  AND U12732 ( .A(n12426), .B(n12425), .Z(n12648) );
  NANDN U12733 ( .A(n17072), .B(n12427), .Z(n12429) );
  XOR U12734 ( .A(b[5]), .B(a[95]), .Z(n12588) );
  NANDN U12735 ( .A(n17223), .B(n12588), .Z(n12428) );
  AND U12736 ( .A(n12429), .B(n12428), .Z(n12646) );
  NANDN U12737 ( .A(n18673), .B(n12430), .Z(n12432) );
  XOR U12738 ( .A(b[19]), .B(a[81]), .Z(n12591) );
  NANDN U12739 ( .A(n18758), .B(n12591), .Z(n12431) );
  NAND U12740 ( .A(n12432), .B(n12431), .Z(n12645) );
  XNOR U12741 ( .A(n12646), .B(n12645), .Z(n12647) );
  XNOR U12742 ( .A(n12648), .B(n12647), .Z(n12639) );
  NANDN U12743 ( .A(n19425), .B(n12433), .Z(n12435) );
  XOR U12744 ( .A(b[31]), .B(a[69]), .Z(n12594) );
  NANDN U12745 ( .A(n19426), .B(n12594), .Z(n12434) );
  AND U12746 ( .A(n12435), .B(n12434), .Z(n12606) );
  NANDN U12747 ( .A(n17067), .B(n12436), .Z(n12438) );
  XOR U12748 ( .A(b[3]), .B(a[97]), .Z(n12597) );
  NANDN U12749 ( .A(n17068), .B(n12597), .Z(n12437) );
  AND U12750 ( .A(n12438), .B(n12437), .Z(n12604) );
  NANDN U12751 ( .A(n18514), .B(n12439), .Z(n12441) );
  XOR U12752 ( .A(b[17]), .B(a[83]), .Z(n12600) );
  NANDN U12753 ( .A(n18585), .B(n12600), .Z(n12440) );
  NAND U12754 ( .A(n12441), .B(n12440), .Z(n12603) );
  XNOR U12755 ( .A(n12604), .B(n12603), .Z(n12605) );
  XOR U12756 ( .A(n12606), .B(n12605), .Z(n12640) );
  XOR U12757 ( .A(n12639), .B(n12640), .Z(n12642) );
  XOR U12758 ( .A(n12641), .B(n12642), .Z(n12574) );
  NANDN U12759 ( .A(n12443), .B(n12442), .Z(n12447) );
  NANDN U12760 ( .A(n12445), .B(n12444), .Z(n12446) );
  AND U12761 ( .A(n12447), .B(n12446), .Z(n12627) );
  NANDN U12762 ( .A(n12449), .B(n12448), .Z(n12453) );
  NANDN U12763 ( .A(n12451), .B(n12450), .Z(n12452) );
  NAND U12764 ( .A(n12453), .B(n12452), .Z(n12628) );
  XNOR U12765 ( .A(n12627), .B(n12628), .Z(n12629) );
  NANDN U12766 ( .A(n12455), .B(n12454), .Z(n12459) );
  NANDN U12767 ( .A(n12457), .B(n12456), .Z(n12458) );
  NAND U12768 ( .A(n12459), .B(n12458), .Z(n12630) );
  XNOR U12769 ( .A(n12629), .B(n12630), .Z(n12573) );
  XNOR U12770 ( .A(n12574), .B(n12573), .Z(n12576) );
  NANDN U12771 ( .A(n12461), .B(n12460), .Z(n12465) );
  NANDN U12772 ( .A(n12463), .B(n12462), .Z(n12464) );
  AND U12773 ( .A(n12465), .B(n12464), .Z(n12575) );
  XOR U12774 ( .A(n12576), .B(n12575), .Z(n12689) );
  NANDN U12775 ( .A(n12467), .B(n12466), .Z(n12471) );
  NANDN U12776 ( .A(n12469), .B(n12468), .Z(n12470) );
  AND U12777 ( .A(n12471), .B(n12470), .Z(n12687) );
  NANDN U12778 ( .A(n12473), .B(n12472), .Z(n12477) );
  NANDN U12779 ( .A(n12475), .B(n12474), .Z(n12476) );
  AND U12780 ( .A(n12477), .B(n12476), .Z(n12570) );
  NANDN U12781 ( .A(n12479), .B(n12478), .Z(n12483) );
  OR U12782 ( .A(n12481), .B(n12480), .Z(n12482) );
  AND U12783 ( .A(n12483), .B(n12482), .Z(n12568) );
  NANDN U12784 ( .A(n12485), .B(n12484), .Z(n12489) );
  NANDN U12785 ( .A(n12487), .B(n12486), .Z(n12488) );
  AND U12786 ( .A(n12489), .B(n12488), .Z(n12634) );
  NANDN U12787 ( .A(n12491), .B(n12490), .Z(n12495) );
  NANDN U12788 ( .A(n12493), .B(n12492), .Z(n12494) );
  NAND U12789 ( .A(n12495), .B(n12494), .Z(n12633) );
  XNOR U12790 ( .A(n12634), .B(n12633), .Z(n12635) );
  NANDN U12791 ( .A(n19394), .B(n12496), .Z(n12498) );
  XOR U12792 ( .A(b[29]), .B(a[71]), .Z(n12660) );
  NANDN U12793 ( .A(n19395), .B(n12660), .Z(n12497) );
  AND U12794 ( .A(n12498), .B(n12497), .Z(n12580) );
  AND U12795 ( .A(b[31]), .B(a[67]), .Z(n12579) );
  XNOR U12796 ( .A(n12580), .B(n12579), .Z(n12581) );
  NAND U12797 ( .A(b[0]), .B(a[99]), .Z(n12499) );
  XNOR U12798 ( .A(b[1]), .B(n12499), .Z(n12501) );
  NANDN U12799 ( .A(b[0]), .B(a[98]), .Z(n12500) );
  NAND U12800 ( .A(n12501), .B(n12500), .Z(n12582) );
  XNOR U12801 ( .A(n12581), .B(n12582), .Z(n12621) );
  NANDN U12802 ( .A(n19005), .B(n12502), .Z(n12504) );
  XOR U12803 ( .A(b[23]), .B(a[77]), .Z(n12663) );
  NANDN U12804 ( .A(n19055), .B(n12663), .Z(n12503) );
  AND U12805 ( .A(n12504), .B(n12503), .Z(n12654) );
  NANDN U12806 ( .A(n17362), .B(n12505), .Z(n12507) );
  XOR U12807 ( .A(b[7]), .B(a[93]), .Z(n12666) );
  NANDN U12808 ( .A(n17522), .B(n12666), .Z(n12506) );
  AND U12809 ( .A(n12507), .B(n12506), .Z(n12652) );
  NANDN U12810 ( .A(n19116), .B(n12508), .Z(n12510) );
  XOR U12811 ( .A(b[25]), .B(a[75]), .Z(n12669) );
  NANDN U12812 ( .A(n19179), .B(n12669), .Z(n12509) );
  NAND U12813 ( .A(n12510), .B(n12509), .Z(n12651) );
  XNOR U12814 ( .A(n12652), .B(n12651), .Z(n12653) );
  XOR U12815 ( .A(n12654), .B(n12653), .Z(n12622) );
  XNOR U12816 ( .A(n12621), .B(n12622), .Z(n12623) );
  NANDN U12817 ( .A(n18113), .B(n12511), .Z(n12513) );
  XOR U12818 ( .A(b[13]), .B(a[87]), .Z(n12672) );
  NANDN U12819 ( .A(n18229), .B(n12672), .Z(n12512) );
  AND U12820 ( .A(n12513), .B(n12512), .Z(n12616) );
  NANDN U12821 ( .A(n17888), .B(n12514), .Z(n12516) );
  XOR U12822 ( .A(b[11]), .B(a[89]), .Z(n12675) );
  NANDN U12823 ( .A(n18025), .B(n12675), .Z(n12515) );
  NAND U12824 ( .A(n12516), .B(n12515), .Z(n12615) );
  XNOR U12825 ( .A(n12616), .B(n12615), .Z(n12617) );
  NANDN U12826 ( .A(n18487), .B(n12517), .Z(n12519) );
  XOR U12827 ( .A(b[15]), .B(a[85]), .Z(n12678) );
  NANDN U12828 ( .A(n18311), .B(n12678), .Z(n12518) );
  AND U12829 ( .A(n12519), .B(n12518), .Z(n12612) );
  NANDN U12830 ( .A(n18853), .B(n12520), .Z(n12522) );
  XOR U12831 ( .A(b[21]), .B(a[79]), .Z(n12681) );
  NANDN U12832 ( .A(n18926), .B(n12681), .Z(n12521) );
  AND U12833 ( .A(n12522), .B(n12521), .Z(n12610) );
  NANDN U12834 ( .A(n17613), .B(n12523), .Z(n12525) );
  XOR U12835 ( .A(b[9]), .B(a[91]), .Z(n12684) );
  NANDN U12836 ( .A(n17739), .B(n12684), .Z(n12524) );
  NAND U12837 ( .A(n12525), .B(n12524), .Z(n12609) );
  XNOR U12838 ( .A(n12610), .B(n12609), .Z(n12611) );
  XOR U12839 ( .A(n12612), .B(n12611), .Z(n12618) );
  XOR U12840 ( .A(n12617), .B(n12618), .Z(n12624) );
  XOR U12841 ( .A(n12623), .B(n12624), .Z(n12636) );
  XNOR U12842 ( .A(n12635), .B(n12636), .Z(n12567) );
  XNOR U12843 ( .A(n12568), .B(n12567), .Z(n12569) );
  XOR U12844 ( .A(n12570), .B(n12569), .Z(n12688) );
  XOR U12845 ( .A(n12687), .B(n12688), .Z(n12690) );
  XOR U12846 ( .A(n12689), .B(n12690), .Z(n12564) );
  NANDN U12847 ( .A(n12527), .B(n12526), .Z(n12531) );
  NAND U12848 ( .A(n12529), .B(n12528), .Z(n12530) );
  AND U12849 ( .A(n12531), .B(n12530), .Z(n12562) );
  NANDN U12850 ( .A(n12533), .B(n12532), .Z(n12537) );
  NANDN U12851 ( .A(n12535), .B(n12534), .Z(n12536) );
  AND U12852 ( .A(n12537), .B(n12536), .Z(n12561) );
  XNOR U12853 ( .A(n12562), .B(n12561), .Z(n12563) );
  XNOR U12854 ( .A(n12564), .B(n12563), .Z(n12555) );
  NANDN U12855 ( .A(n12539), .B(n12538), .Z(n12543) );
  OR U12856 ( .A(n12541), .B(n12540), .Z(n12542) );
  NAND U12857 ( .A(n12543), .B(n12542), .Z(n12556) );
  XNOR U12858 ( .A(n12555), .B(n12556), .Z(n12557) );
  XNOR U12859 ( .A(n12558), .B(n12557), .Z(n12549) );
  XNOR U12860 ( .A(n12550), .B(n12549), .Z(n12551) );
  XNOR U12861 ( .A(n12552), .B(n12551), .Z(n12693) );
  XNOR U12862 ( .A(sreg[195]), .B(n12693), .Z(n12695) );
  NANDN U12863 ( .A(sreg[194]), .B(n12544), .Z(n12548) );
  NAND U12864 ( .A(n12546), .B(n12545), .Z(n12547) );
  NAND U12865 ( .A(n12548), .B(n12547), .Z(n12694) );
  XNOR U12866 ( .A(n12695), .B(n12694), .Z(c[195]) );
  NANDN U12867 ( .A(n12550), .B(n12549), .Z(n12554) );
  NANDN U12868 ( .A(n12552), .B(n12551), .Z(n12553) );
  AND U12869 ( .A(n12554), .B(n12553), .Z(n12701) );
  NANDN U12870 ( .A(n12556), .B(n12555), .Z(n12560) );
  NANDN U12871 ( .A(n12558), .B(n12557), .Z(n12559) );
  AND U12872 ( .A(n12560), .B(n12559), .Z(n12699) );
  NANDN U12873 ( .A(n12562), .B(n12561), .Z(n12566) );
  NANDN U12874 ( .A(n12564), .B(n12563), .Z(n12565) );
  AND U12875 ( .A(n12566), .B(n12565), .Z(n12707) );
  NANDN U12876 ( .A(n12568), .B(n12567), .Z(n12572) );
  NANDN U12877 ( .A(n12570), .B(n12569), .Z(n12571) );
  AND U12878 ( .A(n12572), .B(n12571), .Z(n12711) );
  NANDN U12879 ( .A(n12574), .B(n12573), .Z(n12578) );
  NAND U12880 ( .A(n12576), .B(n12575), .Z(n12577) );
  AND U12881 ( .A(n12578), .B(n12577), .Z(n12710) );
  XNOR U12882 ( .A(n12711), .B(n12710), .Z(n12713) );
  NANDN U12883 ( .A(n12580), .B(n12579), .Z(n12584) );
  NANDN U12884 ( .A(n12582), .B(n12581), .Z(n12583) );
  AND U12885 ( .A(n12584), .B(n12583), .Z(n12788) );
  NANDN U12886 ( .A(n19237), .B(n12585), .Z(n12587) );
  XOR U12887 ( .A(b[27]), .B(a[74]), .Z(n12734) );
  NANDN U12888 ( .A(n19277), .B(n12734), .Z(n12586) );
  AND U12889 ( .A(n12587), .B(n12586), .Z(n12795) );
  NANDN U12890 ( .A(n17072), .B(n12588), .Z(n12590) );
  XOR U12891 ( .A(b[5]), .B(a[96]), .Z(n12737) );
  NANDN U12892 ( .A(n17223), .B(n12737), .Z(n12589) );
  AND U12893 ( .A(n12590), .B(n12589), .Z(n12793) );
  NANDN U12894 ( .A(n18673), .B(n12591), .Z(n12593) );
  XOR U12895 ( .A(b[19]), .B(a[82]), .Z(n12740) );
  NANDN U12896 ( .A(n18758), .B(n12740), .Z(n12592) );
  NAND U12897 ( .A(n12593), .B(n12592), .Z(n12792) );
  XNOR U12898 ( .A(n12793), .B(n12792), .Z(n12794) );
  XNOR U12899 ( .A(n12795), .B(n12794), .Z(n12786) );
  NANDN U12900 ( .A(n19425), .B(n12594), .Z(n12596) );
  XOR U12901 ( .A(b[31]), .B(a[70]), .Z(n12743) );
  NANDN U12902 ( .A(n19426), .B(n12743), .Z(n12595) );
  AND U12903 ( .A(n12596), .B(n12595), .Z(n12755) );
  NANDN U12904 ( .A(n17067), .B(n12597), .Z(n12599) );
  XOR U12905 ( .A(b[3]), .B(a[98]), .Z(n12746) );
  NANDN U12906 ( .A(n17068), .B(n12746), .Z(n12598) );
  AND U12907 ( .A(n12599), .B(n12598), .Z(n12753) );
  NANDN U12908 ( .A(n18514), .B(n12600), .Z(n12602) );
  XOR U12909 ( .A(b[17]), .B(a[84]), .Z(n12749) );
  NANDN U12910 ( .A(n18585), .B(n12749), .Z(n12601) );
  NAND U12911 ( .A(n12602), .B(n12601), .Z(n12752) );
  XNOR U12912 ( .A(n12753), .B(n12752), .Z(n12754) );
  XOR U12913 ( .A(n12755), .B(n12754), .Z(n12787) );
  XOR U12914 ( .A(n12786), .B(n12787), .Z(n12789) );
  XOR U12915 ( .A(n12788), .B(n12789), .Z(n12723) );
  NANDN U12916 ( .A(n12604), .B(n12603), .Z(n12608) );
  NANDN U12917 ( .A(n12606), .B(n12605), .Z(n12607) );
  AND U12918 ( .A(n12608), .B(n12607), .Z(n12776) );
  NANDN U12919 ( .A(n12610), .B(n12609), .Z(n12614) );
  NANDN U12920 ( .A(n12612), .B(n12611), .Z(n12613) );
  NAND U12921 ( .A(n12614), .B(n12613), .Z(n12777) );
  XNOR U12922 ( .A(n12776), .B(n12777), .Z(n12778) );
  NANDN U12923 ( .A(n12616), .B(n12615), .Z(n12620) );
  NANDN U12924 ( .A(n12618), .B(n12617), .Z(n12619) );
  NAND U12925 ( .A(n12620), .B(n12619), .Z(n12779) );
  XNOR U12926 ( .A(n12778), .B(n12779), .Z(n12722) );
  XNOR U12927 ( .A(n12723), .B(n12722), .Z(n12725) );
  NANDN U12928 ( .A(n12622), .B(n12621), .Z(n12626) );
  NANDN U12929 ( .A(n12624), .B(n12623), .Z(n12625) );
  AND U12930 ( .A(n12626), .B(n12625), .Z(n12724) );
  XOR U12931 ( .A(n12725), .B(n12724), .Z(n12837) );
  NANDN U12932 ( .A(n12628), .B(n12627), .Z(n12632) );
  NANDN U12933 ( .A(n12630), .B(n12629), .Z(n12631) );
  AND U12934 ( .A(n12632), .B(n12631), .Z(n12834) );
  NANDN U12935 ( .A(n12634), .B(n12633), .Z(n12638) );
  NANDN U12936 ( .A(n12636), .B(n12635), .Z(n12637) );
  AND U12937 ( .A(n12638), .B(n12637), .Z(n12719) );
  NANDN U12938 ( .A(n12640), .B(n12639), .Z(n12644) );
  OR U12939 ( .A(n12642), .B(n12641), .Z(n12643) );
  AND U12940 ( .A(n12644), .B(n12643), .Z(n12717) );
  NANDN U12941 ( .A(n12646), .B(n12645), .Z(n12650) );
  NANDN U12942 ( .A(n12648), .B(n12647), .Z(n12649) );
  AND U12943 ( .A(n12650), .B(n12649), .Z(n12783) );
  NANDN U12944 ( .A(n12652), .B(n12651), .Z(n12656) );
  NANDN U12945 ( .A(n12654), .B(n12653), .Z(n12655) );
  NAND U12946 ( .A(n12656), .B(n12655), .Z(n12782) );
  XNOR U12947 ( .A(n12783), .B(n12782), .Z(n12785) );
  NAND U12948 ( .A(b[0]), .B(a[100]), .Z(n12657) );
  XNOR U12949 ( .A(b[1]), .B(n12657), .Z(n12659) );
  NANDN U12950 ( .A(b[0]), .B(a[99]), .Z(n12658) );
  NAND U12951 ( .A(n12659), .B(n12658), .Z(n12731) );
  NANDN U12952 ( .A(n19394), .B(n12660), .Z(n12662) );
  XOR U12953 ( .A(b[29]), .B(a[72]), .Z(n12807) );
  NANDN U12954 ( .A(n19395), .B(n12807), .Z(n12661) );
  AND U12955 ( .A(n12662), .B(n12661), .Z(n12729) );
  AND U12956 ( .A(b[31]), .B(a[68]), .Z(n12728) );
  XNOR U12957 ( .A(n12729), .B(n12728), .Z(n12730) );
  XNOR U12958 ( .A(n12731), .B(n12730), .Z(n12771) );
  NANDN U12959 ( .A(n19005), .B(n12663), .Z(n12665) );
  XOR U12960 ( .A(b[23]), .B(a[78]), .Z(n12810) );
  NANDN U12961 ( .A(n19055), .B(n12810), .Z(n12664) );
  AND U12962 ( .A(n12665), .B(n12664), .Z(n12800) );
  NANDN U12963 ( .A(n17362), .B(n12666), .Z(n12668) );
  XOR U12964 ( .A(b[7]), .B(a[94]), .Z(n12813) );
  NANDN U12965 ( .A(n17522), .B(n12813), .Z(n12667) );
  AND U12966 ( .A(n12668), .B(n12667), .Z(n12799) );
  NANDN U12967 ( .A(n19116), .B(n12669), .Z(n12671) );
  XOR U12968 ( .A(b[25]), .B(a[76]), .Z(n12816) );
  NANDN U12969 ( .A(n19179), .B(n12816), .Z(n12670) );
  NAND U12970 ( .A(n12671), .B(n12670), .Z(n12798) );
  XOR U12971 ( .A(n12799), .B(n12798), .Z(n12801) );
  XOR U12972 ( .A(n12800), .B(n12801), .Z(n12770) );
  XOR U12973 ( .A(n12771), .B(n12770), .Z(n12773) );
  NANDN U12974 ( .A(n18113), .B(n12672), .Z(n12674) );
  XOR U12975 ( .A(b[13]), .B(a[88]), .Z(n12819) );
  NANDN U12976 ( .A(n18229), .B(n12819), .Z(n12673) );
  AND U12977 ( .A(n12674), .B(n12673), .Z(n12765) );
  NANDN U12978 ( .A(n17888), .B(n12675), .Z(n12677) );
  XOR U12979 ( .A(b[11]), .B(a[90]), .Z(n12822) );
  NANDN U12980 ( .A(n18025), .B(n12822), .Z(n12676) );
  NAND U12981 ( .A(n12677), .B(n12676), .Z(n12764) );
  XNOR U12982 ( .A(n12765), .B(n12764), .Z(n12767) );
  NANDN U12983 ( .A(n18487), .B(n12678), .Z(n12680) );
  XOR U12984 ( .A(b[15]), .B(a[86]), .Z(n12825) );
  NANDN U12985 ( .A(n18311), .B(n12825), .Z(n12679) );
  AND U12986 ( .A(n12680), .B(n12679), .Z(n12761) );
  NANDN U12987 ( .A(n18853), .B(n12681), .Z(n12683) );
  XOR U12988 ( .A(b[21]), .B(a[80]), .Z(n12828) );
  NANDN U12989 ( .A(n18926), .B(n12828), .Z(n12682) );
  AND U12990 ( .A(n12683), .B(n12682), .Z(n12759) );
  NANDN U12991 ( .A(n17613), .B(n12684), .Z(n12686) );
  XOR U12992 ( .A(b[9]), .B(a[92]), .Z(n12831) );
  NANDN U12993 ( .A(n17739), .B(n12831), .Z(n12685) );
  NAND U12994 ( .A(n12686), .B(n12685), .Z(n12758) );
  XNOR U12995 ( .A(n12759), .B(n12758), .Z(n12760) );
  XNOR U12996 ( .A(n12761), .B(n12760), .Z(n12766) );
  XOR U12997 ( .A(n12767), .B(n12766), .Z(n12772) );
  XOR U12998 ( .A(n12773), .B(n12772), .Z(n12784) );
  XOR U12999 ( .A(n12785), .B(n12784), .Z(n12716) );
  XNOR U13000 ( .A(n12717), .B(n12716), .Z(n12718) );
  XOR U13001 ( .A(n12719), .B(n12718), .Z(n12835) );
  XNOR U13002 ( .A(n12834), .B(n12835), .Z(n12836) );
  XNOR U13003 ( .A(n12837), .B(n12836), .Z(n12712) );
  XOR U13004 ( .A(n12713), .B(n12712), .Z(n12705) );
  NANDN U13005 ( .A(n12688), .B(n12687), .Z(n12692) );
  OR U13006 ( .A(n12690), .B(n12689), .Z(n12691) );
  AND U13007 ( .A(n12692), .B(n12691), .Z(n12704) );
  XNOR U13008 ( .A(n12705), .B(n12704), .Z(n12706) );
  XNOR U13009 ( .A(n12707), .B(n12706), .Z(n12698) );
  XNOR U13010 ( .A(n12699), .B(n12698), .Z(n12700) );
  XNOR U13011 ( .A(n12701), .B(n12700), .Z(n12840) );
  XNOR U13012 ( .A(sreg[196]), .B(n12840), .Z(n12842) );
  NANDN U13013 ( .A(sreg[195]), .B(n12693), .Z(n12697) );
  NAND U13014 ( .A(n12695), .B(n12694), .Z(n12696) );
  NAND U13015 ( .A(n12697), .B(n12696), .Z(n12841) );
  XNOR U13016 ( .A(n12842), .B(n12841), .Z(c[196]) );
  NANDN U13017 ( .A(n12699), .B(n12698), .Z(n12703) );
  NANDN U13018 ( .A(n12701), .B(n12700), .Z(n12702) );
  AND U13019 ( .A(n12703), .B(n12702), .Z(n12848) );
  NANDN U13020 ( .A(n12705), .B(n12704), .Z(n12709) );
  NANDN U13021 ( .A(n12707), .B(n12706), .Z(n12708) );
  AND U13022 ( .A(n12709), .B(n12708), .Z(n12846) );
  NANDN U13023 ( .A(n12711), .B(n12710), .Z(n12715) );
  NAND U13024 ( .A(n12713), .B(n12712), .Z(n12714) );
  AND U13025 ( .A(n12715), .B(n12714), .Z(n12853) );
  NANDN U13026 ( .A(n12717), .B(n12716), .Z(n12721) );
  NANDN U13027 ( .A(n12719), .B(n12718), .Z(n12720) );
  AND U13028 ( .A(n12721), .B(n12720), .Z(n12984) );
  NANDN U13029 ( .A(n12723), .B(n12722), .Z(n12727) );
  NAND U13030 ( .A(n12725), .B(n12724), .Z(n12726) );
  AND U13031 ( .A(n12727), .B(n12726), .Z(n12983) );
  XNOR U13032 ( .A(n12984), .B(n12983), .Z(n12986) );
  NANDN U13033 ( .A(n12729), .B(n12728), .Z(n12733) );
  NANDN U13034 ( .A(n12731), .B(n12730), .Z(n12732) );
  AND U13035 ( .A(n12733), .B(n12732), .Z(n12919) );
  NANDN U13036 ( .A(n19237), .B(n12734), .Z(n12736) );
  XOR U13037 ( .A(b[27]), .B(a[75]), .Z(n12863) );
  NANDN U13038 ( .A(n19277), .B(n12863), .Z(n12735) );
  AND U13039 ( .A(n12736), .B(n12735), .Z(n12926) );
  NANDN U13040 ( .A(n17072), .B(n12737), .Z(n12739) );
  XOR U13041 ( .A(b[5]), .B(a[97]), .Z(n12866) );
  NANDN U13042 ( .A(n17223), .B(n12866), .Z(n12738) );
  AND U13043 ( .A(n12739), .B(n12738), .Z(n12924) );
  NANDN U13044 ( .A(n18673), .B(n12740), .Z(n12742) );
  XOR U13045 ( .A(b[19]), .B(a[83]), .Z(n12869) );
  NANDN U13046 ( .A(n18758), .B(n12869), .Z(n12741) );
  NAND U13047 ( .A(n12742), .B(n12741), .Z(n12923) );
  XNOR U13048 ( .A(n12924), .B(n12923), .Z(n12925) );
  XNOR U13049 ( .A(n12926), .B(n12925), .Z(n12917) );
  NANDN U13050 ( .A(n19425), .B(n12743), .Z(n12745) );
  XOR U13051 ( .A(b[31]), .B(a[71]), .Z(n12872) );
  NANDN U13052 ( .A(n19426), .B(n12872), .Z(n12744) );
  AND U13053 ( .A(n12745), .B(n12744), .Z(n12884) );
  NANDN U13054 ( .A(n17067), .B(n12746), .Z(n12748) );
  XOR U13055 ( .A(b[3]), .B(a[99]), .Z(n12875) );
  NANDN U13056 ( .A(n17068), .B(n12875), .Z(n12747) );
  AND U13057 ( .A(n12748), .B(n12747), .Z(n12882) );
  NANDN U13058 ( .A(n18514), .B(n12749), .Z(n12751) );
  XOR U13059 ( .A(b[17]), .B(a[85]), .Z(n12878) );
  NANDN U13060 ( .A(n18585), .B(n12878), .Z(n12750) );
  NAND U13061 ( .A(n12751), .B(n12750), .Z(n12881) );
  XNOR U13062 ( .A(n12882), .B(n12881), .Z(n12883) );
  XOR U13063 ( .A(n12884), .B(n12883), .Z(n12918) );
  XOR U13064 ( .A(n12917), .B(n12918), .Z(n12920) );
  XOR U13065 ( .A(n12919), .B(n12920), .Z(n12966) );
  NANDN U13066 ( .A(n12753), .B(n12752), .Z(n12757) );
  NANDN U13067 ( .A(n12755), .B(n12754), .Z(n12756) );
  AND U13068 ( .A(n12757), .B(n12756), .Z(n12905) );
  NANDN U13069 ( .A(n12759), .B(n12758), .Z(n12763) );
  NANDN U13070 ( .A(n12761), .B(n12760), .Z(n12762) );
  NAND U13071 ( .A(n12763), .B(n12762), .Z(n12906) );
  XNOR U13072 ( .A(n12905), .B(n12906), .Z(n12907) );
  NANDN U13073 ( .A(n12765), .B(n12764), .Z(n12769) );
  NAND U13074 ( .A(n12767), .B(n12766), .Z(n12768) );
  NAND U13075 ( .A(n12769), .B(n12768), .Z(n12908) );
  XNOR U13076 ( .A(n12907), .B(n12908), .Z(n12965) );
  XNOR U13077 ( .A(n12966), .B(n12965), .Z(n12968) );
  NAND U13078 ( .A(n12771), .B(n12770), .Z(n12775) );
  NAND U13079 ( .A(n12773), .B(n12772), .Z(n12774) );
  AND U13080 ( .A(n12775), .B(n12774), .Z(n12967) );
  XOR U13081 ( .A(n12968), .B(n12967), .Z(n12980) );
  NANDN U13082 ( .A(n12777), .B(n12776), .Z(n12781) );
  NANDN U13083 ( .A(n12779), .B(n12778), .Z(n12780) );
  AND U13084 ( .A(n12781), .B(n12780), .Z(n12977) );
  NANDN U13085 ( .A(n12787), .B(n12786), .Z(n12791) );
  OR U13086 ( .A(n12789), .B(n12788), .Z(n12790) );
  AND U13087 ( .A(n12791), .B(n12790), .Z(n12972) );
  NANDN U13088 ( .A(n12793), .B(n12792), .Z(n12797) );
  NANDN U13089 ( .A(n12795), .B(n12794), .Z(n12796) );
  AND U13090 ( .A(n12797), .B(n12796), .Z(n12912) );
  NANDN U13091 ( .A(n12799), .B(n12798), .Z(n12803) );
  OR U13092 ( .A(n12801), .B(n12800), .Z(n12802) );
  NAND U13093 ( .A(n12803), .B(n12802), .Z(n12911) );
  XNOR U13094 ( .A(n12912), .B(n12911), .Z(n12913) );
  NAND U13095 ( .A(b[0]), .B(a[101]), .Z(n12804) );
  XNOR U13096 ( .A(b[1]), .B(n12804), .Z(n12806) );
  NANDN U13097 ( .A(b[0]), .B(a[100]), .Z(n12805) );
  NAND U13098 ( .A(n12806), .B(n12805), .Z(n12860) );
  NANDN U13099 ( .A(n19394), .B(n12807), .Z(n12809) );
  XOR U13100 ( .A(b[29]), .B(a[73]), .Z(n12935) );
  NANDN U13101 ( .A(n19395), .B(n12935), .Z(n12808) );
  AND U13102 ( .A(n12809), .B(n12808), .Z(n12858) );
  AND U13103 ( .A(b[31]), .B(a[69]), .Z(n12857) );
  XNOR U13104 ( .A(n12858), .B(n12857), .Z(n12859) );
  XNOR U13105 ( .A(n12860), .B(n12859), .Z(n12899) );
  NANDN U13106 ( .A(n19005), .B(n12810), .Z(n12812) );
  XOR U13107 ( .A(b[23]), .B(a[79]), .Z(n12941) );
  NANDN U13108 ( .A(n19055), .B(n12941), .Z(n12811) );
  AND U13109 ( .A(n12812), .B(n12811), .Z(n12932) );
  NANDN U13110 ( .A(n17362), .B(n12813), .Z(n12815) );
  XOR U13111 ( .A(b[7]), .B(a[95]), .Z(n12944) );
  NANDN U13112 ( .A(n17522), .B(n12944), .Z(n12814) );
  AND U13113 ( .A(n12815), .B(n12814), .Z(n12930) );
  NANDN U13114 ( .A(n19116), .B(n12816), .Z(n12818) );
  XOR U13115 ( .A(b[25]), .B(a[77]), .Z(n12947) );
  NANDN U13116 ( .A(n19179), .B(n12947), .Z(n12817) );
  NAND U13117 ( .A(n12818), .B(n12817), .Z(n12929) );
  XNOR U13118 ( .A(n12930), .B(n12929), .Z(n12931) );
  XOR U13119 ( .A(n12932), .B(n12931), .Z(n12900) );
  XNOR U13120 ( .A(n12899), .B(n12900), .Z(n12901) );
  NANDN U13121 ( .A(n18113), .B(n12819), .Z(n12821) );
  XOR U13122 ( .A(b[13]), .B(a[89]), .Z(n12950) );
  NANDN U13123 ( .A(n18229), .B(n12950), .Z(n12820) );
  AND U13124 ( .A(n12821), .B(n12820), .Z(n12894) );
  NANDN U13125 ( .A(n17888), .B(n12822), .Z(n12824) );
  XOR U13126 ( .A(b[11]), .B(a[91]), .Z(n12953) );
  NANDN U13127 ( .A(n18025), .B(n12953), .Z(n12823) );
  NAND U13128 ( .A(n12824), .B(n12823), .Z(n12893) );
  XNOR U13129 ( .A(n12894), .B(n12893), .Z(n12895) );
  NANDN U13130 ( .A(n18487), .B(n12825), .Z(n12827) );
  XOR U13131 ( .A(b[15]), .B(a[87]), .Z(n12956) );
  NANDN U13132 ( .A(n18311), .B(n12956), .Z(n12826) );
  AND U13133 ( .A(n12827), .B(n12826), .Z(n12890) );
  NANDN U13134 ( .A(n18853), .B(n12828), .Z(n12830) );
  XOR U13135 ( .A(b[21]), .B(a[81]), .Z(n12959) );
  NANDN U13136 ( .A(n18926), .B(n12959), .Z(n12829) );
  AND U13137 ( .A(n12830), .B(n12829), .Z(n12888) );
  NANDN U13138 ( .A(n17613), .B(n12831), .Z(n12833) );
  XOR U13139 ( .A(b[9]), .B(a[93]), .Z(n12962) );
  NANDN U13140 ( .A(n17739), .B(n12962), .Z(n12832) );
  NAND U13141 ( .A(n12833), .B(n12832), .Z(n12887) );
  XNOR U13142 ( .A(n12888), .B(n12887), .Z(n12889) );
  XOR U13143 ( .A(n12890), .B(n12889), .Z(n12896) );
  XOR U13144 ( .A(n12895), .B(n12896), .Z(n12902) );
  XOR U13145 ( .A(n12901), .B(n12902), .Z(n12914) );
  XNOR U13146 ( .A(n12913), .B(n12914), .Z(n12971) );
  XNOR U13147 ( .A(n12972), .B(n12971), .Z(n12973) );
  XOR U13148 ( .A(n12974), .B(n12973), .Z(n12978) );
  XNOR U13149 ( .A(n12977), .B(n12978), .Z(n12979) );
  XNOR U13150 ( .A(n12980), .B(n12979), .Z(n12985) );
  XOR U13151 ( .A(n12986), .B(n12985), .Z(n12852) );
  NANDN U13152 ( .A(n12835), .B(n12834), .Z(n12839) );
  NANDN U13153 ( .A(n12837), .B(n12836), .Z(n12838) );
  AND U13154 ( .A(n12839), .B(n12838), .Z(n12851) );
  XOR U13155 ( .A(n12852), .B(n12851), .Z(n12854) );
  XNOR U13156 ( .A(n12853), .B(n12854), .Z(n12845) );
  XNOR U13157 ( .A(n12846), .B(n12845), .Z(n12847) );
  XNOR U13158 ( .A(n12848), .B(n12847), .Z(n12989) );
  XNOR U13159 ( .A(sreg[197]), .B(n12989), .Z(n12991) );
  NANDN U13160 ( .A(sreg[196]), .B(n12840), .Z(n12844) );
  NAND U13161 ( .A(n12842), .B(n12841), .Z(n12843) );
  NAND U13162 ( .A(n12844), .B(n12843), .Z(n12990) );
  XNOR U13163 ( .A(n12991), .B(n12990), .Z(c[197]) );
  NANDN U13164 ( .A(n12846), .B(n12845), .Z(n12850) );
  NANDN U13165 ( .A(n12848), .B(n12847), .Z(n12849) );
  AND U13166 ( .A(n12850), .B(n12849), .Z(n12997) );
  NANDN U13167 ( .A(n12852), .B(n12851), .Z(n12856) );
  NANDN U13168 ( .A(n12854), .B(n12853), .Z(n12855) );
  AND U13169 ( .A(n12856), .B(n12855), .Z(n12995) );
  NANDN U13170 ( .A(n12858), .B(n12857), .Z(n12862) );
  NANDN U13171 ( .A(n12860), .B(n12859), .Z(n12861) );
  AND U13172 ( .A(n12862), .B(n12861), .Z(n13086) );
  NANDN U13173 ( .A(n19237), .B(n12863), .Z(n12865) );
  XOR U13174 ( .A(b[27]), .B(a[76]), .Z(n13030) );
  NANDN U13175 ( .A(n19277), .B(n13030), .Z(n12864) );
  AND U13176 ( .A(n12865), .B(n12864), .Z(n13093) );
  NANDN U13177 ( .A(n17072), .B(n12866), .Z(n12868) );
  XOR U13178 ( .A(b[5]), .B(a[98]), .Z(n13033) );
  NANDN U13179 ( .A(n17223), .B(n13033), .Z(n12867) );
  AND U13180 ( .A(n12868), .B(n12867), .Z(n13091) );
  NANDN U13181 ( .A(n18673), .B(n12869), .Z(n12871) );
  XOR U13182 ( .A(b[19]), .B(a[84]), .Z(n13036) );
  NANDN U13183 ( .A(n18758), .B(n13036), .Z(n12870) );
  NAND U13184 ( .A(n12871), .B(n12870), .Z(n13090) );
  XNOR U13185 ( .A(n13091), .B(n13090), .Z(n13092) );
  XNOR U13186 ( .A(n13093), .B(n13092), .Z(n13084) );
  NANDN U13187 ( .A(n19425), .B(n12872), .Z(n12874) );
  XOR U13188 ( .A(b[31]), .B(a[72]), .Z(n13039) );
  NANDN U13189 ( .A(n19426), .B(n13039), .Z(n12873) );
  AND U13190 ( .A(n12874), .B(n12873), .Z(n13051) );
  NANDN U13191 ( .A(n17067), .B(n12875), .Z(n12877) );
  XOR U13192 ( .A(b[3]), .B(a[100]), .Z(n13042) );
  NANDN U13193 ( .A(n17068), .B(n13042), .Z(n12876) );
  AND U13194 ( .A(n12877), .B(n12876), .Z(n13049) );
  NANDN U13195 ( .A(n18514), .B(n12878), .Z(n12880) );
  XOR U13196 ( .A(b[17]), .B(a[86]), .Z(n13045) );
  NANDN U13197 ( .A(n18585), .B(n13045), .Z(n12879) );
  NAND U13198 ( .A(n12880), .B(n12879), .Z(n13048) );
  XNOR U13199 ( .A(n13049), .B(n13048), .Z(n13050) );
  XOR U13200 ( .A(n13051), .B(n13050), .Z(n13085) );
  XOR U13201 ( .A(n13084), .B(n13085), .Z(n13087) );
  XOR U13202 ( .A(n13086), .B(n13087), .Z(n13019) );
  NANDN U13203 ( .A(n12882), .B(n12881), .Z(n12886) );
  NANDN U13204 ( .A(n12884), .B(n12883), .Z(n12885) );
  AND U13205 ( .A(n12886), .B(n12885), .Z(n13072) );
  NANDN U13206 ( .A(n12888), .B(n12887), .Z(n12892) );
  NANDN U13207 ( .A(n12890), .B(n12889), .Z(n12891) );
  NAND U13208 ( .A(n12892), .B(n12891), .Z(n13073) );
  XNOR U13209 ( .A(n13072), .B(n13073), .Z(n13074) );
  NANDN U13210 ( .A(n12894), .B(n12893), .Z(n12898) );
  NANDN U13211 ( .A(n12896), .B(n12895), .Z(n12897) );
  NAND U13212 ( .A(n12898), .B(n12897), .Z(n13075) );
  XNOR U13213 ( .A(n13074), .B(n13075), .Z(n13018) );
  XNOR U13214 ( .A(n13019), .B(n13018), .Z(n13021) );
  NANDN U13215 ( .A(n12900), .B(n12899), .Z(n12904) );
  NANDN U13216 ( .A(n12902), .B(n12901), .Z(n12903) );
  AND U13217 ( .A(n12904), .B(n12903), .Z(n13020) );
  XOR U13218 ( .A(n13021), .B(n13020), .Z(n13134) );
  NANDN U13219 ( .A(n12906), .B(n12905), .Z(n12910) );
  NANDN U13220 ( .A(n12908), .B(n12907), .Z(n12909) );
  AND U13221 ( .A(n12910), .B(n12909), .Z(n13132) );
  NANDN U13222 ( .A(n12912), .B(n12911), .Z(n12916) );
  NANDN U13223 ( .A(n12914), .B(n12913), .Z(n12915) );
  AND U13224 ( .A(n12916), .B(n12915), .Z(n13015) );
  NANDN U13225 ( .A(n12918), .B(n12917), .Z(n12922) );
  OR U13226 ( .A(n12920), .B(n12919), .Z(n12921) );
  AND U13227 ( .A(n12922), .B(n12921), .Z(n13013) );
  NANDN U13228 ( .A(n12924), .B(n12923), .Z(n12928) );
  NANDN U13229 ( .A(n12926), .B(n12925), .Z(n12927) );
  AND U13230 ( .A(n12928), .B(n12927), .Z(n13079) );
  NANDN U13231 ( .A(n12930), .B(n12929), .Z(n12934) );
  NANDN U13232 ( .A(n12932), .B(n12931), .Z(n12933) );
  NAND U13233 ( .A(n12934), .B(n12933), .Z(n13078) );
  XNOR U13234 ( .A(n13079), .B(n13078), .Z(n13080) );
  NANDN U13235 ( .A(n19394), .B(n12935), .Z(n12937) );
  XOR U13236 ( .A(b[29]), .B(a[74]), .Z(n13105) );
  NANDN U13237 ( .A(n19395), .B(n13105), .Z(n12936) );
  AND U13238 ( .A(n12937), .B(n12936), .Z(n13025) );
  AND U13239 ( .A(b[31]), .B(a[70]), .Z(n13024) );
  XNOR U13240 ( .A(n13025), .B(n13024), .Z(n13026) );
  NAND U13241 ( .A(b[0]), .B(a[102]), .Z(n12938) );
  XNOR U13242 ( .A(b[1]), .B(n12938), .Z(n12940) );
  NANDN U13243 ( .A(b[0]), .B(a[101]), .Z(n12939) );
  NAND U13244 ( .A(n12940), .B(n12939), .Z(n13027) );
  XNOR U13245 ( .A(n13026), .B(n13027), .Z(n13066) );
  NANDN U13246 ( .A(n19005), .B(n12941), .Z(n12943) );
  XOR U13247 ( .A(b[23]), .B(a[80]), .Z(n13108) );
  NANDN U13248 ( .A(n19055), .B(n13108), .Z(n12942) );
  AND U13249 ( .A(n12943), .B(n12942), .Z(n13099) );
  NANDN U13250 ( .A(n17362), .B(n12944), .Z(n12946) );
  XOR U13251 ( .A(b[7]), .B(a[96]), .Z(n13111) );
  NANDN U13252 ( .A(n17522), .B(n13111), .Z(n12945) );
  AND U13253 ( .A(n12946), .B(n12945), .Z(n13097) );
  NANDN U13254 ( .A(n19116), .B(n12947), .Z(n12949) );
  XOR U13255 ( .A(b[25]), .B(a[78]), .Z(n13114) );
  NANDN U13256 ( .A(n19179), .B(n13114), .Z(n12948) );
  NAND U13257 ( .A(n12949), .B(n12948), .Z(n13096) );
  XNOR U13258 ( .A(n13097), .B(n13096), .Z(n13098) );
  XOR U13259 ( .A(n13099), .B(n13098), .Z(n13067) );
  XNOR U13260 ( .A(n13066), .B(n13067), .Z(n13068) );
  NANDN U13261 ( .A(n18113), .B(n12950), .Z(n12952) );
  XOR U13262 ( .A(b[13]), .B(a[90]), .Z(n13117) );
  NANDN U13263 ( .A(n18229), .B(n13117), .Z(n12951) );
  AND U13264 ( .A(n12952), .B(n12951), .Z(n13061) );
  NANDN U13265 ( .A(n17888), .B(n12953), .Z(n12955) );
  XOR U13266 ( .A(b[11]), .B(a[92]), .Z(n13120) );
  NANDN U13267 ( .A(n18025), .B(n13120), .Z(n12954) );
  NAND U13268 ( .A(n12955), .B(n12954), .Z(n13060) );
  XNOR U13269 ( .A(n13061), .B(n13060), .Z(n13062) );
  NANDN U13270 ( .A(n18487), .B(n12956), .Z(n12958) );
  XOR U13271 ( .A(b[15]), .B(a[88]), .Z(n13123) );
  NANDN U13272 ( .A(n18311), .B(n13123), .Z(n12957) );
  AND U13273 ( .A(n12958), .B(n12957), .Z(n13057) );
  NANDN U13274 ( .A(n18853), .B(n12959), .Z(n12961) );
  XOR U13275 ( .A(b[21]), .B(a[82]), .Z(n13126) );
  NANDN U13276 ( .A(n18926), .B(n13126), .Z(n12960) );
  AND U13277 ( .A(n12961), .B(n12960), .Z(n13055) );
  NANDN U13278 ( .A(n17613), .B(n12962), .Z(n12964) );
  XOR U13279 ( .A(b[9]), .B(a[94]), .Z(n13129) );
  NANDN U13280 ( .A(n17739), .B(n13129), .Z(n12963) );
  NAND U13281 ( .A(n12964), .B(n12963), .Z(n13054) );
  XNOR U13282 ( .A(n13055), .B(n13054), .Z(n13056) );
  XOR U13283 ( .A(n13057), .B(n13056), .Z(n13063) );
  XOR U13284 ( .A(n13062), .B(n13063), .Z(n13069) );
  XOR U13285 ( .A(n13068), .B(n13069), .Z(n13081) );
  XNOR U13286 ( .A(n13080), .B(n13081), .Z(n13012) );
  XNOR U13287 ( .A(n13013), .B(n13012), .Z(n13014) );
  XOR U13288 ( .A(n13015), .B(n13014), .Z(n13133) );
  XOR U13289 ( .A(n13132), .B(n13133), .Z(n13135) );
  XOR U13290 ( .A(n13134), .B(n13135), .Z(n13009) );
  NANDN U13291 ( .A(n12966), .B(n12965), .Z(n12970) );
  NAND U13292 ( .A(n12968), .B(n12967), .Z(n12969) );
  AND U13293 ( .A(n12970), .B(n12969), .Z(n13007) );
  NANDN U13294 ( .A(n12972), .B(n12971), .Z(n12976) );
  NANDN U13295 ( .A(n12974), .B(n12973), .Z(n12975) );
  AND U13296 ( .A(n12976), .B(n12975), .Z(n13006) );
  XNOR U13297 ( .A(n13007), .B(n13006), .Z(n13008) );
  XNOR U13298 ( .A(n13009), .B(n13008), .Z(n13000) );
  NANDN U13299 ( .A(n12978), .B(n12977), .Z(n12982) );
  NANDN U13300 ( .A(n12980), .B(n12979), .Z(n12981) );
  NAND U13301 ( .A(n12982), .B(n12981), .Z(n13001) );
  XNOR U13302 ( .A(n13000), .B(n13001), .Z(n13002) );
  NANDN U13303 ( .A(n12984), .B(n12983), .Z(n12988) );
  NAND U13304 ( .A(n12986), .B(n12985), .Z(n12987) );
  NAND U13305 ( .A(n12988), .B(n12987), .Z(n13003) );
  XNOR U13306 ( .A(n13002), .B(n13003), .Z(n12994) );
  XNOR U13307 ( .A(n12995), .B(n12994), .Z(n12996) );
  XNOR U13308 ( .A(n12997), .B(n12996), .Z(n13138) );
  XNOR U13309 ( .A(sreg[198]), .B(n13138), .Z(n13140) );
  NANDN U13310 ( .A(sreg[197]), .B(n12989), .Z(n12993) );
  NAND U13311 ( .A(n12991), .B(n12990), .Z(n12992) );
  NAND U13312 ( .A(n12993), .B(n12992), .Z(n13139) );
  XNOR U13313 ( .A(n13140), .B(n13139), .Z(c[198]) );
  NANDN U13314 ( .A(n12995), .B(n12994), .Z(n12999) );
  NANDN U13315 ( .A(n12997), .B(n12996), .Z(n12998) );
  AND U13316 ( .A(n12999), .B(n12998), .Z(n13146) );
  NANDN U13317 ( .A(n13001), .B(n13000), .Z(n13005) );
  NANDN U13318 ( .A(n13003), .B(n13002), .Z(n13004) );
  AND U13319 ( .A(n13005), .B(n13004), .Z(n13144) );
  NANDN U13320 ( .A(n13007), .B(n13006), .Z(n13011) );
  NANDN U13321 ( .A(n13009), .B(n13008), .Z(n13010) );
  AND U13322 ( .A(n13011), .B(n13010), .Z(n13152) );
  NANDN U13323 ( .A(n13013), .B(n13012), .Z(n13017) );
  NANDN U13324 ( .A(n13015), .B(n13014), .Z(n13016) );
  AND U13325 ( .A(n13017), .B(n13016), .Z(n13156) );
  NANDN U13326 ( .A(n13019), .B(n13018), .Z(n13023) );
  NAND U13327 ( .A(n13021), .B(n13020), .Z(n13022) );
  AND U13328 ( .A(n13023), .B(n13022), .Z(n13155) );
  XNOR U13329 ( .A(n13156), .B(n13155), .Z(n13158) );
  NANDN U13330 ( .A(n13025), .B(n13024), .Z(n13029) );
  NANDN U13331 ( .A(n13027), .B(n13026), .Z(n13028) );
  AND U13332 ( .A(n13029), .B(n13028), .Z(n13235) );
  NANDN U13333 ( .A(n19237), .B(n13030), .Z(n13032) );
  XOR U13334 ( .A(b[27]), .B(a[77]), .Z(n13179) );
  NANDN U13335 ( .A(n19277), .B(n13179), .Z(n13031) );
  AND U13336 ( .A(n13032), .B(n13031), .Z(n13242) );
  NANDN U13337 ( .A(n17072), .B(n13033), .Z(n13035) );
  XOR U13338 ( .A(b[5]), .B(a[99]), .Z(n13182) );
  NANDN U13339 ( .A(n17223), .B(n13182), .Z(n13034) );
  AND U13340 ( .A(n13035), .B(n13034), .Z(n13240) );
  NANDN U13341 ( .A(n18673), .B(n13036), .Z(n13038) );
  XOR U13342 ( .A(b[19]), .B(a[85]), .Z(n13185) );
  NANDN U13343 ( .A(n18758), .B(n13185), .Z(n13037) );
  NAND U13344 ( .A(n13038), .B(n13037), .Z(n13239) );
  XNOR U13345 ( .A(n13240), .B(n13239), .Z(n13241) );
  XNOR U13346 ( .A(n13242), .B(n13241), .Z(n13233) );
  NANDN U13347 ( .A(n19425), .B(n13039), .Z(n13041) );
  XOR U13348 ( .A(b[31]), .B(a[73]), .Z(n13188) );
  NANDN U13349 ( .A(n19426), .B(n13188), .Z(n13040) );
  AND U13350 ( .A(n13041), .B(n13040), .Z(n13200) );
  NANDN U13351 ( .A(n17067), .B(n13042), .Z(n13044) );
  XOR U13352 ( .A(b[3]), .B(a[101]), .Z(n13191) );
  NANDN U13353 ( .A(n17068), .B(n13191), .Z(n13043) );
  AND U13354 ( .A(n13044), .B(n13043), .Z(n13198) );
  NANDN U13355 ( .A(n18514), .B(n13045), .Z(n13047) );
  XOR U13356 ( .A(b[17]), .B(a[87]), .Z(n13194) );
  NANDN U13357 ( .A(n18585), .B(n13194), .Z(n13046) );
  NAND U13358 ( .A(n13047), .B(n13046), .Z(n13197) );
  XNOR U13359 ( .A(n13198), .B(n13197), .Z(n13199) );
  XOR U13360 ( .A(n13200), .B(n13199), .Z(n13234) );
  XOR U13361 ( .A(n13233), .B(n13234), .Z(n13236) );
  XOR U13362 ( .A(n13235), .B(n13236), .Z(n13168) );
  NANDN U13363 ( .A(n13049), .B(n13048), .Z(n13053) );
  NANDN U13364 ( .A(n13051), .B(n13050), .Z(n13052) );
  AND U13365 ( .A(n13053), .B(n13052), .Z(n13221) );
  NANDN U13366 ( .A(n13055), .B(n13054), .Z(n13059) );
  NANDN U13367 ( .A(n13057), .B(n13056), .Z(n13058) );
  NAND U13368 ( .A(n13059), .B(n13058), .Z(n13222) );
  XNOR U13369 ( .A(n13221), .B(n13222), .Z(n13223) );
  NANDN U13370 ( .A(n13061), .B(n13060), .Z(n13065) );
  NANDN U13371 ( .A(n13063), .B(n13062), .Z(n13064) );
  NAND U13372 ( .A(n13065), .B(n13064), .Z(n13224) );
  XNOR U13373 ( .A(n13223), .B(n13224), .Z(n13167) );
  XNOR U13374 ( .A(n13168), .B(n13167), .Z(n13170) );
  NANDN U13375 ( .A(n13067), .B(n13066), .Z(n13071) );
  NANDN U13376 ( .A(n13069), .B(n13068), .Z(n13070) );
  AND U13377 ( .A(n13071), .B(n13070), .Z(n13169) );
  XOR U13378 ( .A(n13170), .B(n13169), .Z(n13284) );
  NANDN U13379 ( .A(n13073), .B(n13072), .Z(n13077) );
  NANDN U13380 ( .A(n13075), .B(n13074), .Z(n13076) );
  AND U13381 ( .A(n13077), .B(n13076), .Z(n13281) );
  NANDN U13382 ( .A(n13079), .B(n13078), .Z(n13083) );
  NANDN U13383 ( .A(n13081), .B(n13080), .Z(n13082) );
  AND U13384 ( .A(n13083), .B(n13082), .Z(n13164) );
  NANDN U13385 ( .A(n13085), .B(n13084), .Z(n13089) );
  OR U13386 ( .A(n13087), .B(n13086), .Z(n13088) );
  AND U13387 ( .A(n13089), .B(n13088), .Z(n13162) );
  NANDN U13388 ( .A(n13091), .B(n13090), .Z(n13095) );
  NANDN U13389 ( .A(n13093), .B(n13092), .Z(n13094) );
  AND U13390 ( .A(n13095), .B(n13094), .Z(n13228) );
  NANDN U13391 ( .A(n13097), .B(n13096), .Z(n13101) );
  NANDN U13392 ( .A(n13099), .B(n13098), .Z(n13100) );
  NAND U13393 ( .A(n13101), .B(n13100), .Z(n13227) );
  XNOR U13394 ( .A(n13228), .B(n13227), .Z(n13229) );
  NAND U13395 ( .A(b[0]), .B(a[103]), .Z(n13102) );
  XNOR U13396 ( .A(b[1]), .B(n13102), .Z(n13104) );
  NANDN U13397 ( .A(b[0]), .B(a[102]), .Z(n13103) );
  NAND U13398 ( .A(n13104), .B(n13103), .Z(n13176) );
  NANDN U13399 ( .A(n19394), .B(n13105), .Z(n13107) );
  XOR U13400 ( .A(b[29]), .B(a[75]), .Z(n13251) );
  NANDN U13401 ( .A(n19395), .B(n13251), .Z(n13106) );
  AND U13402 ( .A(n13107), .B(n13106), .Z(n13174) );
  AND U13403 ( .A(b[31]), .B(a[71]), .Z(n13173) );
  XNOR U13404 ( .A(n13174), .B(n13173), .Z(n13175) );
  XNOR U13405 ( .A(n13176), .B(n13175), .Z(n13215) );
  NANDN U13406 ( .A(n19005), .B(n13108), .Z(n13110) );
  XOR U13407 ( .A(b[23]), .B(a[81]), .Z(n13257) );
  NANDN U13408 ( .A(n19055), .B(n13257), .Z(n13109) );
  AND U13409 ( .A(n13110), .B(n13109), .Z(n13248) );
  NANDN U13410 ( .A(n17362), .B(n13111), .Z(n13113) );
  XOR U13411 ( .A(b[7]), .B(a[97]), .Z(n13260) );
  NANDN U13412 ( .A(n17522), .B(n13260), .Z(n13112) );
  AND U13413 ( .A(n13113), .B(n13112), .Z(n13246) );
  NANDN U13414 ( .A(n19116), .B(n13114), .Z(n13116) );
  XOR U13415 ( .A(b[25]), .B(a[79]), .Z(n13263) );
  NANDN U13416 ( .A(n19179), .B(n13263), .Z(n13115) );
  NAND U13417 ( .A(n13116), .B(n13115), .Z(n13245) );
  XNOR U13418 ( .A(n13246), .B(n13245), .Z(n13247) );
  XOR U13419 ( .A(n13248), .B(n13247), .Z(n13216) );
  XNOR U13420 ( .A(n13215), .B(n13216), .Z(n13217) );
  NANDN U13421 ( .A(n18113), .B(n13117), .Z(n13119) );
  XOR U13422 ( .A(b[13]), .B(a[91]), .Z(n13266) );
  NANDN U13423 ( .A(n18229), .B(n13266), .Z(n13118) );
  AND U13424 ( .A(n13119), .B(n13118), .Z(n13210) );
  NANDN U13425 ( .A(n17888), .B(n13120), .Z(n13122) );
  XOR U13426 ( .A(b[11]), .B(a[93]), .Z(n13269) );
  NANDN U13427 ( .A(n18025), .B(n13269), .Z(n13121) );
  NAND U13428 ( .A(n13122), .B(n13121), .Z(n13209) );
  XNOR U13429 ( .A(n13210), .B(n13209), .Z(n13211) );
  NANDN U13430 ( .A(n18487), .B(n13123), .Z(n13125) );
  XOR U13431 ( .A(b[15]), .B(a[89]), .Z(n13272) );
  NANDN U13432 ( .A(n18311), .B(n13272), .Z(n13124) );
  AND U13433 ( .A(n13125), .B(n13124), .Z(n13206) );
  NANDN U13434 ( .A(n18853), .B(n13126), .Z(n13128) );
  XOR U13435 ( .A(b[21]), .B(a[83]), .Z(n13275) );
  NANDN U13436 ( .A(n18926), .B(n13275), .Z(n13127) );
  AND U13437 ( .A(n13128), .B(n13127), .Z(n13204) );
  NANDN U13438 ( .A(n17613), .B(n13129), .Z(n13131) );
  XOR U13439 ( .A(b[9]), .B(a[95]), .Z(n13278) );
  NANDN U13440 ( .A(n17739), .B(n13278), .Z(n13130) );
  NAND U13441 ( .A(n13131), .B(n13130), .Z(n13203) );
  XNOR U13442 ( .A(n13204), .B(n13203), .Z(n13205) );
  XOR U13443 ( .A(n13206), .B(n13205), .Z(n13212) );
  XOR U13444 ( .A(n13211), .B(n13212), .Z(n13218) );
  XOR U13445 ( .A(n13217), .B(n13218), .Z(n13230) );
  XNOR U13446 ( .A(n13229), .B(n13230), .Z(n13161) );
  XNOR U13447 ( .A(n13162), .B(n13161), .Z(n13163) );
  XOR U13448 ( .A(n13164), .B(n13163), .Z(n13282) );
  XNOR U13449 ( .A(n13281), .B(n13282), .Z(n13283) );
  XNOR U13450 ( .A(n13284), .B(n13283), .Z(n13157) );
  XOR U13451 ( .A(n13158), .B(n13157), .Z(n13150) );
  NANDN U13452 ( .A(n13133), .B(n13132), .Z(n13137) );
  OR U13453 ( .A(n13135), .B(n13134), .Z(n13136) );
  AND U13454 ( .A(n13137), .B(n13136), .Z(n13149) );
  XNOR U13455 ( .A(n13150), .B(n13149), .Z(n13151) );
  XNOR U13456 ( .A(n13152), .B(n13151), .Z(n13143) );
  XNOR U13457 ( .A(n13144), .B(n13143), .Z(n13145) );
  XNOR U13458 ( .A(n13146), .B(n13145), .Z(n13287) );
  XNOR U13459 ( .A(sreg[199]), .B(n13287), .Z(n13289) );
  NANDN U13460 ( .A(sreg[198]), .B(n13138), .Z(n13142) );
  NAND U13461 ( .A(n13140), .B(n13139), .Z(n13141) );
  NAND U13462 ( .A(n13142), .B(n13141), .Z(n13288) );
  XNOR U13463 ( .A(n13289), .B(n13288), .Z(c[199]) );
  NANDN U13464 ( .A(n13144), .B(n13143), .Z(n13148) );
  NANDN U13465 ( .A(n13146), .B(n13145), .Z(n13147) );
  AND U13466 ( .A(n13148), .B(n13147), .Z(n13295) );
  NANDN U13467 ( .A(n13150), .B(n13149), .Z(n13154) );
  NANDN U13468 ( .A(n13152), .B(n13151), .Z(n13153) );
  AND U13469 ( .A(n13154), .B(n13153), .Z(n13293) );
  NANDN U13470 ( .A(n13156), .B(n13155), .Z(n13160) );
  NAND U13471 ( .A(n13158), .B(n13157), .Z(n13159) );
  AND U13472 ( .A(n13160), .B(n13159), .Z(n13300) );
  NANDN U13473 ( .A(n13162), .B(n13161), .Z(n13166) );
  NANDN U13474 ( .A(n13164), .B(n13163), .Z(n13165) );
  AND U13475 ( .A(n13166), .B(n13165), .Z(n13305) );
  NANDN U13476 ( .A(n13168), .B(n13167), .Z(n13172) );
  NAND U13477 ( .A(n13170), .B(n13169), .Z(n13171) );
  AND U13478 ( .A(n13172), .B(n13171), .Z(n13304) );
  XNOR U13479 ( .A(n13305), .B(n13304), .Z(n13307) );
  NANDN U13480 ( .A(n13174), .B(n13173), .Z(n13178) );
  NANDN U13481 ( .A(n13176), .B(n13175), .Z(n13177) );
  AND U13482 ( .A(n13178), .B(n13177), .Z(n13384) );
  NANDN U13483 ( .A(n19237), .B(n13179), .Z(n13181) );
  XOR U13484 ( .A(b[27]), .B(a[78]), .Z(n13328) );
  NANDN U13485 ( .A(n19277), .B(n13328), .Z(n13180) );
  AND U13486 ( .A(n13181), .B(n13180), .Z(n13391) );
  NANDN U13487 ( .A(n17072), .B(n13182), .Z(n13184) );
  XOR U13488 ( .A(b[5]), .B(a[100]), .Z(n13331) );
  NANDN U13489 ( .A(n17223), .B(n13331), .Z(n13183) );
  AND U13490 ( .A(n13184), .B(n13183), .Z(n13389) );
  NANDN U13491 ( .A(n18673), .B(n13185), .Z(n13187) );
  XOR U13492 ( .A(b[19]), .B(a[86]), .Z(n13334) );
  NANDN U13493 ( .A(n18758), .B(n13334), .Z(n13186) );
  NAND U13494 ( .A(n13187), .B(n13186), .Z(n13388) );
  XNOR U13495 ( .A(n13389), .B(n13388), .Z(n13390) );
  XNOR U13496 ( .A(n13391), .B(n13390), .Z(n13382) );
  NANDN U13497 ( .A(n19425), .B(n13188), .Z(n13190) );
  XOR U13498 ( .A(b[31]), .B(a[74]), .Z(n13337) );
  NANDN U13499 ( .A(n19426), .B(n13337), .Z(n13189) );
  AND U13500 ( .A(n13190), .B(n13189), .Z(n13349) );
  NANDN U13501 ( .A(n17067), .B(n13191), .Z(n13193) );
  XOR U13502 ( .A(a[102]), .B(b[3]), .Z(n13340) );
  NANDN U13503 ( .A(n17068), .B(n13340), .Z(n13192) );
  AND U13504 ( .A(n13193), .B(n13192), .Z(n13347) );
  NANDN U13505 ( .A(n18514), .B(n13194), .Z(n13196) );
  XOR U13506 ( .A(b[17]), .B(a[88]), .Z(n13343) );
  NANDN U13507 ( .A(n18585), .B(n13343), .Z(n13195) );
  NAND U13508 ( .A(n13196), .B(n13195), .Z(n13346) );
  XNOR U13509 ( .A(n13347), .B(n13346), .Z(n13348) );
  XOR U13510 ( .A(n13349), .B(n13348), .Z(n13383) );
  XOR U13511 ( .A(n13382), .B(n13383), .Z(n13385) );
  XOR U13512 ( .A(n13384), .B(n13385), .Z(n13317) );
  NANDN U13513 ( .A(n13198), .B(n13197), .Z(n13202) );
  NANDN U13514 ( .A(n13200), .B(n13199), .Z(n13201) );
  AND U13515 ( .A(n13202), .B(n13201), .Z(n13370) );
  NANDN U13516 ( .A(n13204), .B(n13203), .Z(n13208) );
  NANDN U13517 ( .A(n13206), .B(n13205), .Z(n13207) );
  NAND U13518 ( .A(n13208), .B(n13207), .Z(n13371) );
  XNOR U13519 ( .A(n13370), .B(n13371), .Z(n13372) );
  NANDN U13520 ( .A(n13210), .B(n13209), .Z(n13214) );
  NANDN U13521 ( .A(n13212), .B(n13211), .Z(n13213) );
  NAND U13522 ( .A(n13214), .B(n13213), .Z(n13373) );
  XNOR U13523 ( .A(n13372), .B(n13373), .Z(n13316) );
  XNOR U13524 ( .A(n13317), .B(n13316), .Z(n13319) );
  NANDN U13525 ( .A(n13216), .B(n13215), .Z(n13220) );
  NANDN U13526 ( .A(n13218), .B(n13217), .Z(n13219) );
  AND U13527 ( .A(n13220), .B(n13219), .Z(n13318) );
  XOR U13528 ( .A(n13319), .B(n13318), .Z(n13433) );
  NANDN U13529 ( .A(n13222), .B(n13221), .Z(n13226) );
  NANDN U13530 ( .A(n13224), .B(n13223), .Z(n13225) );
  AND U13531 ( .A(n13226), .B(n13225), .Z(n13430) );
  NANDN U13532 ( .A(n13228), .B(n13227), .Z(n13232) );
  NANDN U13533 ( .A(n13230), .B(n13229), .Z(n13231) );
  AND U13534 ( .A(n13232), .B(n13231), .Z(n13313) );
  NANDN U13535 ( .A(n13234), .B(n13233), .Z(n13238) );
  OR U13536 ( .A(n13236), .B(n13235), .Z(n13237) );
  AND U13537 ( .A(n13238), .B(n13237), .Z(n13311) );
  NANDN U13538 ( .A(n13240), .B(n13239), .Z(n13244) );
  NANDN U13539 ( .A(n13242), .B(n13241), .Z(n13243) );
  AND U13540 ( .A(n13244), .B(n13243), .Z(n13377) );
  NANDN U13541 ( .A(n13246), .B(n13245), .Z(n13250) );
  NANDN U13542 ( .A(n13248), .B(n13247), .Z(n13249) );
  NAND U13543 ( .A(n13250), .B(n13249), .Z(n13376) );
  XNOR U13544 ( .A(n13377), .B(n13376), .Z(n13378) );
  NANDN U13545 ( .A(n19394), .B(n13251), .Z(n13253) );
  XOR U13546 ( .A(b[29]), .B(a[76]), .Z(n13400) );
  NANDN U13547 ( .A(n19395), .B(n13400), .Z(n13252) );
  AND U13548 ( .A(n13253), .B(n13252), .Z(n13323) );
  AND U13549 ( .A(b[31]), .B(a[72]), .Z(n13322) );
  XNOR U13550 ( .A(n13323), .B(n13322), .Z(n13324) );
  NAND U13551 ( .A(b[0]), .B(a[104]), .Z(n13254) );
  XNOR U13552 ( .A(b[1]), .B(n13254), .Z(n13256) );
  NANDN U13553 ( .A(b[0]), .B(a[103]), .Z(n13255) );
  NAND U13554 ( .A(n13256), .B(n13255), .Z(n13325) );
  XNOR U13555 ( .A(n13324), .B(n13325), .Z(n13364) );
  NANDN U13556 ( .A(n19005), .B(n13257), .Z(n13259) );
  XOR U13557 ( .A(b[23]), .B(a[82]), .Z(n13406) );
  NANDN U13558 ( .A(n19055), .B(n13406), .Z(n13258) );
  AND U13559 ( .A(n13259), .B(n13258), .Z(n13397) );
  NANDN U13560 ( .A(n17362), .B(n13260), .Z(n13262) );
  XOR U13561 ( .A(b[7]), .B(a[98]), .Z(n13409) );
  NANDN U13562 ( .A(n17522), .B(n13409), .Z(n13261) );
  AND U13563 ( .A(n13262), .B(n13261), .Z(n13395) );
  NANDN U13564 ( .A(n19116), .B(n13263), .Z(n13265) );
  XOR U13565 ( .A(b[25]), .B(a[80]), .Z(n13412) );
  NANDN U13566 ( .A(n19179), .B(n13412), .Z(n13264) );
  NAND U13567 ( .A(n13265), .B(n13264), .Z(n13394) );
  XNOR U13568 ( .A(n13395), .B(n13394), .Z(n13396) );
  XOR U13569 ( .A(n13397), .B(n13396), .Z(n13365) );
  XNOR U13570 ( .A(n13364), .B(n13365), .Z(n13366) );
  NANDN U13571 ( .A(n18113), .B(n13266), .Z(n13268) );
  XOR U13572 ( .A(b[13]), .B(a[92]), .Z(n13415) );
  NANDN U13573 ( .A(n18229), .B(n13415), .Z(n13267) );
  AND U13574 ( .A(n13268), .B(n13267), .Z(n13359) );
  NANDN U13575 ( .A(n17888), .B(n13269), .Z(n13271) );
  XOR U13576 ( .A(b[11]), .B(a[94]), .Z(n13418) );
  NANDN U13577 ( .A(n18025), .B(n13418), .Z(n13270) );
  NAND U13578 ( .A(n13271), .B(n13270), .Z(n13358) );
  XNOR U13579 ( .A(n13359), .B(n13358), .Z(n13360) );
  NANDN U13580 ( .A(n18487), .B(n13272), .Z(n13274) );
  XOR U13581 ( .A(b[15]), .B(a[90]), .Z(n13421) );
  NANDN U13582 ( .A(n18311), .B(n13421), .Z(n13273) );
  AND U13583 ( .A(n13274), .B(n13273), .Z(n13355) );
  NANDN U13584 ( .A(n18853), .B(n13275), .Z(n13277) );
  XOR U13585 ( .A(b[21]), .B(a[84]), .Z(n13424) );
  NANDN U13586 ( .A(n18926), .B(n13424), .Z(n13276) );
  AND U13587 ( .A(n13277), .B(n13276), .Z(n13353) );
  NANDN U13588 ( .A(n17613), .B(n13278), .Z(n13280) );
  XOR U13589 ( .A(b[9]), .B(a[96]), .Z(n13427) );
  NANDN U13590 ( .A(n17739), .B(n13427), .Z(n13279) );
  NAND U13591 ( .A(n13280), .B(n13279), .Z(n13352) );
  XNOR U13592 ( .A(n13353), .B(n13352), .Z(n13354) );
  XOR U13593 ( .A(n13355), .B(n13354), .Z(n13361) );
  XOR U13594 ( .A(n13360), .B(n13361), .Z(n13367) );
  XOR U13595 ( .A(n13366), .B(n13367), .Z(n13379) );
  XNOR U13596 ( .A(n13378), .B(n13379), .Z(n13310) );
  XNOR U13597 ( .A(n13311), .B(n13310), .Z(n13312) );
  XOR U13598 ( .A(n13313), .B(n13312), .Z(n13431) );
  XNOR U13599 ( .A(n13430), .B(n13431), .Z(n13432) );
  XNOR U13600 ( .A(n13433), .B(n13432), .Z(n13306) );
  XOR U13601 ( .A(n13307), .B(n13306), .Z(n13299) );
  NANDN U13602 ( .A(n13282), .B(n13281), .Z(n13286) );
  NANDN U13603 ( .A(n13284), .B(n13283), .Z(n13285) );
  AND U13604 ( .A(n13286), .B(n13285), .Z(n13298) );
  XOR U13605 ( .A(n13299), .B(n13298), .Z(n13301) );
  XNOR U13606 ( .A(n13300), .B(n13301), .Z(n13292) );
  XNOR U13607 ( .A(n13293), .B(n13292), .Z(n13294) );
  XNOR U13608 ( .A(n13295), .B(n13294), .Z(n13436) );
  XNOR U13609 ( .A(sreg[200]), .B(n13436), .Z(n13438) );
  NANDN U13610 ( .A(sreg[199]), .B(n13287), .Z(n13291) );
  NAND U13611 ( .A(n13289), .B(n13288), .Z(n13290) );
  NAND U13612 ( .A(n13291), .B(n13290), .Z(n13437) );
  XNOR U13613 ( .A(n13438), .B(n13437), .Z(c[200]) );
  NANDN U13614 ( .A(n13293), .B(n13292), .Z(n13297) );
  NANDN U13615 ( .A(n13295), .B(n13294), .Z(n13296) );
  AND U13616 ( .A(n13297), .B(n13296), .Z(n13444) );
  NANDN U13617 ( .A(n13299), .B(n13298), .Z(n13303) );
  NANDN U13618 ( .A(n13301), .B(n13300), .Z(n13302) );
  AND U13619 ( .A(n13303), .B(n13302), .Z(n13442) );
  NANDN U13620 ( .A(n13305), .B(n13304), .Z(n13309) );
  NAND U13621 ( .A(n13307), .B(n13306), .Z(n13308) );
  AND U13622 ( .A(n13309), .B(n13308), .Z(n13449) );
  NANDN U13623 ( .A(n13311), .B(n13310), .Z(n13315) );
  NANDN U13624 ( .A(n13313), .B(n13312), .Z(n13314) );
  AND U13625 ( .A(n13315), .B(n13314), .Z(n13454) );
  NANDN U13626 ( .A(n13317), .B(n13316), .Z(n13321) );
  NAND U13627 ( .A(n13319), .B(n13318), .Z(n13320) );
  AND U13628 ( .A(n13321), .B(n13320), .Z(n13453) );
  XNOR U13629 ( .A(n13454), .B(n13453), .Z(n13456) );
  NANDN U13630 ( .A(n13323), .B(n13322), .Z(n13327) );
  NANDN U13631 ( .A(n13325), .B(n13324), .Z(n13326) );
  AND U13632 ( .A(n13327), .B(n13326), .Z(n13533) );
  NANDN U13633 ( .A(n19237), .B(n13328), .Z(n13330) );
  XOR U13634 ( .A(b[27]), .B(a[79]), .Z(n13477) );
  NANDN U13635 ( .A(n19277), .B(n13477), .Z(n13329) );
  AND U13636 ( .A(n13330), .B(n13329), .Z(n13540) );
  NANDN U13637 ( .A(n17072), .B(n13331), .Z(n13333) );
  XOR U13638 ( .A(b[5]), .B(a[101]), .Z(n13480) );
  NANDN U13639 ( .A(n17223), .B(n13480), .Z(n13332) );
  AND U13640 ( .A(n13333), .B(n13332), .Z(n13538) );
  NANDN U13641 ( .A(n18673), .B(n13334), .Z(n13336) );
  XOR U13642 ( .A(b[19]), .B(a[87]), .Z(n13483) );
  NANDN U13643 ( .A(n18758), .B(n13483), .Z(n13335) );
  NAND U13644 ( .A(n13336), .B(n13335), .Z(n13537) );
  XNOR U13645 ( .A(n13538), .B(n13537), .Z(n13539) );
  XNOR U13646 ( .A(n13540), .B(n13539), .Z(n13531) );
  NANDN U13647 ( .A(n19425), .B(n13337), .Z(n13339) );
  XOR U13648 ( .A(b[31]), .B(a[75]), .Z(n13486) );
  NANDN U13649 ( .A(n19426), .B(n13486), .Z(n13338) );
  AND U13650 ( .A(n13339), .B(n13338), .Z(n13498) );
  NANDN U13651 ( .A(n17067), .B(n13340), .Z(n13342) );
  XOR U13652 ( .A(a[103]), .B(b[3]), .Z(n13489) );
  NANDN U13653 ( .A(n17068), .B(n13489), .Z(n13341) );
  AND U13654 ( .A(n13342), .B(n13341), .Z(n13496) );
  NANDN U13655 ( .A(n18514), .B(n13343), .Z(n13345) );
  XOR U13656 ( .A(b[17]), .B(a[89]), .Z(n13492) );
  NANDN U13657 ( .A(n18585), .B(n13492), .Z(n13344) );
  NAND U13658 ( .A(n13345), .B(n13344), .Z(n13495) );
  XNOR U13659 ( .A(n13496), .B(n13495), .Z(n13497) );
  XOR U13660 ( .A(n13498), .B(n13497), .Z(n13532) );
  XOR U13661 ( .A(n13531), .B(n13532), .Z(n13534) );
  XOR U13662 ( .A(n13533), .B(n13534), .Z(n13466) );
  NANDN U13663 ( .A(n13347), .B(n13346), .Z(n13351) );
  NANDN U13664 ( .A(n13349), .B(n13348), .Z(n13350) );
  AND U13665 ( .A(n13351), .B(n13350), .Z(n13519) );
  NANDN U13666 ( .A(n13353), .B(n13352), .Z(n13357) );
  NANDN U13667 ( .A(n13355), .B(n13354), .Z(n13356) );
  NAND U13668 ( .A(n13357), .B(n13356), .Z(n13520) );
  XNOR U13669 ( .A(n13519), .B(n13520), .Z(n13521) );
  NANDN U13670 ( .A(n13359), .B(n13358), .Z(n13363) );
  NANDN U13671 ( .A(n13361), .B(n13360), .Z(n13362) );
  NAND U13672 ( .A(n13363), .B(n13362), .Z(n13522) );
  XNOR U13673 ( .A(n13521), .B(n13522), .Z(n13465) );
  XNOR U13674 ( .A(n13466), .B(n13465), .Z(n13468) );
  NANDN U13675 ( .A(n13365), .B(n13364), .Z(n13369) );
  NANDN U13676 ( .A(n13367), .B(n13366), .Z(n13368) );
  AND U13677 ( .A(n13369), .B(n13368), .Z(n13467) );
  XOR U13678 ( .A(n13468), .B(n13467), .Z(n13582) );
  NANDN U13679 ( .A(n13371), .B(n13370), .Z(n13375) );
  NANDN U13680 ( .A(n13373), .B(n13372), .Z(n13374) );
  AND U13681 ( .A(n13375), .B(n13374), .Z(n13579) );
  NANDN U13682 ( .A(n13377), .B(n13376), .Z(n13381) );
  NANDN U13683 ( .A(n13379), .B(n13378), .Z(n13380) );
  AND U13684 ( .A(n13381), .B(n13380), .Z(n13462) );
  NANDN U13685 ( .A(n13383), .B(n13382), .Z(n13387) );
  OR U13686 ( .A(n13385), .B(n13384), .Z(n13386) );
  AND U13687 ( .A(n13387), .B(n13386), .Z(n13460) );
  NANDN U13688 ( .A(n13389), .B(n13388), .Z(n13393) );
  NANDN U13689 ( .A(n13391), .B(n13390), .Z(n13392) );
  AND U13690 ( .A(n13393), .B(n13392), .Z(n13526) );
  NANDN U13691 ( .A(n13395), .B(n13394), .Z(n13399) );
  NANDN U13692 ( .A(n13397), .B(n13396), .Z(n13398) );
  NAND U13693 ( .A(n13399), .B(n13398), .Z(n13525) );
  XNOR U13694 ( .A(n13526), .B(n13525), .Z(n13527) );
  NANDN U13695 ( .A(n19394), .B(n13400), .Z(n13402) );
  XOR U13696 ( .A(b[29]), .B(a[77]), .Z(n13552) );
  NANDN U13697 ( .A(n19395), .B(n13552), .Z(n13401) );
  AND U13698 ( .A(n13402), .B(n13401), .Z(n13472) );
  AND U13699 ( .A(b[31]), .B(a[73]), .Z(n13471) );
  XNOR U13700 ( .A(n13472), .B(n13471), .Z(n13473) );
  NAND U13701 ( .A(b[0]), .B(a[105]), .Z(n13403) );
  XNOR U13702 ( .A(b[1]), .B(n13403), .Z(n13405) );
  NANDN U13703 ( .A(b[0]), .B(a[104]), .Z(n13404) );
  NAND U13704 ( .A(n13405), .B(n13404), .Z(n13474) );
  XNOR U13705 ( .A(n13473), .B(n13474), .Z(n13513) );
  NANDN U13706 ( .A(n19005), .B(n13406), .Z(n13408) );
  XOR U13707 ( .A(b[23]), .B(a[83]), .Z(n13555) );
  NANDN U13708 ( .A(n19055), .B(n13555), .Z(n13407) );
  AND U13709 ( .A(n13408), .B(n13407), .Z(n13546) );
  NANDN U13710 ( .A(n17362), .B(n13409), .Z(n13411) );
  XOR U13711 ( .A(b[7]), .B(a[99]), .Z(n13558) );
  NANDN U13712 ( .A(n17522), .B(n13558), .Z(n13410) );
  AND U13713 ( .A(n13411), .B(n13410), .Z(n13544) );
  NANDN U13714 ( .A(n19116), .B(n13412), .Z(n13414) );
  XOR U13715 ( .A(b[25]), .B(a[81]), .Z(n13561) );
  NANDN U13716 ( .A(n19179), .B(n13561), .Z(n13413) );
  NAND U13717 ( .A(n13414), .B(n13413), .Z(n13543) );
  XNOR U13718 ( .A(n13544), .B(n13543), .Z(n13545) );
  XOR U13719 ( .A(n13546), .B(n13545), .Z(n13514) );
  XNOR U13720 ( .A(n13513), .B(n13514), .Z(n13515) );
  NANDN U13721 ( .A(n18113), .B(n13415), .Z(n13417) );
  XOR U13722 ( .A(b[13]), .B(a[93]), .Z(n13564) );
  NANDN U13723 ( .A(n18229), .B(n13564), .Z(n13416) );
  AND U13724 ( .A(n13417), .B(n13416), .Z(n13508) );
  NANDN U13725 ( .A(n17888), .B(n13418), .Z(n13420) );
  XOR U13726 ( .A(b[11]), .B(a[95]), .Z(n13567) );
  NANDN U13727 ( .A(n18025), .B(n13567), .Z(n13419) );
  NAND U13728 ( .A(n13420), .B(n13419), .Z(n13507) );
  XNOR U13729 ( .A(n13508), .B(n13507), .Z(n13509) );
  NANDN U13730 ( .A(n18487), .B(n13421), .Z(n13423) );
  XOR U13731 ( .A(b[15]), .B(a[91]), .Z(n13570) );
  NANDN U13732 ( .A(n18311), .B(n13570), .Z(n13422) );
  AND U13733 ( .A(n13423), .B(n13422), .Z(n13504) );
  NANDN U13734 ( .A(n18853), .B(n13424), .Z(n13426) );
  XOR U13735 ( .A(b[21]), .B(a[85]), .Z(n13573) );
  NANDN U13736 ( .A(n18926), .B(n13573), .Z(n13425) );
  AND U13737 ( .A(n13426), .B(n13425), .Z(n13502) );
  NANDN U13738 ( .A(n17613), .B(n13427), .Z(n13429) );
  XOR U13739 ( .A(b[9]), .B(a[97]), .Z(n13576) );
  NANDN U13740 ( .A(n17739), .B(n13576), .Z(n13428) );
  NAND U13741 ( .A(n13429), .B(n13428), .Z(n13501) );
  XNOR U13742 ( .A(n13502), .B(n13501), .Z(n13503) );
  XOR U13743 ( .A(n13504), .B(n13503), .Z(n13510) );
  XOR U13744 ( .A(n13509), .B(n13510), .Z(n13516) );
  XOR U13745 ( .A(n13515), .B(n13516), .Z(n13528) );
  XNOR U13746 ( .A(n13527), .B(n13528), .Z(n13459) );
  XNOR U13747 ( .A(n13460), .B(n13459), .Z(n13461) );
  XOR U13748 ( .A(n13462), .B(n13461), .Z(n13580) );
  XNOR U13749 ( .A(n13579), .B(n13580), .Z(n13581) );
  XNOR U13750 ( .A(n13582), .B(n13581), .Z(n13455) );
  XOR U13751 ( .A(n13456), .B(n13455), .Z(n13448) );
  NANDN U13752 ( .A(n13431), .B(n13430), .Z(n13435) );
  NANDN U13753 ( .A(n13433), .B(n13432), .Z(n13434) );
  AND U13754 ( .A(n13435), .B(n13434), .Z(n13447) );
  XOR U13755 ( .A(n13448), .B(n13447), .Z(n13450) );
  XNOR U13756 ( .A(n13449), .B(n13450), .Z(n13441) );
  XNOR U13757 ( .A(n13442), .B(n13441), .Z(n13443) );
  XNOR U13758 ( .A(n13444), .B(n13443), .Z(n13585) );
  XNOR U13759 ( .A(sreg[201]), .B(n13585), .Z(n13587) );
  NANDN U13760 ( .A(sreg[200]), .B(n13436), .Z(n13440) );
  NAND U13761 ( .A(n13438), .B(n13437), .Z(n13439) );
  NAND U13762 ( .A(n13440), .B(n13439), .Z(n13586) );
  XNOR U13763 ( .A(n13587), .B(n13586), .Z(c[201]) );
  NANDN U13764 ( .A(n13442), .B(n13441), .Z(n13446) );
  NANDN U13765 ( .A(n13444), .B(n13443), .Z(n13445) );
  AND U13766 ( .A(n13446), .B(n13445), .Z(n13593) );
  NANDN U13767 ( .A(n13448), .B(n13447), .Z(n13452) );
  NANDN U13768 ( .A(n13450), .B(n13449), .Z(n13451) );
  AND U13769 ( .A(n13452), .B(n13451), .Z(n13591) );
  NANDN U13770 ( .A(n13454), .B(n13453), .Z(n13458) );
  NAND U13771 ( .A(n13456), .B(n13455), .Z(n13457) );
  AND U13772 ( .A(n13458), .B(n13457), .Z(n13598) );
  NANDN U13773 ( .A(n13460), .B(n13459), .Z(n13464) );
  NANDN U13774 ( .A(n13462), .B(n13461), .Z(n13463) );
  AND U13775 ( .A(n13464), .B(n13463), .Z(n13603) );
  NANDN U13776 ( .A(n13466), .B(n13465), .Z(n13470) );
  NAND U13777 ( .A(n13468), .B(n13467), .Z(n13469) );
  AND U13778 ( .A(n13470), .B(n13469), .Z(n13602) );
  XNOR U13779 ( .A(n13603), .B(n13602), .Z(n13605) );
  NANDN U13780 ( .A(n13472), .B(n13471), .Z(n13476) );
  NANDN U13781 ( .A(n13474), .B(n13473), .Z(n13475) );
  AND U13782 ( .A(n13476), .B(n13475), .Z(n13682) );
  NANDN U13783 ( .A(n19237), .B(n13477), .Z(n13479) );
  XOR U13784 ( .A(b[27]), .B(a[80]), .Z(n13626) );
  NANDN U13785 ( .A(n19277), .B(n13626), .Z(n13478) );
  AND U13786 ( .A(n13479), .B(n13478), .Z(n13689) );
  NANDN U13787 ( .A(n17072), .B(n13480), .Z(n13482) );
  XOR U13788 ( .A(b[5]), .B(a[102]), .Z(n13629) );
  NANDN U13789 ( .A(n17223), .B(n13629), .Z(n13481) );
  AND U13790 ( .A(n13482), .B(n13481), .Z(n13687) );
  NANDN U13791 ( .A(n18673), .B(n13483), .Z(n13485) );
  XOR U13792 ( .A(b[19]), .B(a[88]), .Z(n13632) );
  NANDN U13793 ( .A(n18758), .B(n13632), .Z(n13484) );
  NAND U13794 ( .A(n13485), .B(n13484), .Z(n13686) );
  XNOR U13795 ( .A(n13687), .B(n13686), .Z(n13688) );
  XNOR U13796 ( .A(n13689), .B(n13688), .Z(n13680) );
  NANDN U13797 ( .A(n19425), .B(n13486), .Z(n13488) );
  XOR U13798 ( .A(b[31]), .B(a[76]), .Z(n13635) );
  NANDN U13799 ( .A(n19426), .B(n13635), .Z(n13487) );
  AND U13800 ( .A(n13488), .B(n13487), .Z(n13647) );
  NANDN U13801 ( .A(n17067), .B(n13489), .Z(n13491) );
  XOR U13802 ( .A(a[104]), .B(b[3]), .Z(n13638) );
  NANDN U13803 ( .A(n17068), .B(n13638), .Z(n13490) );
  AND U13804 ( .A(n13491), .B(n13490), .Z(n13645) );
  NANDN U13805 ( .A(n18514), .B(n13492), .Z(n13494) );
  XOR U13806 ( .A(b[17]), .B(a[90]), .Z(n13641) );
  NANDN U13807 ( .A(n18585), .B(n13641), .Z(n13493) );
  NAND U13808 ( .A(n13494), .B(n13493), .Z(n13644) );
  XNOR U13809 ( .A(n13645), .B(n13644), .Z(n13646) );
  XOR U13810 ( .A(n13647), .B(n13646), .Z(n13681) );
  XOR U13811 ( .A(n13680), .B(n13681), .Z(n13683) );
  XOR U13812 ( .A(n13682), .B(n13683), .Z(n13615) );
  NANDN U13813 ( .A(n13496), .B(n13495), .Z(n13500) );
  NANDN U13814 ( .A(n13498), .B(n13497), .Z(n13499) );
  AND U13815 ( .A(n13500), .B(n13499), .Z(n13668) );
  NANDN U13816 ( .A(n13502), .B(n13501), .Z(n13506) );
  NANDN U13817 ( .A(n13504), .B(n13503), .Z(n13505) );
  NAND U13818 ( .A(n13506), .B(n13505), .Z(n13669) );
  XNOR U13819 ( .A(n13668), .B(n13669), .Z(n13670) );
  NANDN U13820 ( .A(n13508), .B(n13507), .Z(n13512) );
  NANDN U13821 ( .A(n13510), .B(n13509), .Z(n13511) );
  NAND U13822 ( .A(n13512), .B(n13511), .Z(n13671) );
  XNOR U13823 ( .A(n13670), .B(n13671), .Z(n13614) );
  XNOR U13824 ( .A(n13615), .B(n13614), .Z(n13617) );
  NANDN U13825 ( .A(n13514), .B(n13513), .Z(n13518) );
  NANDN U13826 ( .A(n13516), .B(n13515), .Z(n13517) );
  AND U13827 ( .A(n13518), .B(n13517), .Z(n13616) );
  XOR U13828 ( .A(n13617), .B(n13616), .Z(n13731) );
  NANDN U13829 ( .A(n13520), .B(n13519), .Z(n13524) );
  NANDN U13830 ( .A(n13522), .B(n13521), .Z(n13523) );
  AND U13831 ( .A(n13524), .B(n13523), .Z(n13728) );
  NANDN U13832 ( .A(n13526), .B(n13525), .Z(n13530) );
  NANDN U13833 ( .A(n13528), .B(n13527), .Z(n13529) );
  AND U13834 ( .A(n13530), .B(n13529), .Z(n13611) );
  NANDN U13835 ( .A(n13532), .B(n13531), .Z(n13536) );
  OR U13836 ( .A(n13534), .B(n13533), .Z(n13535) );
  AND U13837 ( .A(n13536), .B(n13535), .Z(n13609) );
  NANDN U13838 ( .A(n13538), .B(n13537), .Z(n13542) );
  NANDN U13839 ( .A(n13540), .B(n13539), .Z(n13541) );
  AND U13840 ( .A(n13542), .B(n13541), .Z(n13675) );
  NANDN U13841 ( .A(n13544), .B(n13543), .Z(n13548) );
  NANDN U13842 ( .A(n13546), .B(n13545), .Z(n13547) );
  NAND U13843 ( .A(n13548), .B(n13547), .Z(n13674) );
  XNOR U13844 ( .A(n13675), .B(n13674), .Z(n13676) );
  NAND U13845 ( .A(b[0]), .B(a[106]), .Z(n13549) );
  XNOR U13846 ( .A(b[1]), .B(n13549), .Z(n13551) );
  NANDN U13847 ( .A(b[0]), .B(a[105]), .Z(n13550) );
  NAND U13848 ( .A(n13551), .B(n13550), .Z(n13623) );
  NANDN U13849 ( .A(n19394), .B(n13552), .Z(n13554) );
  XOR U13850 ( .A(b[29]), .B(a[78]), .Z(n13701) );
  NANDN U13851 ( .A(n19395), .B(n13701), .Z(n13553) );
  AND U13852 ( .A(n13554), .B(n13553), .Z(n13621) );
  AND U13853 ( .A(b[31]), .B(a[74]), .Z(n13620) );
  XNOR U13854 ( .A(n13621), .B(n13620), .Z(n13622) );
  XNOR U13855 ( .A(n13623), .B(n13622), .Z(n13662) );
  NANDN U13856 ( .A(n19005), .B(n13555), .Z(n13557) );
  XOR U13857 ( .A(b[23]), .B(a[84]), .Z(n13704) );
  NANDN U13858 ( .A(n19055), .B(n13704), .Z(n13556) );
  AND U13859 ( .A(n13557), .B(n13556), .Z(n13695) );
  NANDN U13860 ( .A(n17362), .B(n13558), .Z(n13560) );
  XOR U13861 ( .A(b[7]), .B(a[100]), .Z(n13707) );
  NANDN U13862 ( .A(n17522), .B(n13707), .Z(n13559) );
  AND U13863 ( .A(n13560), .B(n13559), .Z(n13693) );
  NANDN U13864 ( .A(n19116), .B(n13561), .Z(n13563) );
  XOR U13865 ( .A(b[25]), .B(a[82]), .Z(n13710) );
  NANDN U13866 ( .A(n19179), .B(n13710), .Z(n13562) );
  NAND U13867 ( .A(n13563), .B(n13562), .Z(n13692) );
  XNOR U13868 ( .A(n13693), .B(n13692), .Z(n13694) );
  XOR U13869 ( .A(n13695), .B(n13694), .Z(n13663) );
  XNOR U13870 ( .A(n13662), .B(n13663), .Z(n13664) );
  NANDN U13871 ( .A(n18113), .B(n13564), .Z(n13566) );
  XOR U13872 ( .A(b[13]), .B(a[94]), .Z(n13713) );
  NANDN U13873 ( .A(n18229), .B(n13713), .Z(n13565) );
  AND U13874 ( .A(n13566), .B(n13565), .Z(n13657) );
  NANDN U13875 ( .A(n17888), .B(n13567), .Z(n13569) );
  XOR U13876 ( .A(b[11]), .B(a[96]), .Z(n13716) );
  NANDN U13877 ( .A(n18025), .B(n13716), .Z(n13568) );
  NAND U13878 ( .A(n13569), .B(n13568), .Z(n13656) );
  XNOR U13879 ( .A(n13657), .B(n13656), .Z(n13658) );
  NANDN U13880 ( .A(n18487), .B(n13570), .Z(n13572) );
  XOR U13881 ( .A(b[15]), .B(a[92]), .Z(n13719) );
  NANDN U13882 ( .A(n18311), .B(n13719), .Z(n13571) );
  AND U13883 ( .A(n13572), .B(n13571), .Z(n13653) );
  NANDN U13884 ( .A(n18853), .B(n13573), .Z(n13575) );
  XOR U13885 ( .A(b[21]), .B(a[86]), .Z(n13722) );
  NANDN U13886 ( .A(n18926), .B(n13722), .Z(n13574) );
  AND U13887 ( .A(n13575), .B(n13574), .Z(n13651) );
  NANDN U13888 ( .A(n17613), .B(n13576), .Z(n13578) );
  XOR U13889 ( .A(b[9]), .B(a[98]), .Z(n13725) );
  NANDN U13890 ( .A(n17739), .B(n13725), .Z(n13577) );
  NAND U13891 ( .A(n13578), .B(n13577), .Z(n13650) );
  XNOR U13892 ( .A(n13651), .B(n13650), .Z(n13652) );
  XOR U13893 ( .A(n13653), .B(n13652), .Z(n13659) );
  XOR U13894 ( .A(n13658), .B(n13659), .Z(n13665) );
  XOR U13895 ( .A(n13664), .B(n13665), .Z(n13677) );
  XNOR U13896 ( .A(n13676), .B(n13677), .Z(n13608) );
  XNOR U13897 ( .A(n13609), .B(n13608), .Z(n13610) );
  XOR U13898 ( .A(n13611), .B(n13610), .Z(n13729) );
  XNOR U13899 ( .A(n13728), .B(n13729), .Z(n13730) );
  XNOR U13900 ( .A(n13731), .B(n13730), .Z(n13604) );
  XOR U13901 ( .A(n13605), .B(n13604), .Z(n13597) );
  NANDN U13902 ( .A(n13580), .B(n13579), .Z(n13584) );
  NANDN U13903 ( .A(n13582), .B(n13581), .Z(n13583) );
  AND U13904 ( .A(n13584), .B(n13583), .Z(n13596) );
  XOR U13905 ( .A(n13597), .B(n13596), .Z(n13599) );
  XNOR U13906 ( .A(n13598), .B(n13599), .Z(n13590) );
  XNOR U13907 ( .A(n13591), .B(n13590), .Z(n13592) );
  XNOR U13908 ( .A(n13593), .B(n13592), .Z(n13734) );
  XNOR U13909 ( .A(sreg[202]), .B(n13734), .Z(n13736) );
  NANDN U13910 ( .A(sreg[201]), .B(n13585), .Z(n13589) );
  NAND U13911 ( .A(n13587), .B(n13586), .Z(n13588) );
  NAND U13912 ( .A(n13589), .B(n13588), .Z(n13735) );
  XNOR U13913 ( .A(n13736), .B(n13735), .Z(c[202]) );
  NANDN U13914 ( .A(n13591), .B(n13590), .Z(n13595) );
  NANDN U13915 ( .A(n13593), .B(n13592), .Z(n13594) );
  AND U13916 ( .A(n13595), .B(n13594), .Z(n13742) );
  NANDN U13917 ( .A(n13597), .B(n13596), .Z(n13601) );
  NANDN U13918 ( .A(n13599), .B(n13598), .Z(n13600) );
  AND U13919 ( .A(n13601), .B(n13600), .Z(n13740) );
  NANDN U13920 ( .A(n13603), .B(n13602), .Z(n13607) );
  NAND U13921 ( .A(n13605), .B(n13604), .Z(n13606) );
  AND U13922 ( .A(n13607), .B(n13606), .Z(n13747) );
  NANDN U13923 ( .A(n13609), .B(n13608), .Z(n13613) );
  NANDN U13924 ( .A(n13611), .B(n13610), .Z(n13612) );
  AND U13925 ( .A(n13613), .B(n13612), .Z(n13876) );
  NANDN U13926 ( .A(n13615), .B(n13614), .Z(n13619) );
  NAND U13927 ( .A(n13617), .B(n13616), .Z(n13618) );
  AND U13928 ( .A(n13619), .B(n13618), .Z(n13875) );
  XNOR U13929 ( .A(n13876), .B(n13875), .Z(n13878) );
  NANDN U13930 ( .A(n13621), .B(n13620), .Z(n13625) );
  NANDN U13931 ( .A(n13623), .B(n13622), .Z(n13624) );
  AND U13932 ( .A(n13625), .B(n13624), .Z(n13823) );
  NANDN U13933 ( .A(n19237), .B(n13626), .Z(n13628) );
  XOR U13934 ( .A(b[27]), .B(a[81]), .Z(n13769) );
  NANDN U13935 ( .A(n19277), .B(n13769), .Z(n13627) );
  AND U13936 ( .A(n13628), .B(n13627), .Z(n13830) );
  NANDN U13937 ( .A(n17072), .B(n13629), .Z(n13631) );
  XOR U13938 ( .A(b[5]), .B(a[103]), .Z(n13772) );
  NANDN U13939 ( .A(n17223), .B(n13772), .Z(n13630) );
  AND U13940 ( .A(n13631), .B(n13630), .Z(n13828) );
  NANDN U13941 ( .A(n18673), .B(n13632), .Z(n13634) );
  XOR U13942 ( .A(b[19]), .B(a[89]), .Z(n13775) );
  NANDN U13943 ( .A(n18758), .B(n13775), .Z(n13633) );
  NAND U13944 ( .A(n13634), .B(n13633), .Z(n13827) );
  XNOR U13945 ( .A(n13828), .B(n13827), .Z(n13829) );
  XNOR U13946 ( .A(n13830), .B(n13829), .Z(n13821) );
  NANDN U13947 ( .A(n19425), .B(n13635), .Z(n13637) );
  XOR U13948 ( .A(b[31]), .B(a[77]), .Z(n13778) );
  NANDN U13949 ( .A(n19426), .B(n13778), .Z(n13636) );
  AND U13950 ( .A(n13637), .B(n13636), .Z(n13790) );
  NANDN U13951 ( .A(n17067), .B(n13638), .Z(n13640) );
  XOR U13952 ( .A(a[105]), .B(b[3]), .Z(n13781) );
  NANDN U13953 ( .A(n17068), .B(n13781), .Z(n13639) );
  AND U13954 ( .A(n13640), .B(n13639), .Z(n13788) );
  NANDN U13955 ( .A(n18514), .B(n13641), .Z(n13643) );
  XOR U13956 ( .A(b[17]), .B(a[91]), .Z(n13784) );
  NANDN U13957 ( .A(n18585), .B(n13784), .Z(n13642) );
  NAND U13958 ( .A(n13643), .B(n13642), .Z(n13787) );
  XNOR U13959 ( .A(n13788), .B(n13787), .Z(n13789) );
  XOR U13960 ( .A(n13790), .B(n13789), .Z(n13822) );
  XOR U13961 ( .A(n13821), .B(n13822), .Z(n13824) );
  XOR U13962 ( .A(n13823), .B(n13824), .Z(n13758) );
  NANDN U13963 ( .A(n13645), .B(n13644), .Z(n13649) );
  NANDN U13964 ( .A(n13647), .B(n13646), .Z(n13648) );
  AND U13965 ( .A(n13649), .B(n13648), .Z(n13811) );
  NANDN U13966 ( .A(n13651), .B(n13650), .Z(n13655) );
  NANDN U13967 ( .A(n13653), .B(n13652), .Z(n13654) );
  NAND U13968 ( .A(n13655), .B(n13654), .Z(n13812) );
  XNOR U13969 ( .A(n13811), .B(n13812), .Z(n13813) );
  NANDN U13970 ( .A(n13657), .B(n13656), .Z(n13661) );
  NANDN U13971 ( .A(n13659), .B(n13658), .Z(n13660) );
  NAND U13972 ( .A(n13661), .B(n13660), .Z(n13814) );
  XNOR U13973 ( .A(n13813), .B(n13814), .Z(n13757) );
  XNOR U13974 ( .A(n13758), .B(n13757), .Z(n13760) );
  NANDN U13975 ( .A(n13663), .B(n13662), .Z(n13667) );
  NANDN U13976 ( .A(n13665), .B(n13664), .Z(n13666) );
  AND U13977 ( .A(n13667), .B(n13666), .Z(n13759) );
  XOR U13978 ( .A(n13760), .B(n13759), .Z(n13872) );
  NANDN U13979 ( .A(n13669), .B(n13668), .Z(n13673) );
  NANDN U13980 ( .A(n13671), .B(n13670), .Z(n13672) );
  AND U13981 ( .A(n13673), .B(n13672), .Z(n13869) );
  NANDN U13982 ( .A(n13675), .B(n13674), .Z(n13679) );
  NANDN U13983 ( .A(n13677), .B(n13676), .Z(n13678) );
  AND U13984 ( .A(n13679), .B(n13678), .Z(n13754) );
  NANDN U13985 ( .A(n13681), .B(n13680), .Z(n13685) );
  OR U13986 ( .A(n13683), .B(n13682), .Z(n13684) );
  AND U13987 ( .A(n13685), .B(n13684), .Z(n13752) );
  NANDN U13988 ( .A(n13687), .B(n13686), .Z(n13691) );
  NANDN U13989 ( .A(n13689), .B(n13688), .Z(n13690) );
  AND U13990 ( .A(n13691), .B(n13690), .Z(n13818) );
  NANDN U13991 ( .A(n13693), .B(n13692), .Z(n13697) );
  NANDN U13992 ( .A(n13695), .B(n13694), .Z(n13696) );
  NAND U13993 ( .A(n13697), .B(n13696), .Z(n13817) );
  XNOR U13994 ( .A(n13818), .B(n13817), .Z(n13820) );
  NAND U13995 ( .A(b[0]), .B(a[107]), .Z(n13698) );
  XNOR U13996 ( .A(b[1]), .B(n13698), .Z(n13700) );
  NANDN U13997 ( .A(b[0]), .B(a[106]), .Z(n13699) );
  NAND U13998 ( .A(n13700), .B(n13699), .Z(n13766) );
  NANDN U13999 ( .A(n19394), .B(n13701), .Z(n13703) );
  XOR U14000 ( .A(b[29]), .B(a[79]), .Z(n13842) );
  NANDN U14001 ( .A(n19395), .B(n13842), .Z(n13702) );
  AND U14002 ( .A(n13703), .B(n13702), .Z(n13764) );
  AND U14003 ( .A(b[31]), .B(a[75]), .Z(n13763) );
  XNOR U14004 ( .A(n13764), .B(n13763), .Z(n13765) );
  XNOR U14005 ( .A(n13766), .B(n13765), .Z(n13806) );
  NANDN U14006 ( .A(n19005), .B(n13704), .Z(n13706) );
  XOR U14007 ( .A(b[23]), .B(a[85]), .Z(n13845) );
  NANDN U14008 ( .A(n19055), .B(n13845), .Z(n13705) );
  AND U14009 ( .A(n13706), .B(n13705), .Z(n13835) );
  NANDN U14010 ( .A(n17362), .B(n13707), .Z(n13709) );
  XOR U14011 ( .A(b[7]), .B(a[101]), .Z(n13848) );
  NANDN U14012 ( .A(n17522), .B(n13848), .Z(n13708) );
  AND U14013 ( .A(n13709), .B(n13708), .Z(n13834) );
  NANDN U14014 ( .A(n19116), .B(n13710), .Z(n13712) );
  XOR U14015 ( .A(b[25]), .B(a[83]), .Z(n13851) );
  NANDN U14016 ( .A(n19179), .B(n13851), .Z(n13711) );
  NAND U14017 ( .A(n13712), .B(n13711), .Z(n13833) );
  XOR U14018 ( .A(n13834), .B(n13833), .Z(n13836) );
  XOR U14019 ( .A(n13835), .B(n13836), .Z(n13805) );
  XOR U14020 ( .A(n13806), .B(n13805), .Z(n13808) );
  NANDN U14021 ( .A(n18113), .B(n13713), .Z(n13715) );
  XOR U14022 ( .A(b[13]), .B(a[95]), .Z(n13854) );
  NANDN U14023 ( .A(n18229), .B(n13854), .Z(n13714) );
  AND U14024 ( .A(n13715), .B(n13714), .Z(n13800) );
  NANDN U14025 ( .A(n17888), .B(n13716), .Z(n13718) );
  XOR U14026 ( .A(b[11]), .B(a[97]), .Z(n13857) );
  NANDN U14027 ( .A(n18025), .B(n13857), .Z(n13717) );
  NAND U14028 ( .A(n13718), .B(n13717), .Z(n13799) );
  XNOR U14029 ( .A(n13800), .B(n13799), .Z(n13802) );
  NANDN U14030 ( .A(n18487), .B(n13719), .Z(n13721) );
  XOR U14031 ( .A(b[15]), .B(a[93]), .Z(n13860) );
  NANDN U14032 ( .A(n18311), .B(n13860), .Z(n13720) );
  AND U14033 ( .A(n13721), .B(n13720), .Z(n13796) );
  NANDN U14034 ( .A(n18853), .B(n13722), .Z(n13724) );
  XOR U14035 ( .A(b[21]), .B(a[87]), .Z(n13863) );
  NANDN U14036 ( .A(n18926), .B(n13863), .Z(n13723) );
  AND U14037 ( .A(n13724), .B(n13723), .Z(n13794) );
  NANDN U14038 ( .A(n17613), .B(n13725), .Z(n13727) );
  XOR U14039 ( .A(b[9]), .B(a[99]), .Z(n13866) );
  NANDN U14040 ( .A(n17739), .B(n13866), .Z(n13726) );
  NAND U14041 ( .A(n13727), .B(n13726), .Z(n13793) );
  XNOR U14042 ( .A(n13794), .B(n13793), .Z(n13795) );
  XNOR U14043 ( .A(n13796), .B(n13795), .Z(n13801) );
  XOR U14044 ( .A(n13802), .B(n13801), .Z(n13807) );
  XOR U14045 ( .A(n13808), .B(n13807), .Z(n13819) );
  XOR U14046 ( .A(n13820), .B(n13819), .Z(n13751) );
  XNOR U14047 ( .A(n13752), .B(n13751), .Z(n13753) );
  XOR U14048 ( .A(n13754), .B(n13753), .Z(n13870) );
  XNOR U14049 ( .A(n13869), .B(n13870), .Z(n13871) );
  XNOR U14050 ( .A(n13872), .B(n13871), .Z(n13877) );
  XOR U14051 ( .A(n13878), .B(n13877), .Z(n13746) );
  NANDN U14052 ( .A(n13729), .B(n13728), .Z(n13733) );
  NANDN U14053 ( .A(n13731), .B(n13730), .Z(n13732) );
  AND U14054 ( .A(n13733), .B(n13732), .Z(n13745) );
  XOR U14055 ( .A(n13746), .B(n13745), .Z(n13748) );
  XNOR U14056 ( .A(n13747), .B(n13748), .Z(n13739) );
  XNOR U14057 ( .A(n13740), .B(n13739), .Z(n13741) );
  XNOR U14058 ( .A(n13742), .B(n13741), .Z(n13881) );
  XNOR U14059 ( .A(sreg[203]), .B(n13881), .Z(n13883) );
  NANDN U14060 ( .A(sreg[202]), .B(n13734), .Z(n13738) );
  NAND U14061 ( .A(n13736), .B(n13735), .Z(n13737) );
  NAND U14062 ( .A(n13738), .B(n13737), .Z(n13882) );
  XNOR U14063 ( .A(n13883), .B(n13882), .Z(c[203]) );
  NANDN U14064 ( .A(n13740), .B(n13739), .Z(n13744) );
  NANDN U14065 ( .A(n13742), .B(n13741), .Z(n13743) );
  AND U14066 ( .A(n13744), .B(n13743), .Z(n13889) );
  NANDN U14067 ( .A(n13746), .B(n13745), .Z(n13750) );
  NANDN U14068 ( .A(n13748), .B(n13747), .Z(n13749) );
  AND U14069 ( .A(n13750), .B(n13749), .Z(n13887) );
  NANDN U14070 ( .A(n13752), .B(n13751), .Z(n13756) );
  NANDN U14071 ( .A(n13754), .B(n13753), .Z(n13755) );
  AND U14072 ( .A(n13756), .B(n13755), .Z(n14025) );
  NANDN U14073 ( .A(n13758), .B(n13757), .Z(n13762) );
  NAND U14074 ( .A(n13760), .B(n13759), .Z(n13761) );
  AND U14075 ( .A(n13762), .B(n13761), .Z(n14024) );
  XNOR U14076 ( .A(n14025), .B(n14024), .Z(n14027) );
  NANDN U14077 ( .A(n13764), .B(n13763), .Z(n13768) );
  NANDN U14078 ( .A(n13766), .B(n13765), .Z(n13767) );
  AND U14079 ( .A(n13768), .B(n13767), .Z(n13960) );
  NANDN U14080 ( .A(n19237), .B(n13769), .Z(n13771) );
  XOR U14081 ( .A(b[27]), .B(a[82]), .Z(n13904) );
  NANDN U14082 ( .A(n19277), .B(n13904), .Z(n13770) );
  AND U14083 ( .A(n13771), .B(n13770), .Z(n13967) );
  NANDN U14084 ( .A(n17072), .B(n13772), .Z(n13774) );
  XOR U14085 ( .A(a[104]), .B(b[5]), .Z(n13907) );
  NANDN U14086 ( .A(n17223), .B(n13907), .Z(n13773) );
  AND U14087 ( .A(n13774), .B(n13773), .Z(n13965) );
  NANDN U14088 ( .A(n18673), .B(n13775), .Z(n13777) );
  XOR U14089 ( .A(b[19]), .B(a[90]), .Z(n13910) );
  NANDN U14090 ( .A(n18758), .B(n13910), .Z(n13776) );
  NAND U14091 ( .A(n13777), .B(n13776), .Z(n13964) );
  XNOR U14092 ( .A(n13965), .B(n13964), .Z(n13966) );
  XNOR U14093 ( .A(n13967), .B(n13966), .Z(n13958) );
  NANDN U14094 ( .A(n19425), .B(n13778), .Z(n13780) );
  XOR U14095 ( .A(b[31]), .B(a[78]), .Z(n13913) );
  NANDN U14096 ( .A(n19426), .B(n13913), .Z(n13779) );
  AND U14097 ( .A(n13780), .B(n13779), .Z(n13925) );
  NANDN U14098 ( .A(n17067), .B(n13781), .Z(n13783) );
  XOR U14099 ( .A(a[106]), .B(b[3]), .Z(n13916) );
  NANDN U14100 ( .A(n17068), .B(n13916), .Z(n13782) );
  AND U14101 ( .A(n13783), .B(n13782), .Z(n13923) );
  NANDN U14102 ( .A(n18514), .B(n13784), .Z(n13786) );
  XOR U14103 ( .A(b[17]), .B(a[92]), .Z(n13919) );
  NANDN U14104 ( .A(n18585), .B(n13919), .Z(n13785) );
  NAND U14105 ( .A(n13786), .B(n13785), .Z(n13922) );
  XNOR U14106 ( .A(n13923), .B(n13922), .Z(n13924) );
  XOR U14107 ( .A(n13925), .B(n13924), .Z(n13959) );
  XOR U14108 ( .A(n13958), .B(n13959), .Z(n13961) );
  XOR U14109 ( .A(n13960), .B(n13961), .Z(n14007) );
  NANDN U14110 ( .A(n13788), .B(n13787), .Z(n13792) );
  NANDN U14111 ( .A(n13790), .B(n13789), .Z(n13791) );
  AND U14112 ( .A(n13792), .B(n13791), .Z(n13946) );
  NANDN U14113 ( .A(n13794), .B(n13793), .Z(n13798) );
  NANDN U14114 ( .A(n13796), .B(n13795), .Z(n13797) );
  NAND U14115 ( .A(n13798), .B(n13797), .Z(n13947) );
  XNOR U14116 ( .A(n13946), .B(n13947), .Z(n13948) );
  NANDN U14117 ( .A(n13800), .B(n13799), .Z(n13804) );
  NAND U14118 ( .A(n13802), .B(n13801), .Z(n13803) );
  NAND U14119 ( .A(n13804), .B(n13803), .Z(n13949) );
  XNOR U14120 ( .A(n13948), .B(n13949), .Z(n14006) );
  XNOR U14121 ( .A(n14007), .B(n14006), .Z(n14009) );
  NAND U14122 ( .A(n13806), .B(n13805), .Z(n13810) );
  NAND U14123 ( .A(n13808), .B(n13807), .Z(n13809) );
  AND U14124 ( .A(n13810), .B(n13809), .Z(n14008) );
  XOR U14125 ( .A(n14009), .B(n14008), .Z(n14021) );
  NANDN U14126 ( .A(n13812), .B(n13811), .Z(n13816) );
  NANDN U14127 ( .A(n13814), .B(n13813), .Z(n13815) );
  AND U14128 ( .A(n13816), .B(n13815), .Z(n14018) );
  NANDN U14129 ( .A(n13822), .B(n13821), .Z(n13826) );
  OR U14130 ( .A(n13824), .B(n13823), .Z(n13825) );
  AND U14131 ( .A(n13826), .B(n13825), .Z(n14013) );
  NANDN U14132 ( .A(n13828), .B(n13827), .Z(n13832) );
  NANDN U14133 ( .A(n13830), .B(n13829), .Z(n13831) );
  AND U14134 ( .A(n13832), .B(n13831), .Z(n13953) );
  NANDN U14135 ( .A(n13834), .B(n13833), .Z(n13838) );
  OR U14136 ( .A(n13836), .B(n13835), .Z(n13837) );
  NAND U14137 ( .A(n13838), .B(n13837), .Z(n13952) );
  XNOR U14138 ( .A(n13953), .B(n13952), .Z(n13954) );
  NAND U14139 ( .A(b[0]), .B(a[108]), .Z(n13839) );
  XNOR U14140 ( .A(b[1]), .B(n13839), .Z(n13841) );
  NANDN U14141 ( .A(b[0]), .B(a[107]), .Z(n13840) );
  NAND U14142 ( .A(n13841), .B(n13840), .Z(n13901) );
  NANDN U14143 ( .A(n19394), .B(n13842), .Z(n13844) );
  XOR U14144 ( .A(b[29]), .B(a[80]), .Z(n13979) );
  NANDN U14145 ( .A(n19395), .B(n13979), .Z(n13843) );
  AND U14146 ( .A(n13844), .B(n13843), .Z(n13899) );
  AND U14147 ( .A(b[31]), .B(a[76]), .Z(n13898) );
  XNOR U14148 ( .A(n13899), .B(n13898), .Z(n13900) );
  XNOR U14149 ( .A(n13901), .B(n13900), .Z(n13940) );
  NANDN U14150 ( .A(n19005), .B(n13845), .Z(n13847) );
  XOR U14151 ( .A(b[23]), .B(a[86]), .Z(n13982) );
  NANDN U14152 ( .A(n19055), .B(n13982), .Z(n13846) );
  AND U14153 ( .A(n13847), .B(n13846), .Z(n13973) );
  NANDN U14154 ( .A(n17362), .B(n13848), .Z(n13850) );
  XOR U14155 ( .A(b[7]), .B(a[102]), .Z(n13985) );
  NANDN U14156 ( .A(n17522), .B(n13985), .Z(n13849) );
  AND U14157 ( .A(n13850), .B(n13849), .Z(n13971) );
  NANDN U14158 ( .A(n19116), .B(n13851), .Z(n13853) );
  XOR U14159 ( .A(b[25]), .B(a[84]), .Z(n13988) );
  NANDN U14160 ( .A(n19179), .B(n13988), .Z(n13852) );
  NAND U14161 ( .A(n13853), .B(n13852), .Z(n13970) );
  XNOR U14162 ( .A(n13971), .B(n13970), .Z(n13972) );
  XOR U14163 ( .A(n13973), .B(n13972), .Z(n13941) );
  XNOR U14164 ( .A(n13940), .B(n13941), .Z(n13942) );
  NANDN U14165 ( .A(n18113), .B(n13854), .Z(n13856) );
  XOR U14166 ( .A(b[13]), .B(a[96]), .Z(n13991) );
  NANDN U14167 ( .A(n18229), .B(n13991), .Z(n13855) );
  AND U14168 ( .A(n13856), .B(n13855), .Z(n13935) );
  NANDN U14169 ( .A(n17888), .B(n13857), .Z(n13859) );
  XOR U14170 ( .A(b[11]), .B(a[98]), .Z(n13994) );
  NANDN U14171 ( .A(n18025), .B(n13994), .Z(n13858) );
  NAND U14172 ( .A(n13859), .B(n13858), .Z(n13934) );
  XNOR U14173 ( .A(n13935), .B(n13934), .Z(n13936) );
  NANDN U14174 ( .A(n18487), .B(n13860), .Z(n13862) );
  XOR U14175 ( .A(b[15]), .B(a[94]), .Z(n13997) );
  NANDN U14176 ( .A(n18311), .B(n13997), .Z(n13861) );
  AND U14177 ( .A(n13862), .B(n13861), .Z(n13931) );
  NANDN U14178 ( .A(n18853), .B(n13863), .Z(n13865) );
  XOR U14179 ( .A(b[21]), .B(a[88]), .Z(n14000) );
  NANDN U14180 ( .A(n18926), .B(n14000), .Z(n13864) );
  AND U14181 ( .A(n13865), .B(n13864), .Z(n13929) );
  NANDN U14182 ( .A(n17613), .B(n13866), .Z(n13868) );
  XOR U14183 ( .A(b[9]), .B(a[100]), .Z(n14003) );
  NANDN U14184 ( .A(n17739), .B(n14003), .Z(n13867) );
  NAND U14185 ( .A(n13868), .B(n13867), .Z(n13928) );
  XNOR U14186 ( .A(n13929), .B(n13928), .Z(n13930) );
  XOR U14187 ( .A(n13931), .B(n13930), .Z(n13937) );
  XOR U14188 ( .A(n13936), .B(n13937), .Z(n13943) );
  XOR U14189 ( .A(n13942), .B(n13943), .Z(n13955) );
  XNOR U14190 ( .A(n13954), .B(n13955), .Z(n14012) );
  XNOR U14191 ( .A(n14013), .B(n14012), .Z(n14014) );
  XOR U14192 ( .A(n14015), .B(n14014), .Z(n14019) );
  XNOR U14193 ( .A(n14018), .B(n14019), .Z(n14020) );
  XNOR U14194 ( .A(n14021), .B(n14020), .Z(n14026) );
  XOR U14195 ( .A(n14027), .B(n14026), .Z(n13893) );
  NANDN U14196 ( .A(n13870), .B(n13869), .Z(n13874) );
  NANDN U14197 ( .A(n13872), .B(n13871), .Z(n13873) );
  AND U14198 ( .A(n13874), .B(n13873), .Z(n13892) );
  XNOR U14199 ( .A(n13893), .B(n13892), .Z(n13894) );
  NANDN U14200 ( .A(n13876), .B(n13875), .Z(n13880) );
  NAND U14201 ( .A(n13878), .B(n13877), .Z(n13879) );
  NAND U14202 ( .A(n13880), .B(n13879), .Z(n13895) );
  XNOR U14203 ( .A(n13894), .B(n13895), .Z(n13886) );
  XNOR U14204 ( .A(n13887), .B(n13886), .Z(n13888) );
  XNOR U14205 ( .A(n13889), .B(n13888), .Z(n14030) );
  XNOR U14206 ( .A(sreg[204]), .B(n14030), .Z(n14032) );
  NANDN U14207 ( .A(sreg[203]), .B(n13881), .Z(n13885) );
  NAND U14208 ( .A(n13883), .B(n13882), .Z(n13884) );
  NAND U14209 ( .A(n13885), .B(n13884), .Z(n14031) );
  XNOR U14210 ( .A(n14032), .B(n14031), .Z(c[204]) );
  NANDN U14211 ( .A(n13887), .B(n13886), .Z(n13891) );
  NANDN U14212 ( .A(n13889), .B(n13888), .Z(n13890) );
  AND U14213 ( .A(n13891), .B(n13890), .Z(n14038) );
  NANDN U14214 ( .A(n13893), .B(n13892), .Z(n13897) );
  NANDN U14215 ( .A(n13895), .B(n13894), .Z(n13896) );
  AND U14216 ( .A(n13897), .B(n13896), .Z(n14036) );
  NANDN U14217 ( .A(n13899), .B(n13898), .Z(n13903) );
  NANDN U14218 ( .A(n13901), .B(n13900), .Z(n13902) );
  AND U14219 ( .A(n13903), .B(n13902), .Z(n14125) );
  NANDN U14220 ( .A(n19237), .B(n13904), .Z(n13906) );
  XOR U14221 ( .A(b[27]), .B(a[83]), .Z(n14071) );
  NANDN U14222 ( .A(n19277), .B(n14071), .Z(n13905) );
  AND U14223 ( .A(n13906), .B(n13905), .Z(n14132) );
  NANDN U14224 ( .A(n17072), .B(n13907), .Z(n13909) );
  XOR U14225 ( .A(a[105]), .B(b[5]), .Z(n14074) );
  NANDN U14226 ( .A(n17223), .B(n14074), .Z(n13908) );
  AND U14227 ( .A(n13909), .B(n13908), .Z(n14130) );
  NANDN U14228 ( .A(n18673), .B(n13910), .Z(n13912) );
  XOR U14229 ( .A(b[19]), .B(a[91]), .Z(n14077) );
  NANDN U14230 ( .A(n18758), .B(n14077), .Z(n13911) );
  NAND U14231 ( .A(n13912), .B(n13911), .Z(n14129) );
  XNOR U14232 ( .A(n14130), .B(n14129), .Z(n14131) );
  XNOR U14233 ( .A(n14132), .B(n14131), .Z(n14123) );
  NANDN U14234 ( .A(n19425), .B(n13913), .Z(n13915) );
  XOR U14235 ( .A(b[31]), .B(a[79]), .Z(n14080) );
  NANDN U14236 ( .A(n19426), .B(n14080), .Z(n13914) );
  AND U14237 ( .A(n13915), .B(n13914), .Z(n14092) );
  NANDN U14238 ( .A(n17067), .B(n13916), .Z(n13918) );
  XOR U14239 ( .A(a[107]), .B(b[3]), .Z(n14083) );
  NANDN U14240 ( .A(n17068), .B(n14083), .Z(n13917) );
  AND U14241 ( .A(n13918), .B(n13917), .Z(n14090) );
  NANDN U14242 ( .A(n18514), .B(n13919), .Z(n13921) );
  XOR U14243 ( .A(b[17]), .B(a[93]), .Z(n14086) );
  NANDN U14244 ( .A(n18585), .B(n14086), .Z(n13920) );
  NAND U14245 ( .A(n13921), .B(n13920), .Z(n14089) );
  XNOR U14246 ( .A(n14090), .B(n14089), .Z(n14091) );
  XOR U14247 ( .A(n14092), .B(n14091), .Z(n14124) );
  XOR U14248 ( .A(n14123), .B(n14124), .Z(n14126) );
  XOR U14249 ( .A(n14125), .B(n14126), .Z(n14060) );
  NANDN U14250 ( .A(n13923), .B(n13922), .Z(n13927) );
  NANDN U14251 ( .A(n13925), .B(n13924), .Z(n13926) );
  AND U14252 ( .A(n13927), .B(n13926), .Z(n14113) );
  NANDN U14253 ( .A(n13929), .B(n13928), .Z(n13933) );
  NANDN U14254 ( .A(n13931), .B(n13930), .Z(n13932) );
  NAND U14255 ( .A(n13933), .B(n13932), .Z(n14114) );
  XNOR U14256 ( .A(n14113), .B(n14114), .Z(n14115) );
  NANDN U14257 ( .A(n13935), .B(n13934), .Z(n13939) );
  NANDN U14258 ( .A(n13937), .B(n13936), .Z(n13938) );
  NAND U14259 ( .A(n13939), .B(n13938), .Z(n14116) );
  XNOR U14260 ( .A(n14115), .B(n14116), .Z(n14059) );
  XNOR U14261 ( .A(n14060), .B(n14059), .Z(n14062) );
  NANDN U14262 ( .A(n13941), .B(n13940), .Z(n13945) );
  NANDN U14263 ( .A(n13943), .B(n13942), .Z(n13944) );
  AND U14264 ( .A(n13945), .B(n13944), .Z(n14061) );
  XOR U14265 ( .A(n14062), .B(n14061), .Z(n14173) );
  NANDN U14266 ( .A(n13947), .B(n13946), .Z(n13951) );
  NANDN U14267 ( .A(n13949), .B(n13948), .Z(n13950) );
  AND U14268 ( .A(n13951), .B(n13950), .Z(n14171) );
  NANDN U14269 ( .A(n13953), .B(n13952), .Z(n13957) );
  NANDN U14270 ( .A(n13955), .B(n13954), .Z(n13956) );
  AND U14271 ( .A(n13957), .B(n13956), .Z(n14056) );
  NANDN U14272 ( .A(n13959), .B(n13958), .Z(n13963) );
  OR U14273 ( .A(n13961), .B(n13960), .Z(n13962) );
  AND U14274 ( .A(n13963), .B(n13962), .Z(n14054) );
  NANDN U14275 ( .A(n13965), .B(n13964), .Z(n13969) );
  NANDN U14276 ( .A(n13967), .B(n13966), .Z(n13968) );
  AND U14277 ( .A(n13969), .B(n13968), .Z(n14120) );
  NANDN U14278 ( .A(n13971), .B(n13970), .Z(n13975) );
  NANDN U14279 ( .A(n13973), .B(n13972), .Z(n13974) );
  NAND U14280 ( .A(n13975), .B(n13974), .Z(n14119) );
  XNOR U14281 ( .A(n14120), .B(n14119), .Z(n14122) );
  NAND U14282 ( .A(b[0]), .B(a[109]), .Z(n13976) );
  XNOR U14283 ( .A(b[1]), .B(n13976), .Z(n13978) );
  NANDN U14284 ( .A(b[0]), .B(a[108]), .Z(n13977) );
  NAND U14285 ( .A(n13978), .B(n13977), .Z(n14068) );
  NANDN U14286 ( .A(n19394), .B(n13979), .Z(n13981) );
  XOR U14287 ( .A(b[29]), .B(a[81]), .Z(n14144) );
  NANDN U14288 ( .A(n19395), .B(n14144), .Z(n13980) );
  AND U14289 ( .A(n13981), .B(n13980), .Z(n14066) );
  AND U14290 ( .A(b[31]), .B(a[77]), .Z(n14065) );
  XNOR U14291 ( .A(n14066), .B(n14065), .Z(n14067) );
  XNOR U14292 ( .A(n14068), .B(n14067), .Z(n14108) );
  NANDN U14293 ( .A(n19005), .B(n13982), .Z(n13984) );
  XOR U14294 ( .A(b[23]), .B(a[87]), .Z(n14147) );
  NANDN U14295 ( .A(n19055), .B(n14147), .Z(n13983) );
  AND U14296 ( .A(n13984), .B(n13983), .Z(n14137) );
  NANDN U14297 ( .A(n17362), .B(n13985), .Z(n13987) );
  XOR U14298 ( .A(b[7]), .B(a[103]), .Z(n14150) );
  NANDN U14299 ( .A(n17522), .B(n14150), .Z(n13986) );
  AND U14300 ( .A(n13987), .B(n13986), .Z(n14136) );
  NANDN U14301 ( .A(n19116), .B(n13988), .Z(n13990) );
  XOR U14302 ( .A(b[25]), .B(a[85]), .Z(n14153) );
  NANDN U14303 ( .A(n19179), .B(n14153), .Z(n13989) );
  NAND U14304 ( .A(n13990), .B(n13989), .Z(n14135) );
  XOR U14305 ( .A(n14136), .B(n14135), .Z(n14138) );
  XOR U14306 ( .A(n14137), .B(n14138), .Z(n14107) );
  XOR U14307 ( .A(n14108), .B(n14107), .Z(n14110) );
  NANDN U14308 ( .A(n18113), .B(n13991), .Z(n13993) );
  XOR U14309 ( .A(b[13]), .B(a[97]), .Z(n14156) );
  NANDN U14310 ( .A(n18229), .B(n14156), .Z(n13992) );
  AND U14311 ( .A(n13993), .B(n13992), .Z(n14102) );
  NANDN U14312 ( .A(n17888), .B(n13994), .Z(n13996) );
  XOR U14313 ( .A(b[11]), .B(a[99]), .Z(n14159) );
  NANDN U14314 ( .A(n18025), .B(n14159), .Z(n13995) );
  NAND U14315 ( .A(n13996), .B(n13995), .Z(n14101) );
  XNOR U14316 ( .A(n14102), .B(n14101), .Z(n14104) );
  NANDN U14317 ( .A(n18487), .B(n13997), .Z(n13999) );
  XOR U14318 ( .A(b[15]), .B(a[95]), .Z(n14162) );
  NANDN U14319 ( .A(n18311), .B(n14162), .Z(n13998) );
  AND U14320 ( .A(n13999), .B(n13998), .Z(n14098) );
  NANDN U14321 ( .A(n18853), .B(n14000), .Z(n14002) );
  XOR U14322 ( .A(b[21]), .B(a[89]), .Z(n14165) );
  NANDN U14323 ( .A(n18926), .B(n14165), .Z(n14001) );
  AND U14324 ( .A(n14002), .B(n14001), .Z(n14096) );
  NANDN U14325 ( .A(n17613), .B(n14003), .Z(n14005) );
  XOR U14326 ( .A(b[9]), .B(a[101]), .Z(n14168) );
  NANDN U14327 ( .A(n17739), .B(n14168), .Z(n14004) );
  NAND U14328 ( .A(n14005), .B(n14004), .Z(n14095) );
  XNOR U14329 ( .A(n14096), .B(n14095), .Z(n14097) );
  XNOR U14330 ( .A(n14098), .B(n14097), .Z(n14103) );
  XOR U14331 ( .A(n14104), .B(n14103), .Z(n14109) );
  XOR U14332 ( .A(n14110), .B(n14109), .Z(n14121) );
  XOR U14333 ( .A(n14122), .B(n14121), .Z(n14053) );
  XNOR U14334 ( .A(n14054), .B(n14053), .Z(n14055) );
  XOR U14335 ( .A(n14056), .B(n14055), .Z(n14172) );
  XOR U14336 ( .A(n14171), .B(n14172), .Z(n14174) );
  XOR U14337 ( .A(n14173), .B(n14174), .Z(n14050) );
  NANDN U14338 ( .A(n14007), .B(n14006), .Z(n14011) );
  NAND U14339 ( .A(n14009), .B(n14008), .Z(n14010) );
  AND U14340 ( .A(n14011), .B(n14010), .Z(n14048) );
  NANDN U14341 ( .A(n14013), .B(n14012), .Z(n14017) );
  NANDN U14342 ( .A(n14015), .B(n14014), .Z(n14016) );
  AND U14343 ( .A(n14017), .B(n14016), .Z(n14047) );
  XNOR U14344 ( .A(n14048), .B(n14047), .Z(n14049) );
  XNOR U14345 ( .A(n14050), .B(n14049), .Z(n14041) );
  NANDN U14346 ( .A(n14019), .B(n14018), .Z(n14023) );
  NANDN U14347 ( .A(n14021), .B(n14020), .Z(n14022) );
  NAND U14348 ( .A(n14023), .B(n14022), .Z(n14042) );
  XNOR U14349 ( .A(n14041), .B(n14042), .Z(n14043) );
  NANDN U14350 ( .A(n14025), .B(n14024), .Z(n14029) );
  NAND U14351 ( .A(n14027), .B(n14026), .Z(n14028) );
  NAND U14352 ( .A(n14029), .B(n14028), .Z(n14044) );
  XNOR U14353 ( .A(n14043), .B(n14044), .Z(n14035) );
  XNOR U14354 ( .A(n14036), .B(n14035), .Z(n14037) );
  XNOR U14355 ( .A(n14038), .B(n14037), .Z(n14177) );
  XNOR U14356 ( .A(sreg[205]), .B(n14177), .Z(n14179) );
  NANDN U14357 ( .A(sreg[204]), .B(n14030), .Z(n14034) );
  NAND U14358 ( .A(n14032), .B(n14031), .Z(n14033) );
  NAND U14359 ( .A(n14034), .B(n14033), .Z(n14178) );
  XNOR U14360 ( .A(n14179), .B(n14178), .Z(c[205]) );
  NANDN U14361 ( .A(n14036), .B(n14035), .Z(n14040) );
  NANDN U14362 ( .A(n14038), .B(n14037), .Z(n14039) );
  AND U14363 ( .A(n14040), .B(n14039), .Z(n14185) );
  NANDN U14364 ( .A(n14042), .B(n14041), .Z(n14046) );
  NANDN U14365 ( .A(n14044), .B(n14043), .Z(n14045) );
  AND U14366 ( .A(n14046), .B(n14045), .Z(n14183) );
  NANDN U14367 ( .A(n14048), .B(n14047), .Z(n14052) );
  NANDN U14368 ( .A(n14050), .B(n14049), .Z(n14051) );
  AND U14369 ( .A(n14052), .B(n14051), .Z(n14191) );
  NANDN U14370 ( .A(n14054), .B(n14053), .Z(n14058) );
  NANDN U14371 ( .A(n14056), .B(n14055), .Z(n14057) );
  AND U14372 ( .A(n14058), .B(n14057), .Z(n14195) );
  NANDN U14373 ( .A(n14060), .B(n14059), .Z(n14064) );
  NAND U14374 ( .A(n14062), .B(n14061), .Z(n14063) );
  AND U14375 ( .A(n14064), .B(n14063), .Z(n14194) );
  XNOR U14376 ( .A(n14195), .B(n14194), .Z(n14197) );
  NANDN U14377 ( .A(n14066), .B(n14065), .Z(n14070) );
  NANDN U14378 ( .A(n14068), .B(n14067), .Z(n14069) );
  AND U14379 ( .A(n14070), .B(n14069), .Z(n14260) );
  NANDN U14380 ( .A(n19237), .B(n14071), .Z(n14073) );
  XOR U14381 ( .A(b[27]), .B(a[84]), .Z(n14206) );
  NANDN U14382 ( .A(n19277), .B(n14206), .Z(n14072) );
  AND U14383 ( .A(n14073), .B(n14072), .Z(n14267) );
  NANDN U14384 ( .A(n17072), .B(n14074), .Z(n14076) );
  XOR U14385 ( .A(a[106]), .B(b[5]), .Z(n14209) );
  NANDN U14386 ( .A(n17223), .B(n14209), .Z(n14075) );
  AND U14387 ( .A(n14076), .B(n14075), .Z(n14265) );
  NANDN U14388 ( .A(n18673), .B(n14077), .Z(n14079) );
  XOR U14389 ( .A(b[19]), .B(a[92]), .Z(n14212) );
  NANDN U14390 ( .A(n18758), .B(n14212), .Z(n14078) );
  NAND U14391 ( .A(n14079), .B(n14078), .Z(n14264) );
  XNOR U14392 ( .A(n14265), .B(n14264), .Z(n14266) );
  XNOR U14393 ( .A(n14267), .B(n14266), .Z(n14258) );
  NANDN U14394 ( .A(n19425), .B(n14080), .Z(n14082) );
  XOR U14395 ( .A(b[31]), .B(a[80]), .Z(n14215) );
  NANDN U14396 ( .A(n19426), .B(n14215), .Z(n14081) );
  AND U14397 ( .A(n14082), .B(n14081), .Z(n14227) );
  NANDN U14398 ( .A(n17067), .B(n14083), .Z(n14085) );
  XOR U14399 ( .A(a[108]), .B(b[3]), .Z(n14218) );
  NANDN U14400 ( .A(n17068), .B(n14218), .Z(n14084) );
  AND U14401 ( .A(n14085), .B(n14084), .Z(n14225) );
  NANDN U14402 ( .A(n18514), .B(n14086), .Z(n14088) );
  XOR U14403 ( .A(b[17]), .B(a[94]), .Z(n14221) );
  NANDN U14404 ( .A(n18585), .B(n14221), .Z(n14087) );
  NAND U14405 ( .A(n14088), .B(n14087), .Z(n14224) );
  XNOR U14406 ( .A(n14225), .B(n14224), .Z(n14226) );
  XOR U14407 ( .A(n14227), .B(n14226), .Z(n14259) );
  XOR U14408 ( .A(n14258), .B(n14259), .Z(n14261) );
  XOR U14409 ( .A(n14260), .B(n14261), .Z(n14307) );
  NANDN U14410 ( .A(n14090), .B(n14089), .Z(n14094) );
  NANDN U14411 ( .A(n14092), .B(n14091), .Z(n14093) );
  AND U14412 ( .A(n14094), .B(n14093), .Z(n14248) );
  NANDN U14413 ( .A(n14096), .B(n14095), .Z(n14100) );
  NANDN U14414 ( .A(n14098), .B(n14097), .Z(n14099) );
  NAND U14415 ( .A(n14100), .B(n14099), .Z(n14249) );
  XNOR U14416 ( .A(n14248), .B(n14249), .Z(n14250) );
  NANDN U14417 ( .A(n14102), .B(n14101), .Z(n14106) );
  NAND U14418 ( .A(n14104), .B(n14103), .Z(n14105) );
  NAND U14419 ( .A(n14106), .B(n14105), .Z(n14251) );
  XNOR U14420 ( .A(n14250), .B(n14251), .Z(n14306) );
  XNOR U14421 ( .A(n14307), .B(n14306), .Z(n14309) );
  NAND U14422 ( .A(n14108), .B(n14107), .Z(n14112) );
  NAND U14423 ( .A(n14110), .B(n14109), .Z(n14111) );
  AND U14424 ( .A(n14112), .B(n14111), .Z(n14308) );
  XOR U14425 ( .A(n14309), .B(n14308), .Z(n14321) );
  NANDN U14426 ( .A(n14114), .B(n14113), .Z(n14118) );
  NANDN U14427 ( .A(n14116), .B(n14115), .Z(n14117) );
  AND U14428 ( .A(n14118), .B(n14117), .Z(n14318) );
  NANDN U14429 ( .A(n14124), .B(n14123), .Z(n14128) );
  OR U14430 ( .A(n14126), .B(n14125), .Z(n14127) );
  AND U14431 ( .A(n14128), .B(n14127), .Z(n14313) );
  NANDN U14432 ( .A(n14130), .B(n14129), .Z(n14134) );
  NANDN U14433 ( .A(n14132), .B(n14131), .Z(n14133) );
  AND U14434 ( .A(n14134), .B(n14133), .Z(n14255) );
  NANDN U14435 ( .A(n14136), .B(n14135), .Z(n14140) );
  OR U14436 ( .A(n14138), .B(n14137), .Z(n14139) );
  NAND U14437 ( .A(n14140), .B(n14139), .Z(n14254) );
  XNOR U14438 ( .A(n14255), .B(n14254), .Z(n14257) );
  AND U14439 ( .A(a[110]), .B(b[0]), .Z(n14141) );
  XOR U14440 ( .A(b[1]), .B(n14141), .Z(n14143) );
  NANDN U14441 ( .A(b[0]), .B(a[109]), .Z(n14142) );
  AND U14442 ( .A(n14143), .B(n14142), .Z(n14202) );
  NANDN U14443 ( .A(n19394), .B(n14144), .Z(n14146) );
  XOR U14444 ( .A(b[29]), .B(a[82]), .Z(n14279) );
  NANDN U14445 ( .A(n19395), .B(n14279), .Z(n14145) );
  AND U14446 ( .A(n14146), .B(n14145), .Z(n14201) );
  AND U14447 ( .A(b[31]), .B(a[78]), .Z(n14200) );
  XOR U14448 ( .A(n14201), .B(n14200), .Z(n14203) );
  XNOR U14449 ( .A(n14202), .B(n14203), .Z(n14243) );
  NANDN U14450 ( .A(n19005), .B(n14147), .Z(n14149) );
  XOR U14451 ( .A(b[23]), .B(a[88]), .Z(n14282) );
  NANDN U14452 ( .A(n19055), .B(n14282), .Z(n14148) );
  AND U14453 ( .A(n14149), .B(n14148), .Z(n14272) );
  NANDN U14454 ( .A(n17362), .B(n14150), .Z(n14152) );
  XOR U14455 ( .A(a[104]), .B(b[7]), .Z(n14285) );
  NANDN U14456 ( .A(n17522), .B(n14285), .Z(n14151) );
  AND U14457 ( .A(n14152), .B(n14151), .Z(n14271) );
  NANDN U14458 ( .A(n19116), .B(n14153), .Z(n14155) );
  XOR U14459 ( .A(b[25]), .B(a[86]), .Z(n14288) );
  NANDN U14460 ( .A(n19179), .B(n14288), .Z(n14154) );
  NAND U14461 ( .A(n14155), .B(n14154), .Z(n14270) );
  XOR U14462 ( .A(n14271), .B(n14270), .Z(n14273) );
  XOR U14463 ( .A(n14272), .B(n14273), .Z(n14242) );
  XOR U14464 ( .A(n14243), .B(n14242), .Z(n14245) );
  NANDN U14465 ( .A(n18113), .B(n14156), .Z(n14158) );
  XOR U14466 ( .A(b[13]), .B(a[98]), .Z(n14291) );
  NANDN U14467 ( .A(n18229), .B(n14291), .Z(n14157) );
  AND U14468 ( .A(n14158), .B(n14157), .Z(n14237) );
  NANDN U14469 ( .A(n17888), .B(n14159), .Z(n14161) );
  XOR U14470 ( .A(b[11]), .B(a[100]), .Z(n14294) );
  NANDN U14471 ( .A(n18025), .B(n14294), .Z(n14160) );
  NAND U14472 ( .A(n14161), .B(n14160), .Z(n14236) );
  XNOR U14473 ( .A(n14237), .B(n14236), .Z(n14239) );
  NANDN U14474 ( .A(n18487), .B(n14162), .Z(n14164) );
  XOR U14475 ( .A(b[15]), .B(a[96]), .Z(n14297) );
  NANDN U14476 ( .A(n18311), .B(n14297), .Z(n14163) );
  AND U14477 ( .A(n14164), .B(n14163), .Z(n14233) );
  NANDN U14478 ( .A(n18853), .B(n14165), .Z(n14167) );
  XOR U14479 ( .A(b[21]), .B(a[90]), .Z(n14300) );
  NANDN U14480 ( .A(n18926), .B(n14300), .Z(n14166) );
  AND U14481 ( .A(n14167), .B(n14166), .Z(n14231) );
  NANDN U14482 ( .A(n17613), .B(n14168), .Z(n14170) );
  XOR U14483 ( .A(b[9]), .B(a[102]), .Z(n14303) );
  NANDN U14484 ( .A(n17739), .B(n14303), .Z(n14169) );
  NAND U14485 ( .A(n14170), .B(n14169), .Z(n14230) );
  XNOR U14486 ( .A(n14231), .B(n14230), .Z(n14232) );
  XNOR U14487 ( .A(n14233), .B(n14232), .Z(n14238) );
  XOR U14488 ( .A(n14239), .B(n14238), .Z(n14244) );
  XOR U14489 ( .A(n14245), .B(n14244), .Z(n14256) );
  XOR U14490 ( .A(n14257), .B(n14256), .Z(n14312) );
  XNOR U14491 ( .A(n14313), .B(n14312), .Z(n14314) );
  XOR U14492 ( .A(n14315), .B(n14314), .Z(n14319) );
  XNOR U14493 ( .A(n14318), .B(n14319), .Z(n14320) );
  XNOR U14494 ( .A(n14321), .B(n14320), .Z(n14196) );
  XOR U14495 ( .A(n14197), .B(n14196), .Z(n14189) );
  NANDN U14496 ( .A(n14172), .B(n14171), .Z(n14176) );
  OR U14497 ( .A(n14174), .B(n14173), .Z(n14175) );
  AND U14498 ( .A(n14176), .B(n14175), .Z(n14188) );
  XNOR U14499 ( .A(n14189), .B(n14188), .Z(n14190) );
  XNOR U14500 ( .A(n14191), .B(n14190), .Z(n14182) );
  XNOR U14501 ( .A(n14183), .B(n14182), .Z(n14184) );
  XNOR U14502 ( .A(n14185), .B(n14184), .Z(n14324) );
  XNOR U14503 ( .A(sreg[206]), .B(n14324), .Z(n14326) );
  NANDN U14504 ( .A(sreg[205]), .B(n14177), .Z(n14181) );
  NAND U14505 ( .A(n14179), .B(n14178), .Z(n14180) );
  NAND U14506 ( .A(n14181), .B(n14180), .Z(n14325) );
  XNOR U14507 ( .A(n14326), .B(n14325), .Z(c[206]) );
  NANDN U14508 ( .A(n14183), .B(n14182), .Z(n14187) );
  NANDN U14509 ( .A(n14185), .B(n14184), .Z(n14186) );
  AND U14510 ( .A(n14187), .B(n14186), .Z(n14332) );
  NANDN U14511 ( .A(n14189), .B(n14188), .Z(n14193) );
  NANDN U14512 ( .A(n14191), .B(n14190), .Z(n14192) );
  AND U14513 ( .A(n14193), .B(n14192), .Z(n14330) );
  NANDN U14514 ( .A(n14195), .B(n14194), .Z(n14199) );
  NAND U14515 ( .A(n14197), .B(n14196), .Z(n14198) );
  AND U14516 ( .A(n14199), .B(n14198), .Z(n14337) );
  NANDN U14517 ( .A(n14201), .B(n14200), .Z(n14205) );
  NANDN U14518 ( .A(n14203), .B(n14202), .Z(n14204) );
  AND U14519 ( .A(n14205), .B(n14204), .Z(n14409) );
  NANDN U14520 ( .A(n19237), .B(n14206), .Z(n14208) );
  XOR U14521 ( .A(b[27]), .B(a[85]), .Z(n14353) );
  NANDN U14522 ( .A(n19277), .B(n14353), .Z(n14207) );
  AND U14523 ( .A(n14208), .B(n14207), .Z(n14416) );
  NANDN U14524 ( .A(n17072), .B(n14209), .Z(n14211) );
  XOR U14525 ( .A(a[107]), .B(b[5]), .Z(n14356) );
  NANDN U14526 ( .A(n17223), .B(n14356), .Z(n14210) );
  AND U14527 ( .A(n14211), .B(n14210), .Z(n14414) );
  NANDN U14528 ( .A(n18673), .B(n14212), .Z(n14214) );
  XOR U14529 ( .A(b[19]), .B(a[93]), .Z(n14359) );
  NANDN U14530 ( .A(n18758), .B(n14359), .Z(n14213) );
  NAND U14531 ( .A(n14214), .B(n14213), .Z(n14413) );
  XNOR U14532 ( .A(n14414), .B(n14413), .Z(n14415) );
  XNOR U14533 ( .A(n14416), .B(n14415), .Z(n14407) );
  NANDN U14534 ( .A(n19425), .B(n14215), .Z(n14217) );
  XOR U14535 ( .A(b[31]), .B(a[81]), .Z(n14362) );
  NANDN U14536 ( .A(n19426), .B(n14362), .Z(n14216) );
  AND U14537 ( .A(n14217), .B(n14216), .Z(n14374) );
  NANDN U14538 ( .A(n17067), .B(n14218), .Z(n14220) );
  XOR U14539 ( .A(a[109]), .B(b[3]), .Z(n14365) );
  NANDN U14540 ( .A(n17068), .B(n14365), .Z(n14219) );
  AND U14541 ( .A(n14220), .B(n14219), .Z(n14372) );
  NANDN U14542 ( .A(n18514), .B(n14221), .Z(n14223) );
  XOR U14543 ( .A(b[17]), .B(a[95]), .Z(n14368) );
  NANDN U14544 ( .A(n18585), .B(n14368), .Z(n14222) );
  NAND U14545 ( .A(n14223), .B(n14222), .Z(n14371) );
  XNOR U14546 ( .A(n14372), .B(n14371), .Z(n14373) );
  XOR U14547 ( .A(n14374), .B(n14373), .Z(n14408) );
  XOR U14548 ( .A(n14407), .B(n14408), .Z(n14410) );
  XOR U14549 ( .A(n14409), .B(n14410), .Z(n14456) );
  NANDN U14550 ( .A(n14225), .B(n14224), .Z(n14229) );
  NANDN U14551 ( .A(n14227), .B(n14226), .Z(n14228) );
  AND U14552 ( .A(n14229), .B(n14228), .Z(n14395) );
  NANDN U14553 ( .A(n14231), .B(n14230), .Z(n14235) );
  NANDN U14554 ( .A(n14233), .B(n14232), .Z(n14234) );
  NAND U14555 ( .A(n14235), .B(n14234), .Z(n14396) );
  XNOR U14556 ( .A(n14395), .B(n14396), .Z(n14397) );
  NANDN U14557 ( .A(n14237), .B(n14236), .Z(n14241) );
  NAND U14558 ( .A(n14239), .B(n14238), .Z(n14240) );
  NAND U14559 ( .A(n14241), .B(n14240), .Z(n14398) );
  XNOR U14560 ( .A(n14397), .B(n14398), .Z(n14455) );
  XNOR U14561 ( .A(n14456), .B(n14455), .Z(n14458) );
  NAND U14562 ( .A(n14243), .B(n14242), .Z(n14247) );
  NAND U14563 ( .A(n14245), .B(n14244), .Z(n14246) );
  AND U14564 ( .A(n14247), .B(n14246), .Z(n14457) );
  XOR U14565 ( .A(n14458), .B(n14457), .Z(n14469) );
  NANDN U14566 ( .A(n14249), .B(n14248), .Z(n14253) );
  NANDN U14567 ( .A(n14251), .B(n14250), .Z(n14252) );
  AND U14568 ( .A(n14253), .B(n14252), .Z(n14467) );
  NANDN U14569 ( .A(n14259), .B(n14258), .Z(n14263) );
  OR U14570 ( .A(n14261), .B(n14260), .Z(n14262) );
  AND U14571 ( .A(n14263), .B(n14262), .Z(n14462) );
  NANDN U14572 ( .A(n14265), .B(n14264), .Z(n14269) );
  NANDN U14573 ( .A(n14267), .B(n14266), .Z(n14268) );
  AND U14574 ( .A(n14269), .B(n14268), .Z(n14402) );
  NANDN U14575 ( .A(n14271), .B(n14270), .Z(n14275) );
  OR U14576 ( .A(n14273), .B(n14272), .Z(n14274) );
  NAND U14577 ( .A(n14275), .B(n14274), .Z(n14401) );
  XNOR U14578 ( .A(n14402), .B(n14401), .Z(n14403) );
  NAND U14579 ( .A(b[0]), .B(a[111]), .Z(n14276) );
  XNOR U14580 ( .A(b[1]), .B(n14276), .Z(n14278) );
  NANDN U14581 ( .A(b[0]), .B(a[110]), .Z(n14277) );
  NAND U14582 ( .A(n14278), .B(n14277), .Z(n14350) );
  NANDN U14583 ( .A(n19394), .B(n14279), .Z(n14281) );
  XOR U14584 ( .A(b[29]), .B(a[83]), .Z(n14428) );
  NANDN U14585 ( .A(n19395), .B(n14428), .Z(n14280) );
  AND U14586 ( .A(n14281), .B(n14280), .Z(n14348) );
  AND U14587 ( .A(b[31]), .B(a[79]), .Z(n14347) );
  XNOR U14588 ( .A(n14348), .B(n14347), .Z(n14349) );
  XNOR U14589 ( .A(n14350), .B(n14349), .Z(n14389) );
  NANDN U14590 ( .A(n19005), .B(n14282), .Z(n14284) );
  XOR U14591 ( .A(b[23]), .B(a[89]), .Z(n14431) );
  NANDN U14592 ( .A(n19055), .B(n14431), .Z(n14283) );
  AND U14593 ( .A(n14284), .B(n14283), .Z(n14422) );
  NANDN U14594 ( .A(n17362), .B(n14285), .Z(n14287) );
  XOR U14595 ( .A(b[7]), .B(a[105]), .Z(n14434) );
  NANDN U14596 ( .A(n17522), .B(n14434), .Z(n14286) );
  AND U14597 ( .A(n14287), .B(n14286), .Z(n14420) );
  NANDN U14598 ( .A(n19116), .B(n14288), .Z(n14290) );
  XOR U14599 ( .A(b[25]), .B(a[87]), .Z(n14437) );
  NANDN U14600 ( .A(n19179), .B(n14437), .Z(n14289) );
  NAND U14601 ( .A(n14290), .B(n14289), .Z(n14419) );
  XNOR U14602 ( .A(n14420), .B(n14419), .Z(n14421) );
  XOR U14603 ( .A(n14422), .B(n14421), .Z(n14390) );
  XNOR U14604 ( .A(n14389), .B(n14390), .Z(n14391) );
  NANDN U14605 ( .A(n18113), .B(n14291), .Z(n14293) );
  XOR U14606 ( .A(b[13]), .B(a[99]), .Z(n14440) );
  NANDN U14607 ( .A(n18229), .B(n14440), .Z(n14292) );
  AND U14608 ( .A(n14293), .B(n14292), .Z(n14384) );
  NANDN U14609 ( .A(n17888), .B(n14294), .Z(n14296) );
  XOR U14610 ( .A(b[11]), .B(a[101]), .Z(n14443) );
  NANDN U14611 ( .A(n18025), .B(n14443), .Z(n14295) );
  NAND U14612 ( .A(n14296), .B(n14295), .Z(n14383) );
  XNOR U14613 ( .A(n14384), .B(n14383), .Z(n14385) );
  NANDN U14614 ( .A(n18487), .B(n14297), .Z(n14299) );
  XOR U14615 ( .A(b[15]), .B(a[97]), .Z(n14446) );
  NANDN U14616 ( .A(n18311), .B(n14446), .Z(n14298) );
  AND U14617 ( .A(n14299), .B(n14298), .Z(n14380) );
  NANDN U14618 ( .A(n18853), .B(n14300), .Z(n14302) );
  XOR U14619 ( .A(b[21]), .B(a[91]), .Z(n14449) );
  NANDN U14620 ( .A(n18926), .B(n14449), .Z(n14301) );
  AND U14621 ( .A(n14302), .B(n14301), .Z(n14378) );
  NANDN U14622 ( .A(n17613), .B(n14303), .Z(n14305) );
  XOR U14623 ( .A(b[9]), .B(a[103]), .Z(n14452) );
  NANDN U14624 ( .A(n17739), .B(n14452), .Z(n14304) );
  NAND U14625 ( .A(n14305), .B(n14304), .Z(n14377) );
  XNOR U14626 ( .A(n14378), .B(n14377), .Z(n14379) );
  XOR U14627 ( .A(n14380), .B(n14379), .Z(n14386) );
  XOR U14628 ( .A(n14385), .B(n14386), .Z(n14392) );
  XOR U14629 ( .A(n14391), .B(n14392), .Z(n14404) );
  XNOR U14630 ( .A(n14403), .B(n14404), .Z(n14461) );
  XNOR U14631 ( .A(n14462), .B(n14461), .Z(n14463) );
  XOR U14632 ( .A(n14464), .B(n14463), .Z(n14468) );
  XOR U14633 ( .A(n14467), .B(n14468), .Z(n14470) );
  XOR U14634 ( .A(n14469), .B(n14470), .Z(n14344) );
  NANDN U14635 ( .A(n14307), .B(n14306), .Z(n14311) );
  NAND U14636 ( .A(n14309), .B(n14308), .Z(n14310) );
  AND U14637 ( .A(n14311), .B(n14310), .Z(n14342) );
  NANDN U14638 ( .A(n14313), .B(n14312), .Z(n14317) );
  NANDN U14639 ( .A(n14315), .B(n14314), .Z(n14316) );
  AND U14640 ( .A(n14317), .B(n14316), .Z(n14341) );
  XNOR U14641 ( .A(n14342), .B(n14341), .Z(n14343) );
  XNOR U14642 ( .A(n14344), .B(n14343), .Z(n14335) );
  NANDN U14643 ( .A(n14319), .B(n14318), .Z(n14323) );
  NANDN U14644 ( .A(n14321), .B(n14320), .Z(n14322) );
  NAND U14645 ( .A(n14323), .B(n14322), .Z(n14336) );
  XOR U14646 ( .A(n14335), .B(n14336), .Z(n14338) );
  XNOR U14647 ( .A(n14337), .B(n14338), .Z(n14329) );
  XNOR U14648 ( .A(n14330), .B(n14329), .Z(n14331) );
  XNOR U14649 ( .A(n14332), .B(n14331), .Z(n14473) );
  XNOR U14650 ( .A(sreg[207]), .B(n14473), .Z(n14475) );
  NANDN U14651 ( .A(sreg[206]), .B(n14324), .Z(n14328) );
  NAND U14652 ( .A(n14326), .B(n14325), .Z(n14327) );
  NAND U14653 ( .A(n14328), .B(n14327), .Z(n14474) );
  XNOR U14654 ( .A(n14475), .B(n14474), .Z(c[207]) );
  NANDN U14655 ( .A(n14330), .B(n14329), .Z(n14334) );
  NANDN U14656 ( .A(n14332), .B(n14331), .Z(n14333) );
  AND U14657 ( .A(n14334), .B(n14333), .Z(n14481) );
  NANDN U14658 ( .A(n14336), .B(n14335), .Z(n14340) );
  NANDN U14659 ( .A(n14338), .B(n14337), .Z(n14339) );
  AND U14660 ( .A(n14340), .B(n14339), .Z(n14479) );
  NANDN U14661 ( .A(n14342), .B(n14341), .Z(n14346) );
  NANDN U14662 ( .A(n14344), .B(n14343), .Z(n14345) );
  AND U14663 ( .A(n14346), .B(n14345), .Z(n14487) );
  NANDN U14664 ( .A(n14348), .B(n14347), .Z(n14352) );
  NANDN U14665 ( .A(n14350), .B(n14349), .Z(n14351) );
  AND U14666 ( .A(n14352), .B(n14351), .Z(n14570) );
  NANDN U14667 ( .A(n19237), .B(n14353), .Z(n14355) );
  XOR U14668 ( .A(b[27]), .B(a[86]), .Z(n14514) );
  NANDN U14669 ( .A(n19277), .B(n14514), .Z(n14354) );
  AND U14670 ( .A(n14355), .B(n14354), .Z(n14577) );
  NANDN U14671 ( .A(n17072), .B(n14356), .Z(n14358) );
  XOR U14672 ( .A(a[108]), .B(b[5]), .Z(n14517) );
  NANDN U14673 ( .A(n17223), .B(n14517), .Z(n14357) );
  AND U14674 ( .A(n14358), .B(n14357), .Z(n14575) );
  NANDN U14675 ( .A(n18673), .B(n14359), .Z(n14361) );
  XOR U14676 ( .A(b[19]), .B(a[94]), .Z(n14520) );
  NANDN U14677 ( .A(n18758), .B(n14520), .Z(n14360) );
  NAND U14678 ( .A(n14361), .B(n14360), .Z(n14574) );
  XNOR U14679 ( .A(n14575), .B(n14574), .Z(n14576) );
  XNOR U14680 ( .A(n14577), .B(n14576), .Z(n14568) );
  NANDN U14681 ( .A(n19425), .B(n14362), .Z(n14364) );
  XOR U14682 ( .A(b[31]), .B(a[82]), .Z(n14523) );
  NANDN U14683 ( .A(n19426), .B(n14523), .Z(n14363) );
  AND U14684 ( .A(n14364), .B(n14363), .Z(n14535) );
  NANDN U14685 ( .A(n17067), .B(n14365), .Z(n14367) );
  XOR U14686 ( .A(a[110]), .B(b[3]), .Z(n14526) );
  NANDN U14687 ( .A(n17068), .B(n14526), .Z(n14366) );
  AND U14688 ( .A(n14367), .B(n14366), .Z(n14533) );
  NANDN U14689 ( .A(n18514), .B(n14368), .Z(n14370) );
  XOR U14690 ( .A(b[17]), .B(a[96]), .Z(n14529) );
  NANDN U14691 ( .A(n18585), .B(n14529), .Z(n14369) );
  NAND U14692 ( .A(n14370), .B(n14369), .Z(n14532) );
  XNOR U14693 ( .A(n14533), .B(n14532), .Z(n14534) );
  XOR U14694 ( .A(n14535), .B(n14534), .Z(n14569) );
  XOR U14695 ( .A(n14568), .B(n14569), .Z(n14571) );
  XOR U14696 ( .A(n14570), .B(n14571), .Z(n14503) );
  NANDN U14697 ( .A(n14372), .B(n14371), .Z(n14376) );
  NANDN U14698 ( .A(n14374), .B(n14373), .Z(n14375) );
  AND U14699 ( .A(n14376), .B(n14375), .Z(n14556) );
  NANDN U14700 ( .A(n14378), .B(n14377), .Z(n14382) );
  NANDN U14701 ( .A(n14380), .B(n14379), .Z(n14381) );
  NAND U14702 ( .A(n14382), .B(n14381), .Z(n14557) );
  XNOR U14703 ( .A(n14556), .B(n14557), .Z(n14558) );
  NANDN U14704 ( .A(n14384), .B(n14383), .Z(n14388) );
  NANDN U14705 ( .A(n14386), .B(n14385), .Z(n14387) );
  NAND U14706 ( .A(n14388), .B(n14387), .Z(n14559) );
  XNOR U14707 ( .A(n14558), .B(n14559), .Z(n14502) );
  XNOR U14708 ( .A(n14503), .B(n14502), .Z(n14505) );
  NANDN U14709 ( .A(n14390), .B(n14389), .Z(n14394) );
  NANDN U14710 ( .A(n14392), .B(n14391), .Z(n14393) );
  AND U14711 ( .A(n14394), .B(n14393), .Z(n14504) );
  XOR U14712 ( .A(n14505), .B(n14504), .Z(n14618) );
  NANDN U14713 ( .A(n14396), .B(n14395), .Z(n14400) );
  NANDN U14714 ( .A(n14398), .B(n14397), .Z(n14399) );
  AND U14715 ( .A(n14400), .B(n14399), .Z(n14616) );
  NANDN U14716 ( .A(n14402), .B(n14401), .Z(n14406) );
  NANDN U14717 ( .A(n14404), .B(n14403), .Z(n14405) );
  AND U14718 ( .A(n14406), .B(n14405), .Z(n14499) );
  NANDN U14719 ( .A(n14408), .B(n14407), .Z(n14412) );
  OR U14720 ( .A(n14410), .B(n14409), .Z(n14411) );
  AND U14721 ( .A(n14412), .B(n14411), .Z(n14497) );
  NANDN U14722 ( .A(n14414), .B(n14413), .Z(n14418) );
  NANDN U14723 ( .A(n14416), .B(n14415), .Z(n14417) );
  AND U14724 ( .A(n14418), .B(n14417), .Z(n14563) );
  NANDN U14725 ( .A(n14420), .B(n14419), .Z(n14424) );
  NANDN U14726 ( .A(n14422), .B(n14421), .Z(n14423) );
  NAND U14727 ( .A(n14424), .B(n14423), .Z(n14562) );
  XNOR U14728 ( .A(n14563), .B(n14562), .Z(n14564) );
  NAND U14729 ( .A(b[0]), .B(a[112]), .Z(n14425) );
  XNOR U14730 ( .A(b[1]), .B(n14425), .Z(n14427) );
  NANDN U14731 ( .A(b[0]), .B(a[111]), .Z(n14426) );
  NAND U14732 ( .A(n14427), .B(n14426), .Z(n14511) );
  NANDN U14733 ( .A(n19394), .B(n14428), .Z(n14430) );
  XOR U14734 ( .A(b[29]), .B(a[84]), .Z(n14589) );
  NANDN U14735 ( .A(n19395), .B(n14589), .Z(n14429) );
  AND U14736 ( .A(n14430), .B(n14429), .Z(n14509) );
  AND U14737 ( .A(b[31]), .B(a[80]), .Z(n14508) );
  XNOR U14738 ( .A(n14509), .B(n14508), .Z(n14510) );
  XNOR U14739 ( .A(n14511), .B(n14510), .Z(n14550) );
  NANDN U14740 ( .A(n19005), .B(n14431), .Z(n14433) );
  XOR U14741 ( .A(b[23]), .B(a[90]), .Z(n14592) );
  NANDN U14742 ( .A(n19055), .B(n14592), .Z(n14432) );
  AND U14743 ( .A(n14433), .B(n14432), .Z(n14583) );
  NANDN U14744 ( .A(n17362), .B(n14434), .Z(n14436) );
  XOR U14745 ( .A(a[106]), .B(b[7]), .Z(n14595) );
  NANDN U14746 ( .A(n17522), .B(n14595), .Z(n14435) );
  AND U14747 ( .A(n14436), .B(n14435), .Z(n14581) );
  NANDN U14748 ( .A(n19116), .B(n14437), .Z(n14439) );
  XOR U14749 ( .A(b[25]), .B(a[88]), .Z(n14598) );
  NANDN U14750 ( .A(n19179), .B(n14598), .Z(n14438) );
  NAND U14751 ( .A(n14439), .B(n14438), .Z(n14580) );
  XNOR U14752 ( .A(n14581), .B(n14580), .Z(n14582) );
  XOR U14753 ( .A(n14583), .B(n14582), .Z(n14551) );
  XNOR U14754 ( .A(n14550), .B(n14551), .Z(n14552) );
  NANDN U14755 ( .A(n18113), .B(n14440), .Z(n14442) );
  XOR U14756 ( .A(b[13]), .B(a[100]), .Z(n14601) );
  NANDN U14757 ( .A(n18229), .B(n14601), .Z(n14441) );
  AND U14758 ( .A(n14442), .B(n14441), .Z(n14545) );
  NANDN U14759 ( .A(n17888), .B(n14443), .Z(n14445) );
  XOR U14760 ( .A(b[11]), .B(a[102]), .Z(n14604) );
  NANDN U14761 ( .A(n18025), .B(n14604), .Z(n14444) );
  NAND U14762 ( .A(n14445), .B(n14444), .Z(n14544) );
  XNOR U14763 ( .A(n14545), .B(n14544), .Z(n14546) );
  NANDN U14764 ( .A(n18487), .B(n14446), .Z(n14448) );
  XOR U14765 ( .A(b[15]), .B(a[98]), .Z(n14607) );
  NANDN U14766 ( .A(n18311), .B(n14607), .Z(n14447) );
  AND U14767 ( .A(n14448), .B(n14447), .Z(n14541) );
  NANDN U14768 ( .A(n18853), .B(n14449), .Z(n14451) );
  XOR U14769 ( .A(b[21]), .B(a[92]), .Z(n14610) );
  NANDN U14770 ( .A(n18926), .B(n14610), .Z(n14450) );
  AND U14771 ( .A(n14451), .B(n14450), .Z(n14539) );
  NANDN U14772 ( .A(n17613), .B(n14452), .Z(n14454) );
  XOR U14773 ( .A(b[9]), .B(a[104]), .Z(n14613) );
  NANDN U14774 ( .A(n17739), .B(n14613), .Z(n14453) );
  NAND U14775 ( .A(n14454), .B(n14453), .Z(n14538) );
  XNOR U14776 ( .A(n14539), .B(n14538), .Z(n14540) );
  XOR U14777 ( .A(n14541), .B(n14540), .Z(n14547) );
  XOR U14778 ( .A(n14546), .B(n14547), .Z(n14553) );
  XOR U14779 ( .A(n14552), .B(n14553), .Z(n14565) );
  XNOR U14780 ( .A(n14564), .B(n14565), .Z(n14496) );
  XNOR U14781 ( .A(n14497), .B(n14496), .Z(n14498) );
  XOR U14782 ( .A(n14499), .B(n14498), .Z(n14617) );
  XOR U14783 ( .A(n14616), .B(n14617), .Z(n14619) );
  XOR U14784 ( .A(n14618), .B(n14619), .Z(n14493) );
  NANDN U14785 ( .A(n14456), .B(n14455), .Z(n14460) );
  NAND U14786 ( .A(n14458), .B(n14457), .Z(n14459) );
  AND U14787 ( .A(n14460), .B(n14459), .Z(n14491) );
  NANDN U14788 ( .A(n14462), .B(n14461), .Z(n14466) );
  NANDN U14789 ( .A(n14464), .B(n14463), .Z(n14465) );
  AND U14790 ( .A(n14466), .B(n14465), .Z(n14490) );
  XNOR U14791 ( .A(n14491), .B(n14490), .Z(n14492) );
  XNOR U14792 ( .A(n14493), .B(n14492), .Z(n14484) );
  NANDN U14793 ( .A(n14468), .B(n14467), .Z(n14472) );
  OR U14794 ( .A(n14470), .B(n14469), .Z(n14471) );
  NAND U14795 ( .A(n14472), .B(n14471), .Z(n14485) );
  XNOR U14796 ( .A(n14484), .B(n14485), .Z(n14486) );
  XNOR U14797 ( .A(n14487), .B(n14486), .Z(n14478) );
  XNOR U14798 ( .A(n14479), .B(n14478), .Z(n14480) );
  XNOR U14799 ( .A(n14481), .B(n14480), .Z(n14622) );
  XNOR U14800 ( .A(sreg[208]), .B(n14622), .Z(n14624) );
  NANDN U14801 ( .A(sreg[207]), .B(n14473), .Z(n14477) );
  NAND U14802 ( .A(n14475), .B(n14474), .Z(n14476) );
  NAND U14803 ( .A(n14477), .B(n14476), .Z(n14623) );
  XNOR U14804 ( .A(n14624), .B(n14623), .Z(c[208]) );
  NANDN U14805 ( .A(n14479), .B(n14478), .Z(n14483) );
  NANDN U14806 ( .A(n14481), .B(n14480), .Z(n14482) );
  AND U14807 ( .A(n14483), .B(n14482), .Z(n14630) );
  NANDN U14808 ( .A(n14485), .B(n14484), .Z(n14489) );
  NANDN U14809 ( .A(n14487), .B(n14486), .Z(n14488) );
  AND U14810 ( .A(n14489), .B(n14488), .Z(n14628) );
  NANDN U14811 ( .A(n14491), .B(n14490), .Z(n14495) );
  NANDN U14812 ( .A(n14493), .B(n14492), .Z(n14494) );
  AND U14813 ( .A(n14495), .B(n14494), .Z(n14636) );
  NANDN U14814 ( .A(n14497), .B(n14496), .Z(n14501) );
  NANDN U14815 ( .A(n14499), .B(n14498), .Z(n14500) );
  AND U14816 ( .A(n14501), .B(n14500), .Z(n14764) );
  NANDN U14817 ( .A(n14503), .B(n14502), .Z(n14507) );
  NAND U14818 ( .A(n14505), .B(n14504), .Z(n14506) );
  AND U14819 ( .A(n14507), .B(n14506), .Z(n14763) );
  XNOR U14820 ( .A(n14764), .B(n14763), .Z(n14766) );
  NANDN U14821 ( .A(n14509), .B(n14508), .Z(n14513) );
  NANDN U14822 ( .A(n14511), .B(n14510), .Z(n14512) );
  AND U14823 ( .A(n14513), .B(n14512), .Z(n14711) );
  NANDN U14824 ( .A(n19237), .B(n14514), .Z(n14516) );
  XOR U14825 ( .A(b[27]), .B(a[87]), .Z(n14657) );
  NANDN U14826 ( .A(n19277), .B(n14657), .Z(n14515) );
  AND U14827 ( .A(n14516), .B(n14515), .Z(n14718) );
  NANDN U14828 ( .A(n17072), .B(n14517), .Z(n14519) );
  XOR U14829 ( .A(a[109]), .B(b[5]), .Z(n14660) );
  NANDN U14830 ( .A(n17223), .B(n14660), .Z(n14518) );
  AND U14831 ( .A(n14519), .B(n14518), .Z(n14716) );
  NANDN U14832 ( .A(n18673), .B(n14520), .Z(n14522) );
  XOR U14833 ( .A(b[19]), .B(a[95]), .Z(n14663) );
  NANDN U14834 ( .A(n18758), .B(n14663), .Z(n14521) );
  NAND U14835 ( .A(n14522), .B(n14521), .Z(n14715) );
  XNOR U14836 ( .A(n14716), .B(n14715), .Z(n14717) );
  XNOR U14837 ( .A(n14718), .B(n14717), .Z(n14709) );
  NANDN U14838 ( .A(n19425), .B(n14523), .Z(n14525) );
  XOR U14839 ( .A(b[31]), .B(a[83]), .Z(n14666) );
  NANDN U14840 ( .A(n19426), .B(n14666), .Z(n14524) );
  AND U14841 ( .A(n14525), .B(n14524), .Z(n14678) );
  NANDN U14842 ( .A(n17067), .B(n14526), .Z(n14528) );
  XOR U14843 ( .A(a[111]), .B(b[3]), .Z(n14669) );
  NANDN U14844 ( .A(n17068), .B(n14669), .Z(n14527) );
  AND U14845 ( .A(n14528), .B(n14527), .Z(n14676) );
  NANDN U14846 ( .A(n18514), .B(n14529), .Z(n14531) );
  XOR U14847 ( .A(b[17]), .B(a[97]), .Z(n14672) );
  NANDN U14848 ( .A(n18585), .B(n14672), .Z(n14530) );
  NAND U14849 ( .A(n14531), .B(n14530), .Z(n14675) );
  XNOR U14850 ( .A(n14676), .B(n14675), .Z(n14677) );
  XOR U14851 ( .A(n14678), .B(n14677), .Z(n14710) );
  XOR U14852 ( .A(n14709), .B(n14710), .Z(n14712) );
  XOR U14853 ( .A(n14711), .B(n14712), .Z(n14646) );
  NANDN U14854 ( .A(n14533), .B(n14532), .Z(n14537) );
  NANDN U14855 ( .A(n14535), .B(n14534), .Z(n14536) );
  AND U14856 ( .A(n14537), .B(n14536), .Z(n14699) );
  NANDN U14857 ( .A(n14539), .B(n14538), .Z(n14543) );
  NANDN U14858 ( .A(n14541), .B(n14540), .Z(n14542) );
  NAND U14859 ( .A(n14543), .B(n14542), .Z(n14700) );
  XNOR U14860 ( .A(n14699), .B(n14700), .Z(n14701) );
  NANDN U14861 ( .A(n14545), .B(n14544), .Z(n14549) );
  NANDN U14862 ( .A(n14547), .B(n14546), .Z(n14548) );
  NAND U14863 ( .A(n14549), .B(n14548), .Z(n14702) );
  XNOR U14864 ( .A(n14701), .B(n14702), .Z(n14645) );
  XNOR U14865 ( .A(n14646), .B(n14645), .Z(n14648) );
  NANDN U14866 ( .A(n14551), .B(n14550), .Z(n14555) );
  NANDN U14867 ( .A(n14553), .B(n14552), .Z(n14554) );
  AND U14868 ( .A(n14555), .B(n14554), .Z(n14647) );
  XOR U14869 ( .A(n14648), .B(n14647), .Z(n14760) );
  NANDN U14870 ( .A(n14557), .B(n14556), .Z(n14561) );
  NANDN U14871 ( .A(n14559), .B(n14558), .Z(n14560) );
  AND U14872 ( .A(n14561), .B(n14560), .Z(n14757) );
  NANDN U14873 ( .A(n14563), .B(n14562), .Z(n14567) );
  NANDN U14874 ( .A(n14565), .B(n14564), .Z(n14566) );
  AND U14875 ( .A(n14567), .B(n14566), .Z(n14642) );
  NANDN U14876 ( .A(n14569), .B(n14568), .Z(n14573) );
  OR U14877 ( .A(n14571), .B(n14570), .Z(n14572) );
  AND U14878 ( .A(n14573), .B(n14572), .Z(n14640) );
  NANDN U14879 ( .A(n14575), .B(n14574), .Z(n14579) );
  NANDN U14880 ( .A(n14577), .B(n14576), .Z(n14578) );
  AND U14881 ( .A(n14579), .B(n14578), .Z(n14706) );
  NANDN U14882 ( .A(n14581), .B(n14580), .Z(n14585) );
  NANDN U14883 ( .A(n14583), .B(n14582), .Z(n14584) );
  NAND U14884 ( .A(n14585), .B(n14584), .Z(n14705) );
  XNOR U14885 ( .A(n14706), .B(n14705), .Z(n14708) );
  NAND U14886 ( .A(b[0]), .B(a[113]), .Z(n14586) );
  XNOR U14887 ( .A(b[1]), .B(n14586), .Z(n14588) );
  NANDN U14888 ( .A(b[0]), .B(a[112]), .Z(n14587) );
  NAND U14889 ( .A(n14588), .B(n14587), .Z(n14654) );
  NANDN U14890 ( .A(n19394), .B(n14589), .Z(n14591) );
  XOR U14891 ( .A(b[29]), .B(a[85]), .Z(n14730) );
  NANDN U14892 ( .A(n19395), .B(n14730), .Z(n14590) );
  AND U14893 ( .A(n14591), .B(n14590), .Z(n14652) );
  AND U14894 ( .A(b[31]), .B(a[81]), .Z(n14651) );
  XNOR U14895 ( .A(n14652), .B(n14651), .Z(n14653) );
  XNOR U14896 ( .A(n14654), .B(n14653), .Z(n14694) );
  NANDN U14897 ( .A(n19005), .B(n14592), .Z(n14594) );
  XOR U14898 ( .A(b[23]), .B(a[91]), .Z(n14733) );
  NANDN U14899 ( .A(n19055), .B(n14733), .Z(n14593) );
  AND U14900 ( .A(n14594), .B(n14593), .Z(n14723) );
  NANDN U14901 ( .A(n17362), .B(n14595), .Z(n14597) );
  XOR U14902 ( .A(a[107]), .B(b[7]), .Z(n14736) );
  NANDN U14903 ( .A(n17522), .B(n14736), .Z(n14596) );
  AND U14904 ( .A(n14597), .B(n14596), .Z(n14722) );
  NANDN U14905 ( .A(n19116), .B(n14598), .Z(n14600) );
  XOR U14906 ( .A(b[25]), .B(a[89]), .Z(n14739) );
  NANDN U14907 ( .A(n19179), .B(n14739), .Z(n14599) );
  NAND U14908 ( .A(n14600), .B(n14599), .Z(n14721) );
  XOR U14909 ( .A(n14722), .B(n14721), .Z(n14724) );
  XOR U14910 ( .A(n14723), .B(n14724), .Z(n14693) );
  XOR U14911 ( .A(n14694), .B(n14693), .Z(n14696) );
  NANDN U14912 ( .A(n18113), .B(n14601), .Z(n14603) );
  XOR U14913 ( .A(b[13]), .B(a[101]), .Z(n14742) );
  NANDN U14914 ( .A(n18229), .B(n14742), .Z(n14602) );
  AND U14915 ( .A(n14603), .B(n14602), .Z(n14688) );
  NANDN U14916 ( .A(n17888), .B(n14604), .Z(n14606) );
  XOR U14917 ( .A(b[11]), .B(a[103]), .Z(n14745) );
  NANDN U14918 ( .A(n18025), .B(n14745), .Z(n14605) );
  NAND U14919 ( .A(n14606), .B(n14605), .Z(n14687) );
  XNOR U14920 ( .A(n14688), .B(n14687), .Z(n14690) );
  NANDN U14921 ( .A(n18487), .B(n14607), .Z(n14609) );
  XOR U14922 ( .A(b[15]), .B(a[99]), .Z(n14748) );
  NANDN U14923 ( .A(n18311), .B(n14748), .Z(n14608) );
  AND U14924 ( .A(n14609), .B(n14608), .Z(n14684) );
  NANDN U14925 ( .A(n18853), .B(n14610), .Z(n14612) );
  XOR U14926 ( .A(b[21]), .B(a[93]), .Z(n14751) );
  NANDN U14927 ( .A(n18926), .B(n14751), .Z(n14611) );
  AND U14928 ( .A(n14612), .B(n14611), .Z(n14682) );
  NANDN U14929 ( .A(n17613), .B(n14613), .Z(n14615) );
  XOR U14930 ( .A(b[9]), .B(a[105]), .Z(n14754) );
  NANDN U14931 ( .A(n17739), .B(n14754), .Z(n14614) );
  NAND U14932 ( .A(n14615), .B(n14614), .Z(n14681) );
  XNOR U14933 ( .A(n14682), .B(n14681), .Z(n14683) );
  XNOR U14934 ( .A(n14684), .B(n14683), .Z(n14689) );
  XOR U14935 ( .A(n14690), .B(n14689), .Z(n14695) );
  XOR U14936 ( .A(n14696), .B(n14695), .Z(n14707) );
  XOR U14937 ( .A(n14708), .B(n14707), .Z(n14639) );
  XNOR U14938 ( .A(n14640), .B(n14639), .Z(n14641) );
  XOR U14939 ( .A(n14642), .B(n14641), .Z(n14758) );
  XNOR U14940 ( .A(n14757), .B(n14758), .Z(n14759) );
  XNOR U14941 ( .A(n14760), .B(n14759), .Z(n14765) );
  XOR U14942 ( .A(n14766), .B(n14765), .Z(n14634) );
  NANDN U14943 ( .A(n14617), .B(n14616), .Z(n14621) );
  OR U14944 ( .A(n14619), .B(n14618), .Z(n14620) );
  AND U14945 ( .A(n14621), .B(n14620), .Z(n14633) );
  XNOR U14946 ( .A(n14634), .B(n14633), .Z(n14635) );
  XNOR U14947 ( .A(n14636), .B(n14635), .Z(n14627) );
  XNOR U14948 ( .A(n14628), .B(n14627), .Z(n14629) );
  XNOR U14949 ( .A(n14630), .B(n14629), .Z(n14769) );
  XNOR U14950 ( .A(sreg[209]), .B(n14769), .Z(n14771) );
  NANDN U14951 ( .A(sreg[208]), .B(n14622), .Z(n14626) );
  NAND U14952 ( .A(n14624), .B(n14623), .Z(n14625) );
  NAND U14953 ( .A(n14626), .B(n14625), .Z(n14770) );
  XNOR U14954 ( .A(n14771), .B(n14770), .Z(c[209]) );
  NANDN U14955 ( .A(n14628), .B(n14627), .Z(n14632) );
  NANDN U14956 ( .A(n14630), .B(n14629), .Z(n14631) );
  AND U14957 ( .A(n14632), .B(n14631), .Z(n14777) );
  NANDN U14958 ( .A(n14634), .B(n14633), .Z(n14638) );
  NANDN U14959 ( .A(n14636), .B(n14635), .Z(n14637) );
  AND U14960 ( .A(n14638), .B(n14637), .Z(n14775) );
  NANDN U14961 ( .A(n14640), .B(n14639), .Z(n14644) );
  NANDN U14962 ( .A(n14642), .B(n14641), .Z(n14643) );
  AND U14963 ( .A(n14644), .B(n14643), .Z(n14913) );
  NANDN U14964 ( .A(n14646), .B(n14645), .Z(n14650) );
  NAND U14965 ( .A(n14648), .B(n14647), .Z(n14649) );
  AND U14966 ( .A(n14650), .B(n14649), .Z(n14912) );
  XNOR U14967 ( .A(n14913), .B(n14912), .Z(n14915) );
  NANDN U14968 ( .A(n14652), .B(n14651), .Z(n14656) );
  NANDN U14969 ( .A(n14654), .B(n14653), .Z(n14655) );
  AND U14970 ( .A(n14656), .B(n14655), .Z(n14848) );
  NANDN U14971 ( .A(n19237), .B(n14657), .Z(n14659) );
  XOR U14972 ( .A(b[27]), .B(a[88]), .Z(n14792) );
  NANDN U14973 ( .A(n19277), .B(n14792), .Z(n14658) );
  AND U14974 ( .A(n14659), .B(n14658), .Z(n14855) );
  NANDN U14975 ( .A(n17072), .B(n14660), .Z(n14662) );
  XOR U14976 ( .A(a[110]), .B(b[5]), .Z(n14795) );
  NANDN U14977 ( .A(n17223), .B(n14795), .Z(n14661) );
  AND U14978 ( .A(n14662), .B(n14661), .Z(n14853) );
  NANDN U14979 ( .A(n18673), .B(n14663), .Z(n14665) );
  XOR U14980 ( .A(b[19]), .B(a[96]), .Z(n14798) );
  NANDN U14981 ( .A(n18758), .B(n14798), .Z(n14664) );
  NAND U14982 ( .A(n14665), .B(n14664), .Z(n14852) );
  XNOR U14983 ( .A(n14853), .B(n14852), .Z(n14854) );
  XNOR U14984 ( .A(n14855), .B(n14854), .Z(n14846) );
  NANDN U14985 ( .A(n19425), .B(n14666), .Z(n14668) );
  XOR U14986 ( .A(b[31]), .B(a[84]), .Z(n14801) );
  NANDN U14987 ( .A(n19426), .B(n14801), .Z(n14667) );
  AND U14988 ( .A(n14668), .B(n14667), .Z(n14813) );
  NANDN U14989 ( .A(n17067), .B(n14669), .Z(n14671) );
  XOR U14990 ( .A(a[112]), .B(b[3]), .Z(n14804) );
  NANDN U14991 ( .A(n17068), .B(n14804), .Z(n14670) );
  AND U14992 ( .A(n14671), .B(n14670), .Z(n14811) );
  NANDN U14993 ( .A(n18514), .B(n14672), .Z(n14674) );
  XOR U14994 ( .A(b[17]), .B(a[98]), .Z(n14807) );
  NANDN U14995 ( .A(n18585), .B(n14807), .Z(n14673) );
  NAND U14996 ( .A(n14674), .B(n14673), .Z(n14810) );
  XNOR U14997 ( .A(n14811), .B(n14810), .Z(n14812) );
  XOR U14998 ( .A(n14813), .B(n14812), .Z(n14847) );
  XOR U14999 ( .A(n14846), .B(n14847), .Z(n14849) );
  XOR U15000 ( .A(n14848), .B(n14849), .Z(n14895) );
  NANDN U15001 ( .A(n14676), .B(n14675), .Z(n14680) );
  NANDN U15002 ( .A(n14678), .B(n14677), .Z(n14679) );
  AND U15003 ( .A(n14680), .B(n14679), .Z(n14834) );
  NANDN U15004 ( .A(n14682), .B(n14681), .Z(n14686) );
  NANDN U15005 ( .A(n14684), .B(n14683), .Z(n14685) );
  NAND U15006 ( .A(n14686), .B(n14685), .Z(n14835) );
  XNOR U15007 ( .A(n14834), .B(n14835), .Z(n14836) );
  NANDN U15008 ( .A(n14688), .B(n14687), .Z(n14692) );
  NAND U15009 ( .A(n14690), .B(n14689), .Z(n14691) );
  NAND U15010 ( .A(n14692), .B(n14691), .Z(n14837) );
  XNOR U15011 ( .A(n14836), .B(n14837), .Z(n14894) );
  XNOR U15012 ( .A(n14895), .B(n14894), .Z(n14897) );
  NAND U15013 ( .A(n14694), .B(n14693), .Z(n14698) );
  NAND U15014 ( .A(n14696), .B(n14695), .Z(n14697) );
  AND U15015 ( .A(n14698), .B(n14697), .Z(n14896) );
  XOR U15016 ( .A(n14897), .B(n14896), .Z(n14909) );
  NANDN U15017 ( .A(n14700), .B(n14699), .Z(n14704) );
  NANDN U15018 ( .A(n14702), .B(n14701), .Z(n14703) );
  AND U15019 ( .A(n14704), .B(n14703), .Z(n14906) );
  NANDN U15020 ( .A(n14710), .B(n14709), .Z(n14714) );
  OR U15021 ( .A(n14712), .B(n14711), .Z(n14713) );
  AND U15022 ( .A(n14714), .B(n14713), .Z(n14901) );
  NANDN U15023 ( .A(n14716), .B(n14715), .Z(n14720) );
  NANDN U15024 ( .A(n14718), .B(n14717), .Z(n14719) );
  AND U15025 ( .A(n14720), .B(n14719), .Z(n14841) );
  NANDN U15026 ( .A(n14722), .B(n14721), .Z(n14726) );
  OR U15027 ( .A(n14724), .B(n14723), .Z(n14725) );
  NAND U15028 ( .A(n14726), .B(n14725), .Z(n14840) );
  XNOR U15029 ( .A(n14841), .B(n14840), .Z(n14842) );
  NAND U15030 ( .A(b[0]), .B(a[114]), .Z(n14727) );
  XNOR U15031 ( .A(b[1]), .B(n14727), .Z(n14729) );
  NANDN U15032 ( .A(b[0]), .B(a[113]), .Z(n14728) );
  NAND U15033 ( .A(n14729), .B(n14728), .Z(n14789) );
  NANDN U15034 ( .A(n19394), .B(n14730), .Z(n14732) );
  XOR U15035 ( .A(b[29]), .B(a[86]), .Z(n14864) );
  NANDN U15036 ( .A(n19395), .B(n14864), .Z(n14731) );
  AND U15037 ( .A(n14732), .B(n14731), .Z(n14787) );
  AND U15038 ( .A(b[31]), .B(a[82]), .Z(n14786) );
  XNOR U15039 ( .A(n14787), .B(n14786), .Z(n14788) );
  XNOR U15040 ( .A(n14789), .B(n14788), .Z(n14828) );
  NANDN U15041 ( .A(n19005), .B(n14733), .Z(n14735) );
  XOR U15042 ( .A(b[23]), .B(a[92]), .Z(n14870) );
  NANDN U15043 ( .A(n19055), .B(n14870), .Z(n14734) );
  AND U15044 ( .A(n14735), .B(n14734), .Z(n14861) );
  NANDN U15045 ( .A(n17362), .B(n14736), .Z(n14738) );
  XOR U15046 ( .A(a[108]), .B(b[7]), .Z(n14873) );
  NANDN U15047 ( .A(n17522), .B(n14873), .Z(n14737) );
  AND U15048 ( .A(n14738), .B(n14737), .Z(n14859) );
  NANDN U15049 ( .A(n19116), .B(n14739), .Z(n14741) );
  XOR U15050 ( .A(b[25]), .B(a[90]), .Z(n14876) );
  NANDN U15051 ( .A(n19179), .B(n14876), .Z(n14740) );
  NAND U15052 ( .A(n14741), .B(n14740), .Z(n14858) );
  XNOR U15053 ( .A(n14859), .B(n14858), .Z(n14860) );
  XOR U15054 ( .A(n14861), .B(n14860), .Z(n14829) );
  XNOR U15055 ( .A(n14828), .B(n14829), .Z(n14830) );
  NANDN U15056 ( .A(n18113), .B(n14742), .Z(n14744) );
  XOR U15057 ( .A(b[13]), .B(a[102]), .Z(n14879) );
  NANDN U15058 ( .A(n18229), .B(n14879), .Z(n14743) );
  AND U15059 ( .A(n14744), .B(n14743), .Z(n14823) );
  NANDN U15060 ( .A(n17888), .B(n14745), .Z(n14747) );
  XOR U15061 ( .A(b[11]), .B(a[104]), .Z(n14882) );
  NANDN U15062 ( .A(n18025), .B(n14882), .Z(n14746) );
  NAND U15063 ( .A(n14747), .B(n14746), .Z(n14822) );
  XNOR U15064 ( .A(n14823), .B(n14822), .Z(n14824) );
  NANDN U15065 ( .A(n18487), .B(n14748), .Z(n14750) );
  XOR U15066 ( .A(b[15]), .B(a[100]), .Z(n14885) );
  NANDN U15067 ( .A(n18311), .B(n14885), .Z(n14749) );
  AND U15068 ( .A(n14750), .B(n14749), .Z(n14819) );
  NANDN U15069 ( .A(n18853), .B(n14751), .Z(n14753) );
  XOR U15070 ( .A(b[21]), .B(a[94]), .Z(n14888) );
  NANDN U15071 ( .A(n18926), .B(n14888), .Z(n14752) );
  AND U15072 ( .A(n14753), .B(n14752), .Z(n14817) );
  NANDN U15073 ( .A(n17613), .B(n14754), .Z(n14756) );
  XOR U15074 ( .A(b[9]), .B(a[106]), .Z(n14891) );
  NANDN U15075 ( .A(n17739), .B(n14891), .Z(n14755) );
  NAND U15076 ( .A(n14756), .B(n14755), .Z(n14816) );
  XNOR U15077 ( .A(n14817), .B(n14816), .Z(n14818) );
  XOR U15078 ( .A(n14819), .B(n14818), .Z(n14825) );
  XOR U15079 ( .A(n14824), .B(n14825), .Z(n14831) );
  XOR U15080 ( .A(n14830), .B(n14831), .Z(n14843) );
  XNOR U15081 ( .A(n14842), .B(n14843), .Z(n14900) );
  XNOR U15082 ( .A(n14901), .B(n14900), .Z(n14902) );
  XOR U15083 ( .A(n14903), .B(n14902), .Z(n14907) );
  XNOR U15084 ( .A(n14906), .B(n14907), .Z(n14908) );
  XNOR U15085 ( .A(n14909), .B(n14908), .Z(n14914) );
  XOR U15086 ( .A(n14915), .B(n14914), .Z(n14781) );
  NANDN U15087 ( .A(n14758), .B(n14757), .Z(n14762) );
  NANDN U15088 ( .A(n14760), .B(n14759), .Z(n14761) );
  AND U15089 ( .A(n14762), .B(n14761), .Z(n14780) );
  XNOR U15090 ( .A(n14781), .B(n14780), .Z(n14782) );
  NANDN U15091 ( .A(n14764), .B(n14763), .Z(n14768) );
  NAND U15092 ( .A(n14766), .B(n14765), .Z(n14767) );
  NAND U15093 ( .A(n14768), .B(n14767), .Z(n14783) );
  XNOR U15094 ( .A(n14782), .B(n14783), .Z(n14774) );
  XNOR U15095 ( .A(n14775), .B(n14774), .Z(n14776) );
  XNOR U15096 ( .A(n14777), .B(n14776), .Z(n14918) );
  XNOR U15097 ( .A(sreg[210]), .B(n14918), .Z(n14920) );
  NANDN U15098 ( .A(sreg[209]), .B(n14769), .Z(n14773) );
  NAND U15099 ( .A(n14771), .B(n14770), .Z(n14772) );
  NAND U15100 ( .A(n14773), .B(n14772), .Z(n14919) );
  XNOR U15101 ( .A(n14920), .B(n14919), .Z(c[210]) );
  NANDN U15102 ( .A(n14775), .B(n14774), .Z(n14779) );
  NANDN U15103 ( .A(n14777), .B(n14776), .Z(n14778) );
  AND U15104 ( .A(n14779), .B(n14778), .Z(n14926) );
  NANDN U15105 ( .A(n14781), .B(n14780), .Z(n14785) );
  NANDN U15106 ( .A(n14783), .B(n14782), .Z(n14784) );
  AND U15107 ( .A(n14785), .B(n14784), .Z(n14924) );
  NANDN U15108 ( .A(n14787), .B(n14786), .Z(n14791) );
  NANDN U15109 ( .A(n14789), .B(n14788), .Z(n14790) );
  AND U15110 ( .A(n14791), .B(n14790), .Z(n15015) );
  NANDN U15111 ( .A(n19237), .B(n14792), .Z(n14794) );
  XOR U15112 ( .A(b[27]), .B(a[89]), .Z(n14959) );
  NANDN U15113 ( .A(n19277), .B(n14959), .Z(n14793) );
  AND U15114 ( .A(n14794), .B(n14793), .Z(n15022) );
  NANDN U15115 ( .A(n17072), .B(n14795), .Z(n14797) );
  XOR U15116 ( .A(a[111]), .B(b[5]), .Z(n14962) );
  NANDN U15117 ( .A(n17223), .B(n14962), .Z(n14796) );
  AND U15118 ( .A(n14797), .B(n14796), .Z(n15020) );
  NANDN U15119 ( .A(n18673), .B(n14798), .Z(n14800) );
  XOR U15120 ( .A(b[19]), .B(a[97]), .Z(n14965) );
  NANDN U15121 ( .A(n18758), .B(n14965), .Z(n14799) );
  NAND U15122 ( .A(n14800), .B(n14799), .Z(n15019) );
  XNOR U15123 ( .A(n15020), .B(n15019), .Z(n15021) );
  XNOR U15124 ( .A(n15022), .B(n15021), .Z(n15013) );
  NANDN U15125 ( .A(n19425), .B(n14801), .Z(n14803) );
  XOR U15126 ( .A(b[31]), .B(a[85]), .Z(n14968) );
  NANDN U15127 ( .A(n19426), .B(n14968), .Z(n14802) );
  AND U15128 ( .A(n14803), .B(n14802), .Z(n14980) );
  NANDN U15129 ( .A(n17067), .B(n14804), .Z(n14806) );
  XOR U15130 ( .A(a[113]), .B(b[3]), .Z(n14971) );
  NANDN U15131 ( .A(n17068), .B(n14971), .Z(n14805) );
  AND U15132 ( .A(n14806), .B(n14805), .Z(n14978) );
  NANDN U15133 ( .A(n18514), .B(n14807), .Z(n14809) );
  XOR U15134 ( .A(b[17]), .B(a[99]), .Z(n14974) );
  NANDN U15135 ( .A(n18585), .B(n14974), .Z(n14808) );
  NAND U15136 ( .A(n14809), .B(n14808), .Z(n14977) );
  XNOR U15137 ( .A(n14978), .B(n14977), .Z(n14979) );
  XOR U15138 ( .A(n14980), .B(n14979), .Z(n15014) );
  XOR U15139 ( .A(n15013), .B(n15014), .Z(n15016) );
  XOR U15140 ( .A(n15015), .B(n15016), .Z(n14948) );
  NANDN U15141 ( .A(n14811), .B(n14810), .Z(n14815) );
  NANDN U15142 ( .A(n14813), .B(n14812), .Z(n14814) );
  AND U15143 ( .A(n14815), .B(n14814), .Z(n15001) );
  NANDN U15144 ( .A(n14817), .B(n14816), .Z(n14821) );
  NANDN U15145 ( .A(n14819), .B(n14818), .Z(n14820) );
  NAND U15146 ( .A(n14821), .B(n14820), .Z(n15002) );
  XNOR U15147 ( .A(n15001), .B(n15002), .Z(n15003) );
  NANDN U15148 ( .A(n14823), .B(n14822), .Z(n14827) );
  NANDN U15149 ( .A(n14825), .B(n14824), .Z(n14826) );
  NAND U15150 ( .A(n14827), .B(n14826), .Z(n15004) );
  XNOR U15151 ( .A(n15003), .B(n15004), .Z(n14947) );
  XNOR U15152 ( .A(n14948), .B(n14947), .Z(n14950) );
  NANDN U15153 ( .A(n14829), .B(n14828), .Z(n14833) );
  NANDN U15154 ( .A(n14831), .B(n14830), .Z(n14832) );
  AND U15155 ( .A(n14833), .B(n14832), .Z(n14949) );
  XOR U15156 ( .A(n14950), .B(n14949), .Z(n15063) );
  NANDN U15157 ( .A(n14835), .B(n14834), .Z(n14839) );
  NANDN U15158 ( .A(n14837), .B(n14836), .Z(n14838) );
  AND U15159 ( .A(n14839), .B(n14838), .Z(n15061) );
  NANDN U15160 ( .A(n14841), .B(n14840), .Z(n14845) );
  NANDN U15161 ( .A(n14843), .B(n14842), .Z(n14844) );
  AND U15162 ( .A(n14845), .B(n14844), .Z(n14944) );
  NANDN U15163 ( .A(n14847), .B(n14846), .Z(n14851) );
  OR U15164 ( .A(n14849), .B(n14848), .Z(n14850) );
  AND U15165 ( .A(n14851), .B(n14850), .Z(n14942) );
  NANDN U15166 ( .A(n14853), .B(n14852), .Z(n14857) );
  NANDN U15167 ( .A(n14855), .B(n14854), .Z(n14856) );
  AND U15168 ( .A(n14857), .B(n14856), .Z(n15008) );
  NANDN U15169 ( .A(n14859), .B(n14858), .Z(n14863) );
  NANDN U15170 ( .A(n14861), .B(n14860), .Z(n14862) );
  NAND U15171 ( .A(n14863), .B(n14862), .Z(n15007) );
  XNOR U15172 ( .A(n15008), .B(n15007), .Z(n15009) );
  NANDN U15173 ( .A(n19394), .B(n14864), .Z(n14866) );
  XOR U15174 ( .A(b[29]), .B(a[87]), .Z(n15031) );
  NANDN U15175 ( .A(n19395), .B(n15031), .Z(n14865) );
  AND U15176 ( .A(n14866), .B(n14865), .Z(n14954) );
  AND U15177 ( .A(b[31]), .B(a[83]), .Z(n14953) );
  XNOR U15178 ( .A(n14954), .B(n14953), .Z(n14955) );
  NAND U15179 ( .A(b[0]), .B(a[115]), .Z(n14867) );
  XNOR U15180 ( .A(b[1]), .B(n14867), .Z(n14869) );
  NANDN U15181 ( .A(b[0]), .B(a[114]), .Z(n14868) );
  NAND U15182 ( .A(n14869), .B(n14868), .Z(n14956) );
  XNOR U15183 ( .A(n14955), .B(n14956), .Z(n14995) );
  NANDN U15184 ( .A(n19005), .B(n14870), .Z(n14872) );
  XOR U15185 ( .A(b[23]), .B(a[93]), .Z(n15037) );
  NANDN U15186 ( .A(n19055), .B(n15037), .Z(n14871) );
  AND U15187 ( .A(n14872), .B(n14871), .Z(n15028) );
  NANDN U15188 ( .A(n17362), .B(n14873), .Z(n14875) );
  XOR U15189 ( .A(a[109]), .B(b[7]), .Z(n15040) );
  NANDN U15190 ( .A(n17522), .B(n15040), .Z(n14874) );
  AND U15191 ( .A(n14875), .B(n14874), .Z(n15026) );
  NANDN U15192 ( .A(n19116), .B(n14876), .Z(n14878) );
  XOR U15193 ( .A(b[25]), .B(a[91]), .Z(n15043) );
  NANDN U15194 ( .A(n19179), .B(n15043), .Z(n14877) );
  NAND U15195 ( .A(n14878), .B(n14877), .Z(n15025) );
  XNOR U15196 ( .A(n15026), .B(n15025), .Z(n15027) );
  XOR U15197 ( .A(n15028), .B(n15027), .Z(n14996) );
  XNOR U15198 ( .A(n14995), .B(n14996), .Z(n14997) );
  NANDN U15199 ( .A(n18113), .B(n14879), .Z(n14881) );
  XOR U15200 ( .A(b[13]), .B(a[103]), .Z(n15046) );
  NANDN U15201 ( .A(n18229), .B(n15046), .Z(n14880) );
  AND U15202 ( .A(n14881), .B(n14880), .Z(n14990) );
  NANDN U15203 ( .A(n17888), .B(n14882), .Z(n14884) );
  XOR U15204 ( .A(b[11]), .B(a[105]), .Z(n15049) );
  NANDN U15205 ( .A(n18025), .B(n15049), .Z(n14883) );
  NAND U15206 ( .A(n14884), .B(n14883), .Z(n14989) );
  XNOR U15207 ( .A(n14990), .B(n14989), .Z(n14991) );
  NANDN U15208 ( .A(n18487), .B(n14885), .Z(n14887) );
  XOR U15209 ( .A(b[15]), .B(a[101]), .Z(n15052) );
  NANDN U15210 ( .A(n18311), .B(n15052), .Z(n14886) );
  AND U15211 ( .A(n14887), .B(n14886), .Z(n14986) );
  NANDN U15212 ( .A(n18853), .B(n14888), .Z(n14890) );
  XOR U15213 ( .A(b[21]), .B(a[95]), .Z(n15055) );
  NANDN U15214 ( .A(n18926), .B(n15055), .Z(n14889) );
  AND U15215 ( .A(n14890), .B(n14889), .Z(n14984) );
  NANDN U15216 ( .A(n17613), .B(n14891), .Z(n14893) );
  XOR U15217 ( .A(b[9]), .B(a[107]), .Z(n15058) );
  NANDN U15218 ( .A(n17739), .B(n15058), .Z(n14892) );
  NAND U15219 ( .A(n14893), .B(n14892), .Z(n14983) );
  XNOR U15220 ( .A(n14984), .B(n14983), .Z(n14985) );
  XOR U15221 ( .A(n14986), .B(n14985), .Z(n14992) );
  XOR U15222 ( .A(n14991), .B(n14992), .Z(n14998) );
  XOR U15223 ( .A(n14997), .B(n14998), .Z(n15010) );
  XNOR U15224 ( .A(n15009), .B(n15010), .Z(n14941) );
  XNOR U15225 ( .A(n14942), .B(n14941), .Z(n14943) );
  XOR U15226 ( .A(n14944), .B(n14943), .Z(n15062) );
  XOR U15227 ( .A(n15061), .B(n15062), .Z(n15064) );
  XOR U15228 ( .A(n15063), .B(n15064), .Z(n14938) );
  NANDN U15229 ( .A(n14895), .B(n14894), .Z(n14899) );
  NAND U15230 ( .A(n14897), .B(n14896), .Z(n14898) );
  AND U15231 ( .A(n14899), .B(n14898), .Z(n14936) );
  NANDN U15232 ( .A(n14901), .B(n14900), .Z(n14905) );
  NANDN U15233 ( .A(n14903), .B(n14902), .Z(n14904) );
  AND U15234 ( .A(n14905), .B(n14904), .Z(n14935) );
  XNOR U15235 ( .A(n14936), .B(n14935), .Z(n14937) );
  XNOR U15236 ( .A(n14938), .B(n14937), .Z(n14929) );
  NANDN U15237 ( .A(n14907), .B(n14906), .Z(n14911) );
  NANDN U15238 ( .A(n14909), .B(n14908), .Z(n14910) );
  NAND U15239 ( .A(n14911), .B(n14910), .Z(n14930) );
  XNOR U15240 ( .A(n14929), .B(n14930), .Z(n14931) );
  NANDN U15241 ( .A(n14913), .B(n14912), .Z(n14917) );
  NAND U15242 ( .A(n14915), .B(n14914), .Z(n14916) );
  NAND U15243 ( .A(n14917), .B(n14916), .Z(n14932) );
  XNOR U15244 ( .A(n14931), .B(n14932), .Z(n14923) );
  XNOR U15245 ( .A(n14924), .B(n14923), .Z(n14925) );
  XNOR U15246 ( .A(n14926), .B(n14925), .Z(n15067) );
  XNOR U15247 ( .A(sreg[211]), .B(n15067), .Z(n15069) );
  NANDN U15248 ( .A(sreg[210]), .B(n14918), .Z(n14922) );
  NAND U15249 ( .A(n14920), .B(n14919), .Z(n14921) );
  NAND U15250 ( .A(n14922), .B(n14921), .Z(n15068) );
  XNOR U15251 ( .A(n15069), .B(n15068), .Z(c[211]) );
  NANDN U15252 ( .A(n14924), .B(n14923), .Z(n14928) );
  NANDN U15253 ( .A(n14926), .B(n14925), .Z(n14927) );
  AND U15254 ( .A(n14928), .B(n14927), .Z(n15075) );
  NANDN U15255 ( .A(n14930), .B(n14929), .Z(n14934) );
  NANDN U15256 ( .A(n14932), .B(n14931), .Z(n14933) );
  AND U15257 ( .A(n14934), .B(n14933), .Z(n15073) );
  NANDN U15258 ( .A(n14936), .B(n14935), .Z(n14940) );
  NANDN U15259 ( .A(n14938), .B(n14937), .Z(n14939) );
  AND U15260 ( .A(n14940), .B(n14939), .Z(n15081) );
  NANDN U15261 ( .A(n14942), .B(n14941), .Z(n14946) );
  NANDN U15262 ( .A(n14944), .B(n14943), .Z(n14945) );
  AND U15263 ( .A(n14946), .B(n14945), .Z(n15211) );
  NANDN U15264 ( .A(n14948), .B(n14947), .Z(n14952) );
  NAND U15265 ( .A(n14950), .B(n14949), .Z(n14951) );
  AND U15266 ( .A(n14952), .B(n14951), .Z(n15210) );
  XNOR U15267 ( .A(n15211), .B(n15210), .Z(n15213) );
  NANDN U15268 ( .A(n14954), .B(n14953), .Z(n14958) );
  NANDN U15269 ( .A(n14956), .B(n14955), .Z(n14957) );
  AND U15270 ( .A(n14958), .B(n14957), .Z(n15158) );
  NANDN U15271 ( .A(n19237), .B(n14959), .Z(n14961) );
  XOR U15272 ( .A(b[27]), .B(a[90]), .Z(n15102) );
  NANDN U15273 ( .A(n19277), .B(n15102), .Z(n14960) );
  AND U15274 ( .A(n14961), .B(n14960), .Z(n15165) );
  NANDN U15275 ( .A(n17072), .B(n14962), .Z(n14964) );
  XOR U15276 ( .A(a[112]), .B(b[5]), .Z(n15105) );
  NANDN U15277 ( .A(n17223), .B(n15105), .Z(n14963) );
  AND U15278 ( .A(n14964), .B(n14963), .Z(n15163) );
  NANDN U15279 ( .A(n18673), .B(n14965), .Z(n14967) );
  XOR U15280 ( .A(b[19]), .B(a[98]), .Z(n15108) );
  NANDN U15281 ( .A(n18758), .B(n15108), .Z(n14966) );
  NAND U15282 ( .A(n14967), .B(n14966), .Z(n15162) );
  XNOR U15283 ( .A(n15163), .B(n15162), .Z(n15164) );
  XNOR U15284 ( .A(n15165), .B(n15164), .Z(n15156) );
  NANDN U15285 ( .A(n19425), .B(n14968), .Z(n14970) );
  XOR U15286 ( .A(b[31]), .B(a[86]), .Z(n15111) );
  NANDN U15287 ( .A(n19426), .B(n15111), .Z(n14969) );
  AND U15288 ( .A(n14970), .B(n14969), .Z(n15123) );
  NANDN U15289 ( .A(n17067), .B(n14971), .Z(n14973) );
  XOR U15290 ( .A(a[114]), .B(b[3]), .Z(n15114) );
  NANDN U15291 ( .A(n17068), .B(n15114), .Z(n14972) );
  AND U15292 ( .A(n14973), .B(n14972), .Z(n15121) );
  NANDN U15293 ( .A(n18514), .B(n14974), .Z(n14976) );
  XOR U15294 ( .A(b[17]), .B(a[100]), .Z(n15117) );
  NANDN U15295 ( .A(n18585), .B(n15117), .Z(n14975) );
  NAND U15296 ( .A(n14976), .B(n14975), .Z(n15120) );
  XNOR U15297 ( .A(n15121), .B(n15120), .Z(n15122) );
  XOR U15298 ( .A(n15123), .B(n15122), .Z(n15157) );
  XOR U15299 ( .A(n15156), .B(n15157), .Z(n15159) );
  XOR U15300 ( .A(n15158), .B(n15159), .Z(n15091) );
  NANDN U15301 ( .A(n14978), .B(n14977), .Z(n14982) );
  NANDN U15302 ( .A(n14980), .B(n14979), .Z(n14981) );
  AND U15303 ( .A(n14982), .B(n14981), .Z(n15144) );
  NANDN U15304 ( .A(n14984), .B(n14983), .Z(n14988) );
  NANDN U15305 ( .A(n14986), .B(n14985), .Z(n14987) );
  NAND U15306 ( .A(n14988), .B(n14987), .Z(n15145) );
  XNOR U15307 ( .A(n15144), .B(n15145), .Z(n15146) );
  NANDN U15308 ( .A(n14990), .B(n14989), .Z(n14994) );
  NANDN U15309 ( .A(n14992), .B(n14991), .Z(n14993) );
  NAND U15310 ( .A(n14994), .B(n14993), .Z(n15147) );
  XNOR U15311 ( .A(n15146), .B(n15147), .Z(n15090) );
  XNOR U15312 ( .A(n15091), .B(n15090), .Z(n15093) );
  NANDN U15313 ( .A(n14996), .B(n14995), .Z(n15000) );
  NANDN U15314 ( .A(n14998), .B(n14997), .Z(n14999) );
  AND U15315 ( .A(n15000), .B(n14999), .Z(n15092) );
  XOR U15316 ( .A(n15093), .B(n15092), .Z(n15207) );
  NANDN U15317 ( .A(n15002), .B(n15001), .Z(n15006) );
  NANDN U15318 ( .A(n15004), .B(n15003), .Z(n15005) );
  AND U15319 ( .A(n15006), .B(n15005), .Z(n15204) );
  NANDN U15320 ( .A(n15008), .B(n15007), .Z(n15012) );
  NANDN U15321 ( .A(n15010), .B(n15009), .Z(n15011) );
  AND U15322 ( .A(n15012), .B(n15011), .Z(n15087) );
  NANDN U15323 ( .A(n15014), .B(n15013), .Z(n15018) );
  OR U15324 ( .A(n15016), .B(n15015), .Z(n15017) );
  AND U15325 ( .A(n15018), .B(n15017), .Z(n15085) );
  NANDN U15326 ( .A(n15020), .B(n15019), .Z(n15024) );
  NANDN U15327 ( .A(n15022), .B(n15021), .Z(n15023) );
  AND U15328 ( .A(n15024), .B(n15023), .Z(n15151) );
  NANDN U15329 ( .A(n15026), .B(n15025), .Z(n15030) );
  NANDN U15330 ( .A(n15028), .B(n15027), .Z(n15029) );
  NAND U15331 ( .A(n15030), .B(n15029), .Z(n15150) );
  XNOR U15332 ( .A(n15151), .B(n15150), .Z(n15152) );
  NANDN U15333 ( .A(n19394), .B(n15031), .Z(n15033) );
  XOR U15334 ( .A(b[29]), .B(a[88]), .Z(n15174) );
  NANDN U15335 ( .A(n19395), .B(n15174), .Z(n15032) );
  AND U15336 ( .A(n15033), .B(n15032), .Z(n15097) );
  AND U15337 ( .A(b[31]), .B(a[84]), .Z(n15096) );
  XNOR U15338 ( .A(n15097), .B(n15096), .Z(n15098) );
  NAND U15339 ( .A(b[0]), .B(a[116]), .Z(n15034) );
  XNOR U15340 ( .A(b[1]), .B(n15034), .Z(n15036) );
  NANDN U15341 ( .A(b[0]), .B(a[115]), .Z(n15035) );
  NAND U15342 ( .A(n15036), .B(n15035), .Z(n15099) );
  XNOR U15343 ( .A(n15098), .B(n15099), .Z(n15138) );
  NANDN U15344 ( .A(n19005), .B(n15037), .Z(n15039) );
  XOR U15345 ( .A(b[23]), .B(a[94]), .Z(n15180) );
  NANDN U15346 ( .A(n19055), .B(n15180), .Z(n15038) );
  AND U15347 ( .A(n15039), .B(n15038), .Z(n15171) );
  NANDN U15348 ( .A(n17362), .B(n15040), .Z(n15042) );
  XOR U15349 ( .A(a[110]), .B(b[7]), .Z(n15183) );
  NANDN U15350 ( .A(n17522), .B(n15183), .Z(n15041) );
  AND U15351 ( .A(n15042), .B(n15041), .Z(n15169) );
  NANDN U15352 ( .A(n19116), .B(n15043), .Z(n15045) );
  XOR U15353 ( .A(b[25]), .B(a[92]), .Z(n15186) );
  NANDN U15354 ( .A(n19179), .B(n15186), .Z(n15044) );
  NAND U15355 ( .A(n15045), .B(n15044), .Z(n15168) );
  XNOR U15356 ( .A(n15169), .B(n15168), .Z(n15170) );
  XOR U15357 ( .A(n15171), .B(n15170), .Z(n15139) );
  XNOR U15358 ( .A(n15138), .B(n15139), .Z(n15140) );
  NANDN U15359 ( .A(n18113), .B(n15046), .Z(n15048) );
  XOR U15360 ( .A(b[13]), .B(a[104]), .Z(n15189) );
  NANDN U15361 ( .A(n18229), .B(n15189), .Z(n15047) );
  AND U15362 ( .A(n15048), .B(n15047), .Z(n15133) );
  NANDN U15363 ( .A(n17888), .B(n15049), .Z(n15051) );
  XOR U15364 ( .A(b[11]), .B(a[106]), .Z(n15192) );
  NANDN U15365 ( .A(n18025), .B(n15192), .Z(n15050) );
  NAND U15366 ( .A(n15051), .B(n15050), .Z(n15132) );
  XNOR U15367 ( .A(n15133), .B(n15132), .Z(n15134) );
  NANDN U15368 ( .A(n18487), .B(n15052), .Z(n15054) );
  XOR U15369 ( .A(b[15]), .B(a[102]), .Z(n15195) );
  NANDN U15370 ( .A(n18311), .B(n15195), .Z(n15053) );
  AND U15371 ( .A(n15054), .B(n15053), .Z(n15129) );
  NANDN U15372 ( .A(n18853), .B(n15055), .Z(n15057) );
  XOR U15373 ( .A(b[21]), .B(a[96]), .Z(n15198) );
  NANDN U15374 ( .A(n18926), .B(n15198), .Z(n15056) );
  AND U15375 ( .A(n15057), .B(n15056), .Z(n15127) );
  NANDN U15376 ( .A(n17613), .B(n15058), .Z(n15060) );
  XOR U15377 ( .A(a[108]), .B(b[9]), .Z(n15201) );
  NANDN U15378 ( .A(n17739), .B(n15201), .Z(n15059) );
  NAND U15379 ( .A(n15060), .B(n15059), .Z(n15126) );
  XNOR U15380 ( .A(n15127), .B(n15126), .Z(n15128) );
  XOR U15381 ( .A(n15129), .B(n15128), .Z(n15135) );
  XOR U15382 ( .A(n15134), .B(n15135), .Z(n15141) );
  XOR U15383 ( .A(n15140), .B(n15141), .Z(n15153) );
  XNOR U15384 ( .A(n15152), .B(n15153), .Z(n15084) );
  XNOR U15385 ( .A(n15085), .B(n15084), .Z(n15086) );
  XOR U15386 ( .A(n15087), .B(n15086), .Z(n15205) );
  XNOR U15387 ( .A(n15204), .B(n15205), .Z(n15206) );
  XNOR U15388 ( .A(n15207), .B(n15206), .Z(n15212) );
  XOR U15389 ( .A(n15213), .B(n15212), .Z(n15079) );
  NANDN U15390 ( .A(n15062), .B(n15061), .Z(n15066) );
  OR U15391 ( .A(n15064), .B(n15063), .Z(n15065) );
  AND U15392 ( .A(n15066), .B(n15065), .Z(n15078) );
  XNOR U15393 ( .A(n15079), .B(n15078), .Z(n15080) );
  XNOR U15394 ( .A(n15081), .B(n15080), .Z(n15072) );
  XNOR U15395 ( .A(n15073), .B(n15072), .Z(n15074) );
  XNOR U15396 ( .A(n15075), .B(n15074), .Z(n15216) );
  XNOR U15397 ( .A(sreg[212]), .B(n15216), .Z(n15218) );
  NANDN U15398 ( .A(sreg[211]), .B(n15067), .Z(n15071) );
  NAND U15399 ( .A(n15069), .B(n15068), .Z(n15070) );
  NAND U15400 ( .A(n15071), .B(n15070), .Z(n15217) );
  XNOR U15401 ( .A(n15218), .B(n15217), .Z(c[212]) );
  NANDN U15402 ( .A(n15073), .B(n15072), .Z(n15077) );
  NANDN U15403 ( .A(n15075), .B(n15074), .Z(n15076) );
  AND U15404 ( .A(n15077), .B(n15076), .Z(n15224) );
  NANDN U15405 ( .A(n15079), .B(n15078), .Z(n15083) );
  NANDN U15406 ( .A(n15081), .B(n15080), .Z(n15082) );
  AND U15407 ( .A(n15083), .B(n15082), .Z(n15222) );
  NANDN U15408 ( .A(n15085), .B(n15084), .Z(n15089) );
  NANDN U15409 ( .A(n15087), .B(n15086), .Z(n15088) );
  AND U15410 ( .A(n15089), .B(n15088), .Z(n15234) );
  NANDN U15411 ( .A(n15091), .B(n15090), .Z(n15095) );
  NAND U15412 ( .A(n15093), .B(n15092), .Z(n15094) );
  AND U15413 ( .A(n15095), .B(n15094), .Z(n15233) );
  XNOR U15414 ( .A(n15234), .B(n15233), .Z(n15236) );
  NANDN U15415 ( .A(n15097), .B(n15096), .Z(n15101) );
  NANDN U15416 ( .A(n15099), .B(n15098), .Z(n15100) );
  AND U15417 ( .A(n15101), .B(n15100), .Z(n15313) );
  NANDN U15418 ( .A(n19237), .B(n15102), .Z(n15104) );
  XOR U15419 ( .A(b[27]), .B(a[91]), .Z(n15257) );
  NANDN U15420 ( .A(n19277), .B(n15257), .Z(n15103) );
  AND U15421 ( .A(n15104), .B(n15103), .Z(n15320) );
  NANDN U15422 ( .A(n17072), .B(n15105), .Z(n15107) );
  XOR U15423 ( .A(a[113]), .B(b[5]), .Z(n15260) );
  NANDN U15424 ( .A(n17223), .B(n15260), .Z(n15106) );
  AND U15425 ( .A(n15107), .B(n15106), .Z(n15318) );
  NANDN U15426 ( .A(n18673), .B(n15108), .Z(n15110) );
  XOR U15427 ( .A(b[19]), .B(a[99]), .Z(n15263) );
  NANDN U15428 ( .A(n18758), .B(n15263), .Z(n15109) );
  NAND U15429 ( .A(n15110), .B(n15109), .Z(n15317) );
  XNOR U15430 ( .A(n15318), .B(n15317), .Z(n15319) );
  XNOR U15431 ( .A(n15320), .B(n15319), .Z(n15311) );
  NANDN U15432 ( .A(n19425), .B(n15111), .Z(n15113) );
  XOR U15433 ( .A(b[31]), .B(a[87]), .Z(n15266) );
  NANDN U15434 ( .A(n19426), .B(n15266), .Z(n15112) );
  AND U15435 ( .A(n15113), .B(n15112), .Z(n15278) );
  NANDN U15436 ( .A(n17067), .B(n15114), .Z(n15116) );
  XOR U15437 ( .A(a[115]), .B(b[3]), .Z(n15269) );
  NANDN U15438 ( .A(n17068), .B(n15269), .Z(n15115) );
  AND U15439 ( .A(n15116), .B(n15115), .Z(n15276) );
  NANDN U15440 ( .A(n18514), .B(n15117), .Z(n15119) );
  XOR U15441 ( .A(b[17]), .B(a[101]), .Z(n15272) );
  NANDN U15442 ( .A(n18585), .B(n15272), .Z(n15118) );
  NAND U15443 ( .A(n15119), .B(n15118), .Z(n15275) );
  XNOR U15444 ( .A(n15276), .B(n15275), .Z(n15277) );
  XOR U15445 ( .A(n15278), .B(n15277), .Z(n15312) );
  XOR U15446 ( .A(n15311), .B(n15312), .Z(n15314) );
  XOR U15447 ( .A(n15313), .B(n15314), .Z(n15246) );
  NANDN U15448 ( .A(n15121), .B(n15120), .Z(n15125) );
  NANDN U15449 ( .A(n15123), .B(n15122), .Z(n15124) );
  AND U15450 ( .A(n15125), .B(n15124), .Z(n15299) );
  NANDN U15451 ( .A(n15127), .B(n15126), .Z(n15131) );
  NANDN U15452 ( .A(n15129), .B(n15128), .Z(n15130) );
  NAND U15453 ( .A(n15131), .B(n15130), .Z(n15300) );
  XNOR U15454 ( .A(n15299), .B(n15300), .Z(n15301) );
  NANDN U15455 ( .A(n15133), .B(n15132), .Z(n15137) );
  NANDN U15456 ( .A(n15135), .B(n15134), .Z(n15136) );
  NAND U15457 ( .A(n15137), .B(n15136), .Z(n15302) );
  XNOR U15458 ( .A(n15301), .B(n15302), .Z(n15245) );
  XNOR U15459 ( .A(n15246), .B(n15245), .Z(n15248) );
  NANDN U15460 ( .A(n15139), .B(n15138), .Z(n15143) );
  NANDN U15461 ( .A(n15141), .B(n15140), .Z(n15142) );
  AND U15462 ( .A(n15143), .B(n15142), .Z(n15247) );
  XOR U15463 ( .A(n15248), .B(n15247), .Z(n15362) );
  NANDN U15464 ( .A(n15145), .B(n15144), .Z(n15149) );
  NANDN U15465 ( .A(n15147), .B(n15146), .Z(n15148) );
  AND U15466 ( .A(n15149), .B(n15148), .Z(n15359) );
  NANDN U15467 ( .A(n15151), .B(n15150), .Z(n15155) );
  NANDN U15468 ( .A(n15153), .B(n15152), .Z(n15154) );
  AND U15469 ( .A(n15155), .B(n15154), .Z(n15242) );
  NANDN U15470 ( .A(n15157), .B(n15156), .Z(n15161) );
  OR U15471 ( .A(n15159), .B(n15158), .Z(n15160) );
  AND U15472 ( .A(n15161), .B(n15160), .Z(n15240) );
  NANDN U15473 ( .A(n15163), .B(n15162), .Z(n15167) );
  NANDN U15474 ( .A(n15165), .B(n15164), .Z(n15166) );
  AND U15475 ( .A(n15167), .B(n15166), .Z(n15306) );
  NANDN U15476 ( .A(n15169), .B(n15168), .Z(n15173) );
  NANDN U15477 ( .A(n15171), .B(n15170), .Z(n15172) );
  NAND U15478 ( .A(n15173), .B(n15172), .Z(n15305) );
  XNOR U15479 ( .A(n15306), .B(n15305), .Z(n15307) );
  NANDN U15480 ( .A(n19394), .B(n15174), .Z(n15176) );
  XOR U15481 ( .A(b[29]), .B(a[89]), .Z(n15332) );
  NANDN U15482 ( .A(n19395), .B(n15332), .Z(n15175) );
  AND U15483 ( .A(n15176), .B(n15175), .Z(n15252) );
  AND U15484 ( .A(b[31]), .B(a[85]), .Z(n15251) );
  XNOR U15485 ( .A(n15252), .B(n15251), .Z(n15253) );
  NAND U15486 ( .A(b[0]), .B(a[117]), .Z(n15177) );
  XNOR U15487 ( .A(b[1]), .B(n15177), .Z(n15179) );
  NANDN U15488 ( .A(b[0]), .B(a[116]), .Z(n15178) );
  NAND U15489 ( .A(n15179), .B(n15178), .Z(n15254) );
  XNOR U15490 ( .A(n15253), .B(n15254), .Z(n15293) );
  NANDN U15491 ( .A(n19005), .B(n15180), .Z(n15182) );
  XOR U15492 ( .A(b[23]), .B(a[95]), .Z(n15335) );
  NANDN U15493 ( .A(n19055), .B(n15335), .Z(n15181) );
  AND U15494 ( .A(n15182), .B(n15181), .Z(n15326) );
  NANDN U15495 ( .A(n17362), .B(n15183), .Z(n15185) );
  XOR U15496 ( .A(a[111]), .B(b[7]), .Z(n15338) );
  NANDN U15497 ( .A(n17522), .B(n15338), .Z(n15184) );
  AND U15498 ( .A(n15185), .B(n15184), .Z(n15324) );
  NANDN U15499 ( .A(n19116), .B(n15186), .Z(n15188) );
  XOR U15500 ( .A(b[25]), .B(a[93]), .Z(n15341) );
  NANDN U15501 ( .A(n19179), .B(n15341), .Z(n15187) );
  NAND U15502 ( .A(n15188), .B(n15187), .Z(n15323) );
  XNOR U15503 ( .A(n15324), .B(n15323), .Z(n15325) );
  XOR U15504 ( .A(n15326), .B(n15325), .Z(n15294) );
  XNOR U15505 ( .A(n15293), .B(n15294), .Z(n15295) );
  NANDN U15506 ( .A(n18113), .B(n15189), .Z(n15191) );
  XOR U15507 ( .A(b[13]), .B(a[105]), .Z(n15344) );
  NANDN U15508 ( .A(n18229), .B(n15344), .Z(n15190) );
  AND U15509 ( .A(n15191), .B(n15190), .Z(n15288) );
  NANDN U15510 ( .A(n17888), .B(n15192), .Z(n15194) );
  XOR U15511 ( .A(b[11]), .B(a[107]), .Z(n15347) );
  NANDN U15512 ( .A(n18025), .B(n15347), .Z(n15193) );
  NAND U15513 ( .A(n15194), .B(n15193), .Z(n15287) );
  XNOR U15514 ( .A(n15288), .B(n15287), .Z(n15289) );
  NANDN U15515 ( .A(n18487), .B(n15195), .Z(n15197) );
  XOR U15516 ( .A(b[15]), .B(a[103]), .Z(n15350) );
  NANDN U15517 ( .A(n18311), .B(n15350), .Z(n15196) );
  AND U15518 ( .A(n15197), .B(n15196), .Z(n15284) );
  NANDN U15519 ( .A(n18853), .B(n15198), .Z(n15200) );
  XOR U15520 ( .A(b[21]), .B(a[97]), .Z(n15353) );
  NANDN U15521 ( .A(n18926), .B(n15353), .Z(n15199) );
  AND U15522 ( .A(n15200), .B(n15199), .Z(n15282) );
  NANDN U15523 ( .A(n17613), .B(n15201), .Z(n15203) );
  XOR U15524 ( .A(a[109]), .B(b[9]), .Z(n15356) );
  NANDN U15525 ( .A(n17739), .B(n15356), .Z(n15202) );
  NAND U15526 ( .A(n15203), .B(n15202), .Z(n15281) );
  XNOR U15527 ( .A(n15282), .B(n15281), .Z(n15283) );
  XOR U15528 ( .A(n15284), .B(n15283), .Z(n15290) );
  XOR U15529 ( .A(n15289), .B(n15290), .Z(n15296) );
  XOR U15530 ( .A(n15295), .B(n15296), .Z(n15308) );
  XNOR U15531 ( .A(n15307), .B(n15308), .Z(n15239) );
  XNOR U15532 ( .A(n15240), .B(n15239), .Z(n15241) );
  XOR U15533 ( .A(n15242), .B(n15241), .Z(n15360) );
  XNOR U15534 ( .A(n15359), .B(n15360), .Z(n15361) );
  XNOR U15535 ( .A(n15362), .B(n15361), .Z(n15235) );
  XOR U15536 ( .A(n15236), .B(n15235), .Z(n15228) );
  NANDN U15537 ( .A(n15205), .B(n15204), .Z(n15209) );
  NANDN U15538 ( .A(n15207), .B(n15206), .Z(n15208) );
  AND U15539 ( .A(n15209), .B(n15208), .Z(n15227) );
  XNOR U15540 ( .A(n15228), .B(n15227), .Z(n15229) );
  NANDN U15541 ( .A(n15211), .B(n15210), .Z(n15215) );
  NAND U15542 ( .A(n15213), .B(n15212), .Z(n15214) );
  NAND U15543 ( .A(n15215), .B(n15214), .Z(n15230) );
  XNOR U15544 ( .A(n15229), .B(n15230), .Z(n15221) );
  XNOR U15545 ( .A(n15222), .B(n15221), .Z(n15223) );
  XNOR U15546 ( .A(n15224), .B(n15223), .Z(n15365) );
  XNOR U15547 ( .A(sreg[213]), .B(n15365), .Z(n15367) );
  NANDN U15548 ( .A(sreg[212]), .B(n15216), .Z(n15220) );
  NAND U15549 ( .A(n15218), .B(n15217), .Z(n15219) );
  NAND U15550 ( .A(n15220), .B(n15219), .Z(n15366) );
  XNOR U15551 ( .A(n15367), .B(n15366), .Z(c[213]) );
  NANDN U15552 ( .A(n15222), .B(n15221), .Z(n15226) );
  NANDN U15553 ( .A(n15224), .B(n15223), .Z(n15225) );
  AND U15554 ( .A(n15226), .B(n15225), .Z(n15373) );
  NANDN U15555 ( .A(n15228), .B(n15227), .Z(n15232) );
  NANDN U15556 ( .A(n15230), .B(n15229), .Z(n15231) );
  AND U15557 ( .A(n15232), .B(n15231), .Z(n15371) );
  NANDN U15558 ( .A(n15234), .B(n15233), .Z(n15238) );
  NAND U15559 ( .A(n15236), .B(n15235), .Z(n15237) );
  AND U15560 ( .A(n15238), .B(n15237), .Z(n15378) );
  NANDN U15561 ( .A(n15240), .B(n15239), .Z(n15244) );
  NANDN U15562 ( .A(n15242), .B(n15241), .Z(n15243) );
  AND U15563 ( .A(n15244), .B(n15243), .Z(n15383) );
  NANDN U15564 ( .A(n15246), .B(n15245), .Z(n15250) );
  NAND U15565 ( .A(n15248), .B(n15247), .Z(n15249) );
  AND U15566 ( .A(n15250), .B(n15249), .Z(n15382) );
  XNOR U15567 ( .A(n15383), .B(n15382), .Z(n15385) );
  NANDN U15568 ( .A(n15252), .B(n15251), .Z(n15256) );
  NANDN U15569 ( .A(n15254), .B(n15253), .Z(n15255) );
  AND U15570 ( .A(n15256), .B(n15255), .Z(n15462) );
  NANDN U15571 ( .A(n19237), .B(n15257), .Z(n15259) );
  XOR U15572 ( .A(b[27]), .B(a[92]), .Z(n15406) );
  NANDN U15573 ( .A(n19277), .B(n15406), .Z(n15258) );
  AND U15574 ( .A(n15259), .B(n15258), .Z(n15469) );
  NANDN U15575 ( .A(n17072), .B(n15260), .Z(n15262) );
  XOR U15576 ( .A(a[114]), .B(b[5]), .Z(n15409) );
  NANDN U15577 ( .A(n17223), .B(n15409), .Z(n15261) );
  AND U15578 ( .A(n15262), .B(n15261), .Z(n15467) );
  NANDN U15579 ( .A(n18673), .B(n15263), .Z(n15265) );
  XOR U15580 ( .A(b[19]), .B(a[100]), .Z(n15412) );
  NANDN U15581 ( .A(n18758), .B(n15412), .Z(n15264) );
  NAND U15582 ( .A(n15265), .B(n15264), .Z(n15466) );
  XNOR U15583 ( .A(n15467), .B(n15466), .Z(n15468) );
  XNOR U15584 ( .A(n15469), .B(n15468), .Z(n15460) );
  NANDN U15585 ( .A(n19425), .B(n15266), .Z(n15268) );
  XOR U15586 ( .A(b[31]), .B(a[88]), .Z(n15415) );
  NANDN U15587 ( .A(n19426), .B(n15415), .Z(n15267) );
  AND U15588 ( .A(n15268), .B(n15267), .Z(n15427) );
  NANDN U15589 ( .A(n17067), .B(n15269), .Z(n15271) );
  XOR U15590 ( .A(a[116]), .B(b[3]), .Z(n15418) );
  NANDN U15591 ( .A(n17068), .B(n15418), .Z(n15270) );
  AND U15592 ( .A(n15271), .B(n15270), .Z(n15425) );
  NANDN U15593 ( .A(n18514), .B(n15272), .Z(n15274) );
  XOR U15594 ( .A(b[17]), .B(a[102]), .Z(n15421) );
  NANDN U15595 ( .A(n18585), .B(n15421), .Z(n15273) );
  NAND U15596 ( .A(n15274), .B(n15273), .Z(n15424) );
  XNOR U15597 ( .A(n15425), .B(n15424), .Z(n15426) );
  XOR U15598 ( .A(n15427), .B(n15426), .Z(n15461) );
  XOR U15599 ( .A(n15460), .B(n15461), .Z(n15463) );
  XOR U15600 ( .A(n15462), .B(n15463), .Z(n15395) );
  NANDN U15601 ( .A(n15276), .B(n15275), .Z(n15280) );
  NANDN U15602 ( .A(n15278), .B(n15277), .Z(n15279) );
  AND U15603 ( .A(n15280), .B(n15279), .Z(n15448) );
  NANDN U15604 ( .A(n15282), .B(n15281), .Z(n15286) );
  NANDN U15605 ( .A(n15284), .B(n15283), .Z(n15285) );
  NAND U15606 ( .A(n15286), .B(n15285), .Z(n15449) );
  XNOR U15607 ( .A(n15448), .B(n15449), .Z(n15450) );
  NANDN U15608 ( .A(n15288), .B(n15287), .Z(n15292) );
  NANDN U15609 ( .A(n15290), .B(n15289), .Z(n15291) );
  NAND U15610 ( .A(n15292), .B(n15291), .Z(n15451) );
  XNOR U15611 ( .A(n15450), .B(n15451), .Z(n15394) );
  XNOR U15612 ( .A(n15395), .B(n15394), .Z(n15397) );
  NANDN U15613 ( .A(n15294), .B(n15293), .Z(n15298) );
  NANDN U15614 ( .A(n15296), .B(n15295), .Z(n15297) );
  AND U15615 ( .A(n15298), .B(n15297), .Z(n15396) );
  XOR U15616 ( .A(n15397), .B(n15396), .Z(n15511) );
  NANDN U15617 ( .A(n15300), .B(n15299), .Z(n15304) );
  NANDN U15618 ( .A(n15302), .B(n15301), .Z(n15303) );
  AND U15619 ( .A(n15304), .B(n15303), .Z(n15508) );
  NANDN U15620 ( .A(n15306), .B(n15305), .Z(n15310) );
  NANDN U15621 ( .A(n15308), .B(n15307), .Z(n15309) );
  AND U15622 ( .A(n15310), .B(n15309), .Z(n15391) );
  NANDN U15623 ( .A(n15312), .B(n15311), .Z(n15316) );
  OR U15624 ( .A(n15314), .B(n15313), .Z(n15315) );
  AND U15625 ( .A(n15316), .B(n15315), .Z(n15389) );
  NANDN U15626 ( .A(n15318), .B(n15317), .Z(n15322) );
  NANDN U15627 ( .A(n15320), .B(n15319), .Z(n15321) );
  AND U15628 ( .A(n15322), .B(n15321), .Z(n15455) );
  NANDN U15629 ( .A(n15324), .B(n15323), .Z(n15328) );
  NANDN U15630 ( .A(n15326), .B(n15325), .Z(n15327) );
  NAND U15631 ( .A(n15328), .B(n15327), .Z(n15454) );
  XNOR U15632 ( .A(n15455), .B(n15454), .Z(n15456) );
  NAND U15633 ( .A(b[0]), .B(a[118]), .Z(n15329) );
  XNOR U15634 ( .A(b[1]), .B(n15329), .Z(n15331) );
  NANDN U15635 ( .A(b[0]), .B(a[117]), .Z(n15330) );
  NAND U15636 ( .A(n15331), .B(n15330), .Z(n15403) );
  NANDN U15637 ( .A(n19394), .B(n15332), .Z(n15334) );
  XOR U15638 ( .A(b[29]), .B(a[90]), .Z(n15481) );
  NANDN U15639 ( .A(n19395), .B(n15481), .Z(n15333) );
  AND U15640 ( .A(n15334), .B(n15333), .Z(n15401) );
  AND U15641 ( .A(b[31]), .B(a[86]), .Z(n15400) );
  XNOR U15642 ( .A(n15401), .B(n15400), .Z(n15402) );
  XNOR U15643 ( .A(n15403), .B(n15402), .Z(n15442) );
  NANDN U15644 ( .A(n19005), .B(n15335), .Z(n15337) );
  XOR U15645 ( .A(b[23]), .B(a[96]), .Z(n15484) );
  NANDN U15646 ( .A(n19055), .B(n15484), .Z(n15336) );
  AND U15647 ( .A(n15337), .B(n15336), .Z(n15475) );
  NANDN U15648 ( .A(n17362), .B(n15338), .Z(n15340) );
  XOR U15649 ( .A(a[112]), .B(b[7]), .Z(n15487) );
  NANDN U15650 ( .A(n17522), .B(n15487), .Z(n15339) );
  AND U15651 ( .A(n15340), .B(n15339), .Z(n15473) );
  NANDN U15652 ( .A(n19116), .B(n15341), .Z(n15343) );
  XOR U15653 ( .A(b[25]), .B(a[94]), .Z(n15490) );
  NANDN U15654 ( .A(n19179), .B(n15490), .Z(n15342) );
  NAND U15655 ( .A(n15343), .B(n15342), .Z(n15472) );
  XNOR U15656 ( .A(n15473), .B(n15472), .Z(n15474) );
  XOR U15657 ( .A(n15475), .B(n15474), .Z(n15443) );
  XNOR U15658 ( .A(n15442), .B(n15443), .Z(n15444) );
  NANDN U15659 ( .A(n18113), .B(n15344), .Z(n15346) );
  XOR U15660 ( .A(b[13]), .B(a[106]), .Z(n15493) );
  NANDN U15661 ( .A(n18229), .B(n15493), .Z(n15345) );
  AND U15662 ( .A(n15346), .B(n15345), .Z(n15437) );
  NANDN U15663 ( .A(n17888), .B(n15347), .Z(n15349) );
  XOR U15664 ( .A(b[11]), .B(a[108]), .Z(n15496) );
  NANDN U15665 ( .A(n18025), .B(n15496), .Z(n15348) );
  NAND U15666 ( .A(n15349), .B(n15348), .Z(n15436) );
  XNOR U15667 ( .A(n15437), .B(n15436), .Z(n15438) );
  NANDN U15668 ( .A(n18487), .B(n15350), .Z(n15352) );
  XOR U15669 ( .A(b[15]), .B(a[104]), .Z(n15499) );
  NANDN U15670 ( .A(n18311), .B(n15499), .Z(n15351) );
  AND U15671 ( .A(n15352), .B(n15351), .Z(n15433) );
  NANDN U15672 ( .A(n18853), .B(n15353), .Z(n15355) );
  XOR U15673 ( .A(b[21]), .B(a[98]), .Z(n15502) );
  NANDN U15674 ( .A(n18926), .B(n15502), .Z(n15354) );
  AND U15675 ( .A(n15355), .B(n15354), .Z(n15431) );
  NANDN U15676 ( .A(n17613), .B(n15356), .Z(n15358) );
  XOR U15677 ( .A(a[110]), .B(b[9]), .Z(n15505) );
  NANDN U15678 ( .A(n17739), .B(n15505), .Z(n15357) );
  NAND U15679 ( .A(n15358), .B(n15357), .Z(n15430) );
  XNOR U15680 ( .A(n15431), .B(n15430), .Z(n15432) );
  XOR U15681 ( .A(n15433), .B(n15432), .Z(n15439) );
  XOR U15682 ( .A(n15438), .B(n15439), .Z(n15445) );
  XOR U15683 ( .A(n15444), .B(n15445), .Z(n15457) );
  XNOR U15684 ( .A(n15456), .B(n15457), .Z(n15388) );
  XNOR U15685 ( .A(n15389), .B(n15388), .Z(n15390) );
  XOR U15686 ( .A(n15391), .B(n15390), .Z(n15509) );
  XNOR U15687 ( .A(n15508), .B(n15509), .Z(n15510) );
  XNOR U15688 ( .A(n15511), .B(n15510), .Z(n15384) );
  XOR U15689 ( .A(n15385), .B(n15384), .Z(n15377) );
  NANDN U15690 ( .A(n15360), .B(n15359), .Z(n15364) );
  NANDN U15691 ( .A(n15362), .B(n15361), .Z(n15363) );
  AND U15692 ( .A(n15364), .B(n15363), .Z(n15376) );
  XOR U15693 ( .A(n15377), .B(n15376), .Z(n15379) );
  XNOR U15694 ( .A(n15378), .B(n15379), .Z(n15370) );
  XNOR U15695 ( .A(n15371), .B(n15370), .Z(n15372) );
  XNOR U15696 ( .A(n15373), .B(n15372), .Z(n15514) );
  XNOR U15697 ( .A(sreg[214]), .B(n15514), .Z(n15516) );
  NANDN U15698 ( .A(sreg[213]), .B(n15365), .Z(n15369) );
  NAND U15699 ( .A(n15367), .B(n15366), .Z(n15368) );
  NAND U15700 ( .A(n15369), .B(n15368), .Z(n15515) );
  XNOR U15701 ( .A(n15516), .B(n15515), .Z(c[214]) );
  NANDN U15702 ( .A(n15371), .B(n15370), .Z(n15375) );
  NANDN U15703 ( .A(n15373), .B(n15372), .Z(n15374) );
  AND U15704 ( .A(n15375), .B(n15374), .Z(n15522) );
  NANDN U15705 ( .A(n15377), .B(n15376), .Z(n15381) );
  NANDN U15706 ( .A(n15379), .B(n15378), .Z(n15380) );
  AND U15707 ( .A(n15381), .B(n15380), .Z(n15520) );
  NANDN U15708 ( .A(n15383), .B(n15382), .Z(n15387) );
  NAND U15709 ( .A(n15385), .B(n15384), .Z(n15386) );
  AND U15710 ( .A(n15387), .B(n15386), .Z(n15527) );
  NANDN U15711 ( .A(n15389), .B(n15388), .Z(n15393) );
  NANDN U15712 ( .A(n15391), .B(n15390), .Z(n15392) );
  AND U15713 ( .A(n15393), .B(n15392), .Z(n15532) );
  NANDN U15714 ( .A(n15395), .B(n15394), .Z(n15399) );
  NAND U15715 ( .A(n15397), .B(n15396), .Z(n15398) );
  AND U15716 ( .A(n15399), .B(n15398), .Z(n15531) );
  XNOR U15717 ( .A(n15532), .B(n15531), .Z(n15534) );
  NANDN U15718 ( .A(n15401), .B(n15400), .Z(n15405) );
  NANDN U15719 ( .A(n15403), .B(n15402), .Z(n15404) );
  AND U15720 ( .A(n15405), .B(n15404), .Z(n15611) );
  NANDN U15721 ( .A(n19237), .B(n15406), .Z(n15408) );
  XOR U15722 ( .A(b[27]), .B(a[93]), .Z(n15555) );
  NANDN U15723 ( .A(n19277), .B(n15555), .Z(n15407) );
  AND U15724 ( .A(n15408), .B(n15407), .Z(n15618) );
  NANDN U15725 ( .A(n17072), .B(n15409), .Z(n15411) );
  XOR U15726 ( .A(a[115]), .B(b[5]), .Z(n15558) );
  NANDN U15727 ( .A(n17223), .B(n15558), .Z(n15410) );
  AND U15728 ( .A(n15411), .B(n15410), .Z(n15616) );
  NANDN U15729 ( .A(n18673), .B(n15412), .Z(n15414) );
  XOR U15730 ( .A(b[19]), .B(a[101]), .Z(n15561) );
  NANDN U15731 ( .A(n18758), .B(n15561), .Z(n15413) );
  NAND U15732 ( .A(n15414), .B(n15413), .Z(n15615) );
  XNOR U15733 ( .A(n15616), .B(n15615), .Z(n15617) );
  XNOR U15734 ( .A(n15618), .B(n15617), .Z(n15609) );
  NANDN U15735 ( .A(n19425), .B(n15415), .Z(n15417) );
  XOR U15736 ( .A(b[31]), .B(a[89]), .Z(n15564) );
  NANDN U15737 ( .A(n19426), .B(n15564), .Z(n15416) );
  AND U15738 ( .A(n15417), .B(n15416), .Z(n15576) );
  NANDN U15739 ( .A(n17067), .B(n15418), .Z(n15420) );
  XOR U15740 ( .A(a[117]), .B(b[3]), .Z(n15567) );
  NANDN U15741 ( .A(n17068), .B(n15567), .Z(n15419) );
  AND U15742 ( .A(n15420), .B(n15419), .Z(n15574) );
  NANDN U15743 ( .A(n18514), .B(n15421), .Z(n15423) );
  XOR U15744 ( .A(b[17]), .B(a[103]), .Z(n15570) );
  NANDN U15745 ( .A(n18585), .B(n15570), .Z(n15422) );
  NAND U15746 ( .A(n15423), .B(n15422), .Z(n15573) );
  XNOR U15747 ( .A(n15574), .B(n15573), .Z(n15575) );
  XOR U15748 ( .A(n15576), .B(n15575), .Z(n15610) );
  XOR U15749 ( .A(n15609), .B(n15610), .Z(n15612) );
  XOR U15750 ( .A(n15611), .B(n15612), .Z(n15544) );
  NANDN U15751 ( .A(n15425), .B(n15424), .Z(n15429) );
  NANDN U15752 ( .A(n15427), .B(n15426), .Z(n15428) );
  AND U15753 ( .A(n15429), .B(n15428), .Z(n15597) );
  NANDN U15754 ( .A(n15431), .B(n15430), .Z(n15435) );
  NANDN U15755 ( .A(n15433), .B(n15432), .Z(n15434) );
  NAND U15756 ( .A(n15435), .B(n15434), .Z(n15598) );
  XNOR U15757 ( .A(n15597), .B(n15598), .Z(n15599) );
  NANDN U15758 ( .A(n15437), .B(n15436), .Z(n15441) );
  NANDN U15759 ( .A(n15439), .B(n15438), .Z(n15440) );
  NAND U15760 ( .A(n15441), .B(n15440), .Z(n15600) );
  XNOR U15761 ( .A(n15599), .B(n15600), .Z(n15543) );
  XNOR U15762 ( .A(n15544), .B(n15543), .Z(n15546) );
  NANDN U15763 ( .A(n15443), .B(n15442), .Z(n15447) );
  NANDN U15764 ( .A(n15445), .B(n15444), .Z(n15446) );
  AND U15765 ( .A(n15447), .B(n15446), .Z(n15545) );
  XOR U15766 ( .A(n15546), .B(n15545), .Z(n15660) );
  NANDN U15767 ( .A(n15449), .B(n15448), .Z(n15453) );
  NANDN U15768 ( .A(n15451), .B(n15450), .Z(n15452) );
  AND U15769 ( .A(n15453), .B(n15452), .Z(n15657) );
  NANDN U15770 ( .A(n15455), .B(n15454), .Z(n15459) );
  NANDN U15771 ( .A(n15457), .B(n15456), .Z(n15458) );
  AND U15772 ( .A(n15459), .B(n15458), .Z(n15540) );
  NANDN U15773 ( .A(n15461), .B(n15460), .Z(n15465) );
  OR U15774 ( .A(n15463), .B(n15462), .Z(n15464) );
  AND U15775 ( .A(n15465), .B(n15464), .Z(n15538) );
  NANDN U15776 ( .A(n15467), .B(n15466), .Z(n15471) );
  NANDN U15777 ( .A(n15469), .B(n15468), .Z(n15470) );
  AND U15778 ( .A(n15471), .B(n15470), .Z(n15604) );
  NANDN U15779 ( .A(n15473), .B(n15472), .Z(n15477) );
  NANDN U15780 ( .A(n15475), .B(n15474), .Z(n15476) );
  NAND U15781 ( .A(n15477), .B(n15476), .Z(n15603) );
  XNOR U15782 ( .A(n15604), .B(n15603), .Z(n15605) );
  NAND U15783 ( .A(b[0]), .B(a[119]), .Z(n15478) );
  XNOR U15784 ( .A(b[1]), .B(n15478), .Z(n15480) );
  NANDN U15785 ( .A(b[0]), .B(a[118]), .Z(n15479) );
  NAND U15786 ( .A(n15480), .B(n15479), .Z(n15552) );
  NANDN U15787 ( .A(n19394), .B(n15481), .Z(n15483) );
  XOR U15788 ( .A(b[29]), .B(a[91]), .Z(n15630) );
  NANDN U15789 ( .A(n19395), .B(n15630), .Z(n15482) );
  AND U15790 ( .A(n15483), .B(n15482), .Z(n15550) );
  AND U15791 ( .A(b[31]), .B(a[87]), .Z(n15549) );
  XNOR U15792 ( .A(n15550), .B(n15549), .Z(n15551) );
  XNOR U15793 ( .A(n15552), .B(n15551), .Z(n15591) );
  NANDN U15794 ( .A(n19005), .B(n15484), .Z(n15486) );
  XOR U15795 ( .A(b[23]), .B(a[97]), .Z(n15633) );
  NANDN U15796 ( .A(n19055), .B(n15633), .Z(n15485) );
  AND U15797 ( .A(n15486), .B(n15485), .Z(n15624) );
  NANDN U15798 ( .A(n17362), .B(n15487), .Z(n15489) );
  XOR U15799 ( .A(a[113]), .B(b[7]), .Z(n15636) );
  NANDN U15800 ( .A(n17522), .B(n15636), .Z(n15488) );
  AND U15801 ( .A(n15489), .B(n15488), .Z(n15622) );
  NANDN U15802 ( .A(n19116), .B(n15490), .Z(n15492) );
  XOR U15803 ( .A(b[25]), .B(a[95]), .Z(n15639) );
  NANDN U15804 ( .A(n19179), .B(n15639), .Z(n15491) );
  NAND U15805 ( .A(n15492), .B(n15491), .Z(n15621) );
  XNOR U15806 ( .A(n15622), .B(n15621), .Z(n15623) );
  XOR U15807 ( .A(n15624), .B(n15623), .Z(n15592) );
  XNOR U15808 ( .A(n15591), .B(n15592), .Z(n15593) );
  NANDN U15809 ( .A(n18113), .B(n15493), .Z(n15495) );
  XOR U15810 ( .A(b[13]), .B(a[107]), .Z(n15642) );
  NANDN U15811 ( .A(n18229), .B(n15642), .Z(n15494) );
  AND U15812 ( .A(n15495), .B(n15494), .Z(n15586) );
  NANDN U15813 ( .A(n17888), .B(n15496), .Z(n15498) );
  XOR U15814 ( .A(b[11]), .B(a[109]), .Z(n15645) );
  NANDN U15815 ( .A(n18025), .B(n15645), .Z(n15497) );
  NAND U15816 ( .A(n15498), .B(n15497), .Z(n15585) );
  XNOR U15817 ( .A(n15586), .B(n15585), .Z(n15587) );
  NANDN U15818 ( .A(n18487), .B(n15499), .Z(n15501) );
  XOR U15819 ( .A(b[15]), .B(a[105]), .Z(n15648) );
  NANDN U15820 ( .A(n18311), .B(n15648), .Z(n15500) );
  AND U15821 ( .A(n15501), .B(n15500), .Z(n15582) );
  NANDN U15822 ( .A(n18853), .B(n15502), .Z(n15504) );
  XOR U15823 ( .A(b[21]), .B(a[99]), .Z(n15651) );
  NANDN U15824 ( .A(n18926), .B(n15651), .Z(n15503) );
  AND U15825 ( .A(n15504), .B(n15503), .Z(n15580) );
  NANDN U15826 ( .A(n17613), .B(n15505), .Z(n15507) );
  XOR U15827 ( .A(a[111]), .B(b[9]), .Z(n15654) );
  NANDN U15828 ( .A(n17739), .B(n15654), .Z(n15506) );
  NAND U15829 ( .A(n15507), .B(n15506), .Z(n15579) );
  XNOR U15830 ( .A(n15580), .B(n15579), .Z(n15581) );
  XOR U15831 ( .A(n15582), .B(n15581), .Z(n15588) );
  XOR U15832 ( .A(n15587), .B(n15588), .Z(n15594) );
  XOR U15833 ( .A(n15593), .B(n15594), .Z(n15606) );
  XNOR U15834 ( .A(n15605), .B(n15606), .Z(n15537) );
  XNOR U15835 ( .A(n15538), .B(n15537), .Z(n15539) );
  XOR U15836 ( .A(n15540), .B(n15539), .Z(n15658) );
  XNOR U15837 ( .A(n15657), .B(n15658), .Z(n15659) );
  XNOR U15838 ( .A(n15660), .B(n15659), .Z(n15533) );
  XOR U15839 ( .A(n15534), .B(n15533), .Z(n15526) );
  NANDN U15840 ( .A(n15509), .B(n15508), .Z(n15513) );
  NANDN U15841 ( .A(n15511), .B(n15510), .Z(n15512) );
  AND U15842 ( .A(n15513), .B(n15512), .Z(n15525) );
  XOR U15843 ( .A(n15526), .B(n15525), .Z(n15528) );
  XNOR U15844 ( .A(n15527), .B(n15528), .Z(n15519) );
  XNOR U15845 ( .A(n15520), .B(n15519), .Z(n15521) );
  XNOR U15846 ( .A(n15522), .B(n15521), .Z(n15663) );
  XNOR U15847 ( .A(sreg[215]), .B(n15663), .Z(n15665) );
  NANDN U15848 ( .A(sreg[214]), .B(n15514), .Z(n15518) );
  NAND U15849 ( .A(n15516), .B(n15515), .Z(n15517) );
  NAND U15850 ( .A(n15518), .B(n15517), .Z(n15664) );
  XNOR U15851 ( .A(n15665), .B(n15664), .Z(c[215]) );
  NANDN U15852 ( .A(n15520), .B(n15519), .Z(n15524) );
  NANDN U15853 ( .A(n15522), .B(n15521), .Z(n15523) );
  AND U15854 ( .A(n15524), .B(n15523), .Z(n15671) );
  NANDN U15855 ( .A(n15526), .B(n15525), .Z(n15530) );
  NANDN U15856 ( .A(n15528), .B(n15527), .Z(n15529) );
  AND U15857 ( .A(n15530), .B(n15529), .Z(n15669) );
  NANDN U15858 ( .A(n15532), .B(n15531), .Z(n15536) );
  NAND U15859 ( .A(n15534), .B(n15533), .Z(n15535) );
  AND U15860 ( .A(n15536), .B(n15535), .Z(n15676) );
  NANDN U15861 ( .A(n15538), .B(n15537), .Z(n15542) );
  NANDN U15862 ( .A(n15540), .B(n15539), .Z(n15541) );
  AND U15863 ( .A(n15542), .B(n15541), .Z(n15681) );
  NANDN U15864 ( .A(n15544), .B(n15543), .Z(n15548) );
  NAND U15865 ( .A(n15546), .B(n15545), .Z(n15547) );
  AND U15866 ( .A(n15548), .B(n15547), .Z(n15680) );
  XNOR U15867 ( .A(n15681), .B(n15680), .Z(n15683) );
  NANDN U15868 ( .A(n15550), .B(n15549), .Z(n15554) );
  NANDN U15869 ( .A(n15552), .B(n15551), .Z(n15553) );
  AND U15870 ( .A(n15554), .B(n15553), .Z(n15760) );
  NANDN U15871 ( .A(n19237), .B(n15555), .Z(n15557) );
  XOR U15872 ( .A(b[27]), .B(a[94]), .Z(n15704) );
  NANDN U15873 ( .A(n19277), .B(n15704), .Z(n15556) );
  AND U15874 ( .A(n15557), .B(n15556), .Z(n15767) );
  NANDN U15875 ( .A(n17072), .B(n15558), .Z(n15560) );
  XOR U15876 ( .A(a[116]), .B(b[5]), .Z(n15707) );
  NANDN U15877 ( .A(n17223), .B(n15707), .Z(n15559) );
  AND U15878 ( .A(n15560), .B(n15559), .Z(n15765) );
  NANDN U15879 ( .A(n18673), .B(n15561), .Z(n15563) );
  XOR U15880 ( .A(b[19]), .B(a[102]), .Z(n15710) );
  NANDN U15881 ( .A(n18758), .B(n15710), .Z(n15562) );
  NAND U15882 ( .A(n15563), .B(n15562), .Z(n15764) );
  XNOR U15883 ( .A(n15765), .B(n15764), .Z(n15766) );
  XNOR U15884 ( .A(n15767), .B(n15766), .Z(n15758) );
  NANDN U15885 ( .A(n19425), .B(n15564), .Z(n15566) );
  XOR U15886 ( .A(b[31]), .B(a[90]), .Z(n15713) );
  NANDN U15887 ( .A(n19426), .B(n15713), .Z(n15565) );
  AND U15888 ( .A(n15566), .B(n15565), .Z(n15725) );
  NANDN U15889 ( .A(n17067), .B(n15567), .Z(n15569) );
  XOR U15890 ( .A(a[118]), .B(b[3]), .Z(n15716) );
  NANDN U15891 ( .A(n17068), .B(n15716), .Z(n15568) );
  AND U15892 ( .A(n15569), .B(n15568), .Z(n15723) );
  NANDN U15893 ( .A(n18514), .B(n15570), .Z(n15572) );
  XOR U15894 ( .A(b[17]), .B(a[104]), .Z(n15719) );
  NANDN U15895 ( .A(n18585), .B(n15719), .Z(n15571) );
  NAND U15896 ( .A(n15572), .B(n15571), .Z(n15722) );
  XNOR U15897 ( .A(n15723), .B(n15722), .Z(n15724) );
  XOR U15898 ( .A(n15725), .B(n15724), .Z(n15759) );
  XOR U15899 ( .A(n15758), .B(n15759), .Z(n15761) );
  XOR U15900 ( .A(n15760), .B(n15761), .Z(n15693) );
  NANDN U15901 ( .A(n15574), .B(n15573), .Z(n15578) );
  NANDN U15902 ( .A(n15576), .B(n15575), .Z(n15577) );
  AND U15903 ( .A(n15578), .B(n15577), .Z(n15746) );
  NANDN U15904 ( .A(n15580), .B(n15579), .Z(n15584) );
  NANDN U15905 ( .A(n15582), .B(n15581), .Z(n15583) );
  NAND U15906 ( .A(n15584), .B(n15583), .Z(n15747) );
  XNOR U15907 ( .A(n15746), .B(n15747), .Z(n15748) );
  NANDN U15908 ( .A(n15586), .B(n15585), .Z(n15590) );
  NANDN U15909 ( .A(n15588), .B(n15587), .Z(n15589) );
  NAND U15910 ( .A(n15590), .B(n15589), .Z(n15749) );
  XNOR U15911 ( .A(n15748), .B(n15749), .Z(n15692) );
  XNOR U15912 ( .A(n15693), .B(n15692), .Z(n15695) );
  NANDN U15913 ( .A(n15592), .B(n15591), .Z(n15596) );
  NANDN U15914 ( .A(n15594), .B(n15593), .Z(n15595) );
  AND U15915 ( .A(n15596), .B(n15595), .Z(n15694) );
  XOR U15916 ( .A(n15695), .B(n15694), .Z(n15809) );
  NANDN U15917 ( .A(n15598), .B(n15597), .Z(n15602) );
  NANDN U15918 ( .A(n15600), .B(n15599), .Z(n15601) );
  AND U15919 ( .A(n15602), .B(n15601), .Z(n15806) );
  NANDN U15920 ( .A(n15604), .B(n15603), .Z(n15608) );
  NANDN U15921 ( .A(n15606), .B(n15605), .Z(n15607) );
  AND U15922 ( .A(n15608), .B(n15607), .Z(n15689) );
  NANDN U15923 ( .A(n15610), .B(n15609), .Z(n15614) );
  OR U15924 ( .A(n15612), .B(n15611), .Z(n15613) );
  AND U15925 ( .A(n15614), .B(n15613), .Z(n15687) );
  NANDN U15926 ( .A(n15616), .B(n15615), .Z(n15620) );
  NANDN U15927 ( .A(n15618), .B(n15617), .Z(n15619) );
  AND U15928 ( .A(n15620), .B(n15619), .Z(n15753) );
  NANDN U15929 ( .A(n15622), .B(n15621), .Z(n15626) );
  NANDN U15930 ( .A(n15624), .B(n15623), .Z(n15625) );
  NAND U15931 ( .A(n15626), .B(n15625), .Z(n15752) );
  XNOR U15932 ( .A(n15753), .B(n15752), .Z(n15754) );
  NAND U15933 ( .A(b[0]), .B(a[120]), .Z(n15627) );
  XNOR U15934 ( .A(b[1]), .B(n15627), .Z(n15629) );
  NANDN U15935 ( .A(b[0]), .B(a[119]), .Z(n15628) );
  NAND U15936 ( .A(n15629), .B(n15628), .Z(n15701) );
  NANDN U15937 ( .A(n19394), .B(n15630), .Z(n15632) );
  XOR U15938 ( .A(b[29]), .B(a[92]), .Z(n15779) );
  NANDN U15939 ( .A(n19395), .B(n15779), .Z(n15631) );
  AND U15940 ( .A(n15632), .B(n15631), .Z(n15699) );
  AND U15941 ( .A(b[31]), .B(a[88]), .Z(n15698) );
  XNOR U15942 ( .A(n15699), .B(n15698), .Z(n15700) );
  XNOR U15943 ( .A(n15701), .B(n15700), .Z(n15740) );
  NANDN U15944 ( .A(n19005), .B(n15633), .Z(n15635) );
  XOR U15945 ( .A(b[23]), .B(a[98]), .Z(n15782) );
  NANDN U15946 ( .A(n19055), .B(n15782), .Z(n15634) );
  AND U15947 ( .A(n15635), .B(n15634), .Z(n15773) );
  NANDN U15948 ( .A(n17362), .B(n15636), .Z(n15638) );
  XOR U15949 ( .A(a[114]), .B(b[7]), .Z(n15785) );
  NANDN U15950 ( .A(n17522), .B(n15785), .Z(n15637) );
  AND U15951 ( .A(n15638), .B(n15637), .Z(n15771) );
  NANDN U15952 ( .A(n19116), .B(n15639), .Z(n15641) );
  XOR U15953 ( .A(b[25]), .B(a[96]), .Z(n15788) );
  NANDN U15954 ( .A(n19179), .B(n15788), .Z(n15640) );
  NAND U15955 ( .A(n15641), .B(n15640), .Z(n15770) );
  XNOR U15956 ( .A(n15771), .B(n15770), .Z(n15772) );
  XOR U15957 ( .A(n15773), .B(n15772), .Z(n15741) );
  XNOR U15958 ( .A(n15740), .B(n15741), .Z(n15742) );
  NANDN U15959 ( .A(n18113), .B(n15642), .Z(n15644) );
  XOR U15960 ( .A(b[13]), .B(a[108]), .Z(n15791) );
  NANDN U15961 ( .A(n18229), .B(n15791), .Z(n15643) );
  AND U15962 ( .A(n15644), .B(n15643), .Z(n15735) );
  NANDN U15963 ( .A(n17888), .B(n15645), .Z(n15647) );
  XOR U15964 ( .A(a[110]), .B(b[11]), .Z(n15794) );
  NANDN U15965 ( .A(n18025), .B(n15794), .Z(n15646) );
  NAND U15966 ( .A(n15647), .B(n15646), .Z(n15734) );
  XNOR U15967 ( .A(n15735), .B(n15734), .Z(n15736) );
  NANDN U15968 ( .A(n18487), .B(n15648), .Z(n15650) );
  XOR U15969 ( .A(b[15]), .B(a[106]), .Z(n15797) );
  NANDN U15970 ( .A(n18311), .B(n15797), .Z(n15649) );
  AND U15971 ( .A(n15650), .B(n15649), .Z(n15731) );
  NANDN U15972 ( .A(n18853), .B(n15651), .Z(n15653) );
  XOR U15973 ( .A(b[21]), .B(a[100]), .Z(n15800) );
  NANDN U15974 ( .A(n18926), .B(n15800), .Z(n15652) );
  AND U15975 ( .A(n15653), .B(n15652), .Z(n15729) );
  NANDN U15976 ( .A(n17613), .B(n15654), .Z(n15656) );
  XOR U15977 ( .A(a[112]), .B(b[9]), .Z(n15803) );
  NANDN U15978 ( .A(n17739), .B(n15803), .Z(n15655) );
  NAND U15979 ( .A(n15656), .B(n15655), .Z(n15728) );
  XNOR U15980 ( .A(n15729), .B(n15728), .Z(n15730) );
  XOR U15981 ( .A(n15731), .B(n15730), .Z(n15737) );
  XOR U15982 ( .A(n15736), .B(n15737), .Z(n15743) );
  XOR U15983 ( .A(n15742), .B(n15743), .Z(n15755) );
  XNOR U15984 ( .A(n15754), .B(n15755), .Z(n15686) );
  XNOR U15985 ( .A(n15687), .B(n15686), .Z(n15688) );
  XOR U15986 ( .A(n15689), .B(n15688), .Z(n15807) );
  XNOR U15987 ( .A(n15806), .B(n15807), .Z(n15808) );
  XNOR U15988 ( .A(n15809), .B(n15808), .Z(n15682) );
  XOR U15989 ( .A(n15683), .B(n15682), .Z(n15675) );
  NANDN U15990 ( .A(n15658), .B(n15657), .Z(n15662) );
  NANDN U15991 ( .A(n15660), .B(n15659), .Z(n15661) );
  AND U15992 ( .A(n15662), .B(n15661), .Z(n15674) );
  XOR U15993 ( .A(n15675), .B(n15674), .Z(n15677) );
  XNOR U15994 ( .A(n15676), .B(n15677), .Z(n15668) );
  XNOR U15995 ( .A(n15669), .B(n15668), .Z(n15670) );
  XNOR U15996 ( .A(n15671), .B(n15670), .Z(n15812) );
  XNOR U15997 ( .A(sreg[216]), .B(n15812), .Z(n15814) );
  NANDN U15998 ( .A(sreg[215]), .B(n15663), .Z(n15667) );
  NAND U15999 ( .A(n15665), .B(n15664), .Z(n15666) );
  NAND U16000 ( .A(n15667), .B(n15666), .Z(n15813) );
  XNOR U16001 ( .A(n15814), .B(n15813), .Z(c[216]) );
  NANDN U16002 ( .A(n15669), .B(n15668), .Z(n15673) );
  NANDN U16003 ( .A(n15671), .B(n15670), .Z(n15672) );
  AND U16004 ( .A(n15673), .B(n15672), .Z(n15820) );
  NANDN U16005 ( .A(n15675), .B(n15674), .Z(n15679) );
  NANDN U16006 ( .A(n15677), .B(n15676), .Z(n15678) );
  AND U16007 ( .A(n15679), .B(n15678), .Z(n15818) );
  NANDN U16008 ( .A(n15681), .B(n15680), .Z(n15685) );
  NAND U16009 ( .A(n15683), .B(n15682), .Z(n15684) );
  AND U16010 ( .A(n15685), .B(n15684), .Z(n15825) );
  NANDN U16011 ( .A(n15687), .B(n15686), .Z(n15691) );
  NANDN U16012 ( .A(n15689), .B(n15688), .Z(n15690) );
  AND U16013 ( .A(n15691), .B(n15690), .Z(n15830) );
  NANDN U16014 ( .A(n15693), .B(n15692), .Z(n15697) );
  NAND U16015 ( .A(n15695), .B(n15694), .Z(n15696) );
  AND U16016 ( .A(n15697), .B(n15696), .Z(n15829) );
  XNOR U16017 ( .A(n15830), .B(n15829), .Z(n15832) );
  NANDN U16018 ( .A(n15699), .B(n15698), .Z(n15703) );
  NANDN U16019 ( .A(n15701), .B(n15700), .Z(n15702) );
  AND U16020 ( .A(n15703), .B(n15702), .Z(n15909) );
  NANDN U16021 ( .A(n19237), .B(n15704), .Z(n15706) );
  XOR U16022 ( .A(b[27]), .B(a[95]), .Z(n15853) );
  NANDN U16023 ( .A(n19277), .B(n15853), .Z(n15705) );
  AND U16024 ( .A(n15706), .B(n15705), .Z(n15916) );
  NANDN U16025 ( .A(n17072), .B(n15707), .Z(n15709) );
  XOR U16026 ( .A(a[117]), .B(b[5]), .Z(n15856) );
  NANDN U16027 ( .A(n17223), .B(n15856), .Z(n15708) );
  AND U16028 ( .A(n15709), .B(n15708), .Z(n15914) );
  NANDN U16029 ( .A(n18673), .B(n15710), .Z(n15712) );
  XOR U16030 ( .A(b[19]), .B(a[103]), .Z(n15859) );
  NANDN U16031 ( .A(n18758), .B(n15859), .Z(n15711) );
  NAND U16032 ( .A(n15712), .B(n15711), .Z(n15913) );
  XNOR U16033 ( .A(n15914), .B(n15913), .Z(n15915) );
  XNOR U16034 ( .A(n15916), .B(n15915), .Z(n15907) );
  NANDN U16035 ( .A(n19425), .B(n15713), .Z(n15715) );
  XOR U16036 ( .A(b[31]), .B(a[91]), .Z(n15862) );
  NANDN U16037 ( .A(n19426), .B(n15862), .Z(n15714) );
  AND U16038 ( .A(n15715), .B(n15714), .Z(n15874) );
  NANDN U16039 ( .A(n17067), .B(n15716), .Z(n15718) );
  XOR U16040 ( .A(a[119]), .B(b[3]), .Z(n15865) );
  NANDN U16041 ( .A(n17068), .B(n15865), .Z(n15717) );
  AND U16042 ( .A(n15718), .B(n15717), .Z(n15872) );
  NANDN U16043 ( .A(n18514), .B(n15719), .Z(n15721) );
  XOR U16044 ( .A(b[17]), .B(a[105]), .Z(n15868) );
  NANDN U16045 ( .A(n18585), .B(n15868), .Z(n15720) );
  NAND U16046 ( .A(n15721), .B(n15720), .Z(n15871) );
  XNOR U16047 ( .A(n15872), .B(n15871), .Z(n15873) );
  XOR U16048 ( .A(n15874), .B(n15873), .Z(n15908) );
  XOR U16049 ( .A(n15907), .B(n15908), .Z(n15910) );
  XOR U16050 ( .A(n15909), .B(n15910), .Z(n15842) );
  NANDN U16051 ( .A(n15723), .B(n15722), .Z(n15727) );
  NANDN U16052 ( .A(n15725), .B(n15724), .Z(n15726) );
  AND U16053 ( .A(n15727), .B(n15726), .Z(n15895) );
  NANDN U16054 ( .A(n15729), .B(n15728), .Z(n15733) );
  NANDN U16055 ( .A(n15731), .B(n15730), .Z(n15732) );
  NAND U16056 ( .A(n15733), .B(n15732), .Z(n15896) );
  XNOR U16057 ( .A(n15895), .B(n15896), .Z(n15897) );
  NANDN U16058 ( .A(n15735), .B(n15734), .Z(n15739) );
  NANDN U16059 ( .A(n15737), .B(n15736), .Z(n15738) );
  NAND U16060 ( .A(n15739), .B(n15738), .Z(n15898) );
  XNOR U16061 ( .A(n15897), .B(n15898), .Z(n15841) );
  XNOR U16062 ( .A(n15842), .B(n15841), .Z(n15844) );
  NANDN U16063 ( .A(n15741), .B(n15740), .Z(n15745) );
  NANDN U16064 ( .A(n15743), .B(n15742), .Z(n15744) );
  AND U16065 ( .A(n15745), .B(n15744), .Z(n15843) );
  XOR U16066 ( .A(n15844), .B(n15843), .Z(n15958) );
  NANDN U16067 ( .A(n15747), .B(n15746), .Z(n15751) );
  NANDN U16068 ( .A(n15749), .B(n15748), .Z(n15750) );
  AND U16069 ( .A(n15751), .B(n15750), .Z(n15955) );
  NANDN U16070 ( .A(n15753), .B(n15752), .Z(n15757) );
  NANDN U16071 ( .A(n15755), .B(n15754), .Z(n15756) );
  AND U16072 ( .A(n15757), .B(n15756), .Z(n15838) );
  NANDN U16073 ( .A(n15759), .B(n15758), .Z(n15763) );
  OR U16074 ( .A(n15761), .B(n15760), .Z(n15762) );
  AND U16075 ( .A(n15763), .B(n15762), .Z(n15836) );
  NANDN U16076 ( .A(n15765), .B(n15764), .Z(n15769) );
  NANDN U16077 ( .A(n15767), .B(n15766), .Z(n15768) );
  AND U16078 ( .A(n15769), .B(n15768), .Z(n15902) );
  NANDN U16079 ( .A(n15771), .B(n15770), .Z(n15775) );
  NANDN U16080 ( .A(n15773), .B(n15772), .Z(n15774) );
  NAND U16081 ( .A(n15775), .B(n15774), .Z(n15901) );
  XNOR U16082 ( .A(n15902), .B(n15901), .Z(n15903) );
  AND U16083 ( .A(a[121]), .B(b[0]), .Z(n15776) );
  XOR U16084 ( .A(b[1]), .B(n15776), .Z(n15778) );
  NANDN U16085 ( .A(b[0]), .B(a[120]), .Z(n15777) );
  AND U16086 ( .A(n15778), .B(n15777), .Z(n15849) );
  NANDN U16087 ( .A(n19394), .B(n15779), .Z(n15781) );
  XOR U16088 ( .A(b[29]), .B(a[93]), .Z(n15928) );
  NANDN U16089 ( .A(n19395), .B(n15928), .Z(n15780) );
  AND U16090 ( .A(n15781), .B(n15780), .Z(n15848) );
  AND U16091 ( .A(b[31]), .B(a[89]), .Z(n15847) );
  XOR U16092 ( .A(n15848), .B(n15847), .Z(n15850) );
  XNOR U16093 ( .A(n15849), .B(n15850), .Z(n15889) );
  NANDN U16094 ( .A(n19005), .B(n15782), .Z(n15784) );
  XOR U16095 ( .A(b[23]), .B(a[99]), .Z(n15931) );
  NANDN U16096 ( .A(n19055), .B(n15931), .Z(n15783) );
  AND U16097 ( .A(n15784), .B(n15783), .Z(n15922) );
  NANDN U16098 ( .A(n17362), .B(n15785), .Z(n15787) );
  XOR U16099 ( .A(a[115]), .B(b[7]), .Z(n15934) );
  NANDN U16100 ( .A(n17522), .B(n15934), .Z(n15786) );
  AND U16101 ( .A(n15787), .B(n15786), .Z(n15920) );
  NANDN U16102 ( .A(n19116), .B(n15788), .Z(n15790) );
  XOR U16103 ( .A(b[25]), .B(a[97]), .Z(n15937) );
  NANDN U16104 ( .A(n19179), .B(n15937), .Z(n15789) );
  NAND U16105 ( .A(n15790), .B(n15789), .Z(n15919) );
  XNOR U16106 ( .A(n15920), .B(n15919), .Z(n15921) );
  XOR U16107 ( .A(n15922), .B(n15921), .Z(n15890) );
  XNOR U16108 ( .A(n15889), .B(n15890), .Z(n15891) );
  NANDN U16109 ( .A(n18113), .B(n15791), .Z(n15793) );
  XOR U16110 ( .A(b[13]), .B(a[109]), .Z(n15940) );
  NANDN U16111 ( .A(n18229), .B(n15940), .Z(n15792) );
  AND U16112 ( .A(n15793), .B(n15792), .Z(n15884) );
  NANDN U16113 ( .A(n17888), .B(n15794), .Z(n15796) );
  XOR U16114 ( .A(a[111]), .B(b[11]), .Z(n15943) );
  NANDN U16115 ( .A(n18025), .B(n15943), .Z(n15795) );
  NAND U16116 ( .A(n15796), .B(n15795), .Z(n15883) );
  XNOR U16117 ( .A(n15884), .B(n15883), .Z(n15885) );
  NANDN U16118 ( .A(n18487), .B(n15797), .Z(n15799) );
  XOR U16119 ( .A(b[15]), .B(a[107]), .Z(n15946) );
  NANDN U16120 ( .A(n18311), .B(n15946), .Z(n15798) );
  AND U16121 ( .A(n15799), .B(n15798), .Z(n15880) );
  NANDN U16122 ( .A(n18853), .B(n15800), .Z(n15802) );
  XOR U16123 ( .A(b[21]), .B(a[101]), .Z(n15949) );
  NANDN U16124 ( .A(n18926), .B(n15949), .Z(n15801) );
  AND U16125 ( .A(n15802), .B(n15801), .Z(n15878) );
  NANDN U16126 ( .A(n17613), .B(n15803), .Z(n15805) );
  XOR U16127 ( .A(a[113]), .B(b[9]), .Z(n15952) );
  NANDN U16128 ( .A(n17739), .B(n15952), .Z(n15804) );
  NAND U16129 ( .A(n15805), .B(n15804), .Z(n15877) );
  XNOR U16130 ( .A(n15878), .B(n15877), .Z(n15879) );
  XOR U16131 ( .A(n15880), .B(n15879), .Z(n15886) );
  XOR U16132 ( .A(n15885), .B(n15886), .Z(n15892) );
  XOR U16133 ( .A(n15891), .B(n15892), .Z(n15904) );
  XNOR U16134 ( .A(n15903), .B(n15904), .Z(n15835) );
  XNOR U16135 ( .A(n15836), .B(n15835), .Z(n15837) );
  XOR U16136 ( .A(n15838), .B(n15837), .Z(n15956) );
  XNOR U16137 ( .A(n15955), .B(n15956), .Z(n15957) );
  XNOR U16138 ( .A(n15958), .B(n15957), .Z(n15831) );
  XOR U16139 ( .A(n15832), .B(n15831), .Z(n15824) );
  NANDN U16140 ( .A(n15807), .B(n15806), .Z(n15811) );
  NANDN U16141 ( .A(n15809), .B(n15808), .Z(n15810) );
  AND U16142 ( .A(n15811), .B(n15810), .Z(n15823) );
  XOR U16143 ( .A(n15824), .B(n15823), .Z(n15826) );
  XNOR U16144 ( .A(n15825), .B(n15826), .Z(n15817) );
  XNOR U16145 ( .A(n15818), .B(n15817), .Z(n15819) );
  XNOR U16146 ( .A(n15820), .B(n15819), .Z(n15961) );
  XNOR U16147 ( .A(sreg[217]), .B(n15961), .Z(n15963) );
  NANDN U16148 ( .A(sreg[216]), .B(n15812), .Z(n15816) );
  NAND U16149 ( .A(n15814), .B(n15813), .Z(n15815) );
  NAND U16150 ( .A(n15816), .B(n15815), .Z(n15962) );
  XNOR U16151 ( .A(n15963), .B(n15962), .Z(c[217]) );
  NANDN U16152 ( .A(n15818), .B(n15817), .Z(n15822) );
  NANDN U16153 ( .A(n15820), .B(n15819), .Z(n15821) );
  AND U16154 ( .A(n15822), .B(n15821), .Z(n15969) );
  NANDN U16155 ( .A(n15824), .B(n15823), .Z(n15828) );
  NANDN U16156 ( .A(n15826), .B(n15825), .Z(n15827) );
  AND U16157 ( .A(n15828), .B(n15827), .Z(n15967) );
  NANDN U16158 ( .A(n15830), .B(n15829), .Z(n15834) );
  NAND U16159 ( .A(n15832), .B(n15831), .Z(n15833) );
  AND U16160 ( .A(n15834), .B(n15833), .Z(n15974) );
  NANDN U16161 ( .A(n15836), .B(n15835), .Z(n15840) );
  NANDN U16162 ( .A(n15838), .B(n15837), .Z(n15839) );
  AND U16163 ( .A(n15840), .B(n15839), .Z(n15979) );
  NANDN U16164 ( .A(n15842), .B(n15841), .Z(n15846) );
  NAND U16165 ( .A(n15844), .B(n15843), .Z(n15845) );
  AND U16166 ( .A(n15846), .B(n15845), .Z(n15978) );
  XNOR U16167 ( .A(n15979), .B(n15978), .Z(n15981) );
  NANDN U16168 ( .A(n15848), .B(n15847), .Z(n15852) );
  NANDN U16169 ( .A(n15850), .B(n15849), .Z(n15851) );
  AND U16170 ( .A(n15852), .B(n15851), .Z(n16058) );
  NANDN U16171 ( .A(n19237), .B(n15853), .Z(n15855) );
  XOR U16172 ( .A(b[27]), .B(a[96]), .Z(n16002) );
  NANDN U16173 ( .A(n19277), .B(n16002), .Z(n15854) );
  AND U16174 ( .A(n15855), .B(n15854), .Z(n16065) );
  NANDN U16175 ( .A(n17072), .B(n15856), .Z(n15858) );
  XOR U16176 ( .A(a[118]), .B(b[5]), .Z(n16005) );
  NANDN U16177 ( .A(n17223), .B(n16005), .Z(n15857) );
  AND U16178 ( .A(n15858), .B(n15857), .Z(n16063) );
  NANDN U16179 ( .A(n18673), .B(n15859), .Z(n15861) );
  XOR U16180 ( .A(b[19]), .B(a[104]), .Z(n16008) );
  NANDN U16181 ( .A(n18758), .B(n16008), .Z(n15860) );
  NAND U16182 ( .A(n15861), .B(n15860), .Z(n16062) );
  XNOR U16183 ( .A(n16063), .B(n16062), .Z(n16064) );
  XNOR U16184 ( .A(n16065), .B(n16064), .Z(n16056) );
  NANDN U16185 ( .A(n19425), .B(n15862), .Z(n15864) );
  XOR U16186 ( .A(b[31]), .B(a[92]), .Z(n16011) );
  NANDN U16187 ( .A(n19426), .B(n16011), .Z(n15863) );
  AND U16188 ( .A(n15864), .B(n15863), .Z(n16023) );
  NANDN U16189 ( .A(n17067), .B(n15865), .Z(n15867) );
  XOR U16190 ( .A(a[120]), .B(b[3]), .Z(n16014) );
  NANDN U16191 ( .A(n17068), .B(n16014), .Z(n15866) );
  AND U16192 ( .A(n15867), .B(n15866), .Z(n16021) );
  NANDN U16193 ( .A(n18514), .B(n15868), .Z(n15870) );
  XOR U16194 ( .A(b[17]), .B(a[106]), .Z(n16017) );
  NANDN U16195 ( .A(n18585), .B(n16017), .Z(n15869) );
  NAND U16196 ( .A(n15870), .B(n15869), .Z(n16020) );
  XNOR U16197 ( .A(n16021), .B(n16020), .Z(n16022) );
  XOR U16198 ( .A(n16023), .B(n16022), .Z(n16057) );
  XOR U16199 ( .A(n16056), .B(n16057), .Z(n16059) );
  XOR U16200 ( .A(n16058), .B(n16059), .Z(n15991) );
  NANDN U16201 ( .A(n15872), .B(n15871), .Z(n15876) );
  NANDN U16202 ( .A(n15874), .B(n15873), .Z(n15875) );
  AND U16203 ( .A(n15876), .B(n15875), .Z(n16044) );
  NANDN U16204 ( .A(n15878), .B(n15877), .Z(n15882) );
  NANDN U16205 ( .A(n15880), .B(n15879), .Z(n15881) );
  NAND U16206 ( .A(n15882), .B(n15881), .Z(n16045) );
  XNOR U16207 ( .A(n16044), .B(n16045), .Z(n16046) );
  NANDN U16208 ( .A(n15884), .B(n15883), .Z(n15888) );
  NANDN U16209 ( .A(n15886), .B(n15885), .Z(n15887) );
  NAND U16210 ( .A(n15888), .B(n15887), .Z(n16047) );
  XNOR U16211 ( .A(n16046), .B(n16047), .Z(n15990) );
  XNOR U16212 ( .A(n15991), .B(n15990), .Z(n15993) );
  NANDN U16213 ( .A(n15890), .B(n15889), .Z(n15894) );
  NANDN U16214 ( .A(n15892), .B(n15891), .Z(n15893) );
  AND U16215 ( .A(n15894), .B(n15893), .Z(n15992) );
  XOR U16216 ( .A(n15993), .B(n15992), .Z(n16107) );
  NANDN U16217 ( .A(n15896), .B(n15895), .Z(n15900) );
  NANDN U16218 ( .A(n15898), .B(n15897), .Z(n15899) );
  AND U16219 ( .A(n15900), .B(n15899), .Z(n16104) );
  NANDN U16220 ( .A(n15902), .B(n15901), .Z(n15906) );
  NANDN U16221 ( .A(n15904), .B(n15903), .Z(n15905) );
  AND U16222 ( .A(n15906), .B(n15905), .Z(n15987) );
  NANDN U16223 ( .A(n15908), .B(n15907), .Z(n15912) );
  OR U16224 ( .A(n15910), .B(n15909), .Z(n15911) );
  AND U16225 ( .A(n15912), .B(n15911), .Z(n15985) );
  NANDN U16226 ( .A(n15914), .B(n15913), .Z(n15918) );
  NANDN U16227 ( .A(n15916), .B(n15915), .Z(n15917) );
  AND U16228 ( .A(n15918), .B(n15917), .Z(n16051) );
  NANDN U16229 ( .A(n15920), .B(n15919), .Z(n15924) );
  NANDN U16230 ( .A(n15922), .B(n15921), .Z(n15923) );
  NAND U16231 ( .A(n15924), .B(n15923), .Z(n16050) );
  XNOR U16232 ( .A(n16051), .B(n16050), .Z(n16052) );
  NAND U16233 ( .A(b[0]), .B(a[122]), .Z(n15925) );
  XNOR U16234 ( .A(b[1]), .B(n15925), .Z(n15927) );
  NANDN U16235 ( .A(b[0]), .B(a[121]), .Z(n15926) );
  NAND U16236 ( .A(n15927), .B(n15926), .Z(n15999) );
  NANDN U16237 ( .A(n19394), .B(n15928), .Z(n15930) );
  XOR U16238 ( .A(b[29]), .B(a[94]), .Z(n16077) );
  NANDN U16239 ( .A(n19395), .B(n16077), .Z(n15929) );
  AND U16240 ( .A(n15930), .B(n15929), .Z(n15997) );
  AND U16241 ( .A(b[31]), .B(a[90]), .Z(n15996) );
  XNOR U16242 ( .A(n15997), .B(n15996), .Z(n15998) );
  XNOR U16243 ( .A(n15999), .B(n15998), .Z(n16038) );
  NANDN U16244 ( .A(n19005), .B(n15931), .Z(n15933) );
  XOR U16245 ( .A(b[23]), .B(a[100]), .Z(n16080) );
  NANDN U16246 ( .A(n19055), .B(n16080), .Z(n15932) );
  AND U16247 ( .A(n15933), .B(n15932), .Z(n16071) );
  NANDN U16248 ( .A(n17362), .B(n15934), .Z(n15936) );
  XOR U16249 ( .A(a[116]), .B(b[7]), .Z(n16083) );
  NANDN U16250 ( .A(n17522), .B(n16083), .Z(n15935) );
  AND U16251 ( .A(n15936), .B(n15935), .Z(n16069) );
  NANDN U16252 ( .A(n19116), .B(n15937), .Z(n15939) );
  XOR U16253 ( .A(b[25]), .B(a[98]), .Z(n16086) );
  NANDN U16254 ( .A(n19179), .B(n16086), .Z(n15938) );
  NAND U16255 ( .A(n15939), .B(n15938), .Z(n16068) );
  XNOR U16256 ( .A(n16069), .B(n16068), .Z(n16070) );
  XOR U16257 ( .A(n16071), .B(n16070), .Z(n16039) );
  XNOR U16258 ( .A(n16038), .B(n16039), .Z(n16040) );
  NANDN U16259 ( .A(n18113), .B(n15940), .Z(n15942) );
  XOR U16260 ( .A(b[13]), .B(a[110]), .Z(n16089) );
  NANDN U16261 ( .A(n18229), .B(n16089), .Z(n15941) );
  AND U16262 ( .A(n15942), .B(n15941), .Z(n16033) );
  NANDN U16263 ( .A(n17888), .B(n15943), .Z(n15945) );
  XOR U16264 ( .A(a[112]), .B(b[11]), .Z(n16092) );
  NANDN U16265 ( .A(n18025), .B(n16092), .Z(n15944) );
  NAND U16266 ( .A(n15945), .B(n15944), .Z(n16032) );
  XNOR U16267 ( .A(n16033), .B(n16032), .Z(n16034) );
  NANDN U16268 ( .A(n18487), .B(n15946), .Z(n15948) );
  XOR U16269 ( .A(b[15]), .B(a[108]), .Z(n16095) );
  NANDN U16270 ( .A(n18311), .B(n16095), .Z(n15947) );
  AND U16271 ( .A(n15948), .B(n15947), .Z(n16029) );
  NANDN U16272 ( .A(n18853), .B(n15949), .Z(n15951) );
  XOR U16273 ( .A(b[21]), .B(a[102]), .Z(n16098) );
  NANDN U16274 ( .A(n18926), .B(n16098), .Z(n15950) );
  AND U16275 ( .A(n15951), .B(n15950), .Z(n16027) );
  NANDN U16276 ( .A(n17613), .B(n15952), .Z(n15954) );
  XOR U16277 ( .A(a[114]), .B(b[9]), .Z(n16101) );
  NANDN U16278 ( .A(n17739), .B(n16101), .Z(n15953) );
  NAND U16279 ( .A(n15954), .B(n15953), .Z(n16026) );
  XNOR U16280 ( .A(n16027), .B(n16026), .Z(n16028) );
  XOR U16281 ( .A(n16029), .B(n16028), .Z(n16035) );
  XOR U16282 ( .A(n16034), .B(n16035), .Z(n16041) );
  XOR U16283 ( .A(n16040), .B(n16041), .Z(n16053) );
  XNOR U16284 ( .A(n16052), .B(n16053), .Z(n15984) );
  XNOR U16285 ( .A(n15985), .B(n15984), .Z(n15986) );
  XOR U16286 ( .A(n15987), .B(n15986), .Z(n16105) );
  XNOR U16287 ( .A(n16104), .B(n16105), .Z(n16106) );
  XNOR U16288 ( .A(n16107), .B(n16106), .Z(n15980) );
  XOR U16289 ( .A(n15981), .B(n15980), .Z(n15973) );
  NANDN U16290 ( .A(n15956), .B(n15955), .Z(n15960) );
  NANDN U16291 ( .A(n15958), .B(n15957), .Z(n15959) );
  AND U16292 ( .A(n15960), .B(n15959), .Z(n15972) );
  XOR U16293 ( .A(n15973), .B(n15972), .Z(n15975) );
  XNOR U16294 ( .A(n15974), .B(n15975), .Z(n15966) );
  XNOR U16295 ( .A(n15967), .B(n15966), .Z(n15968) );
  XNOR U16296 ( .A(n15969), .B(n15968), .Z(n16110) );
  XNOR U16297 ( .A(sreg[218]), .B(n16110), .Z(n16112) );
  NANDN U16298 ( .A(sreg[217]), .B(n15961), .Z(n15965) );
  NAND U16299 ( .A(n15963), .B(n15962), .Z(n15964) );
  NAND U16300 ( .A(n15965), .B(n15964), .Z(n16111) );
  XNOR U16301 ( .A(n16112), .B(n16111), .Z(c[218]) );
  NANDN U16302 ( .A(n15967), .B(n15966), .Z(n15971) );
  NANDN U16303 ( .A(n15969), .B(n15968), .Z(n15970) );
  AND U16304 ( .A(n15971), .B(n15970), .Z(n16118) );
  NANDN U16305 ( .A(n15973), .B(n15972), .Z(n15977) );
  NANDN U16306 ( .A(n15975), .B(n15974), .Z(n15976) );
  AND U16307 ( .A(n15977), .B(n15976), .Z(n16116) );
  NANDN U16308 ( .A(n15979), .B(n15978), .Z(n15983) );
  NAND U16309 ( .A(n15981), .B(n15980), .Z(n15982) );
  AND U16310 ( .A(n15983), .B(n15982), .Z(n16123) );
  NANDN U16311 ( .A(n15985), .B(n15984), .Z(n15989) );
  NANDN U16312 ( .A(n15987), .B(n15986), .Z(n15988) );
  AND U16313 ( .A(n15989), .B(n15988), .Z(n16128) );
  NANDN U16314 ( .A(n15991), .B(n15990), .Z(n15995) );
  NAND U16315 ( .A(n15993), .B(n15992), .Z(n15994) );
  AND U16316 ( .A(n15995), .B(n15994), .Z(n16127) );
  XNOR U16317 ( .A(n16128), .B(n16127), .Z(n16130) );
  NANDN U16318 ( .A(n15997), .B(n15996), .Z(n16001) );
  NANDN U16319 ( .A(n15999), .B(n15998), .Z(n16000) );
  AND U16320 ( .A(n16001), .B(n16000), .Z(n16207) );
  NANDN U16321 ( .A(n19237), .B(n16002), .Z(n16004) );
  XOR U16322 ( .A(b[27]), .B(a[97]), .Z(n16151) );
  NANDN U16323 ( .A(n19277), .B(n16151), .Z(n16003) );
  AND U16324 ( .A(n16004), .B(n16003), .Z(n16214) );
  NANDN U16325 ( .A(n17072), .B(n16005), .Z(n16007) );
  XOR U16326 ( .A(a[119]), .B(b[5]), .Z(n16154) );
  NANDN U16327 ( .A(n17223), .B(n16154), .Z(n16006) );
  AND U16328 ( .A(n16007), .B(n16006), .Z(n16212) );
  NANDN U16329 ( .A(n18673), .B(n16008), .Z(n16010) );
  XOR U16330 ( .A(b[19]), .B(a[105]), .Z(n16157) );
  NANDN U16331 ( .A(n18758), .B(n16157), .Z(n16009) );
  NAND U16332 ( .A(n16010), .B(n16009), .Z(n16211) );
  XNOR U16333 ( .A(n16212), .B(n16211), .Z(n16213) );
  XNOR U16334 ( .A(n16214), .B(n16213), .Z(n16205) );
  NANDN U16335 ( .A(n19425), .B(n16011), .Z(n16013) );
  XOR U16336 ( .A(b[31]), .B(a[93]), .Z(n16160) );
  NANDN U16337 ( .A(n19426), .B(n16160), .Z(n16012) );
  AND U16338 ( .A(n16013), .B(n16012), .Z(n16172) );
  NANDN U16339 ( .A(n17067), .B(n16014), .Z(n16016) );
  XOR U16340 ( .A(a[121]), .B(b[3]), .Z(n16163) );
  NANDN U16341 ( .A(n17068), .B(n16163), .Z(n16015) );
  AND U16342 ( .A(n16016), .B(n16015), .Z(n16170) );
  NANDN U16343 ( .A(n18514), .B(n16017), .Z(n16019) );
  XOR U16344 ( .A(b[17]), .B(a[107]), .Z(n16166) );
  NANDN U16345 ( .A(n18585), .B(n16166), .Z(n16018) );
  NAND U16346 ( .A(n16019), .B(n16018), .Z(n16169) );
  XNOR U16347 ( .A(n16170), .B(n16169), .Z(n16171) );
  XOR U16348 ( .A(n16172), .B(n16171), .Z(n16206) );
  XOR U16349 ( .A(n16205), .B(n16206), .Z(n16208) );
  XOR U16350 ( .A(n16207), .B(n16208), .Z(n16140) );
  NANDN U16351 ( .A(n16021), .B(n16020), .Z(n16025) );
  NANDN U16352 ( .A(n16023), .B(n16022), .Z(n16024) );
  AND U16353 ( .A(n16025), .B(n16024), .Z(n16193) );
  NANDN U16354 ( .A(n16027), .B(n16026), .Z(n16031) );
  NANDN U16355 ( .A(n16029), .B(n16028), .Z(n16030) );
  NAND U16356 ( .A(n16031), .B(n16030), .Z(n16194) );
  XNOR U16357 ( .A(n16193), .B(n16194), .Z(n16195) );
  NANDN U16358 ( .A(n16033), .B(n16032), .Z(n16037) );
  NANDN U16359 ( .A(n16035), .B(n16034), .Z(n16036) );
  NAND U16360 ( .A(n16037), .B(n16036), .Z(n16196) );
  XNOR U16361 ( .A(n16195), .B(n16196), .Z(n16139) );
  XNOR U16362 ( .A(n16140), .B(n16139), .Z(n16142) );
  NANDN U16363 ( .A(n16039), .B(n16038), .Z(n16043) );
  NANDN U16364 ( .A(n16041), .B(n16040), .Z(n16042) );
  AND U16365 ( .A(n16043), .B(n16042), .Z(n16141) );
  XOR U16366 ( .A(n16142), .B(n16141), .Z(n16256) );
  NANDN U16367 ( .A(n16045), .B(n16044), .Z(n16049) );
  NANDN U16368 ( .A(n16047), .B(n16046), .Z(n16048) );
  AND U16369 ( .A(n16049), .B(n16048), .Z(n16253) );
  NANDN U16370 ( .A(n16051), .B(n16050), .Z(n16055) );
  NANDN U16371 ( .A(n16053), .B(n16052), .Z(n16054) );
  AND U16372 ( .A(n16055), .B(n16054), .Z(n16136) );
  NANDN U16373 ( .A(n16057), .B(n16056), .Z(n16061) );
  OR U16374 ( .A(n16059), .B(n16058), .Z(n16060) );
  AND U16375 ( .A(n16061), .B(n16060), .Z(n16134) );
  NANDN U16376 ( .A(n16063), .B(n16062), .Z(n16067) );
  NANDN U16377 ( .A(n16065), .B(n16064), .Z(n16066) );
  AND U16378 ( .A(n16067), .B(n16066), .Z(n16200) );
  NANDN U16379 ( .A(n16069), .B(n16068), .Z(n16073) );
  NANDN U16380 ( .A(n16071), .B(n16070), .Z(n16072) );
  NAND U16381 ( .A(n16073), .B(n16072), .Z(n16199) );
  XNOR U16382 ( .A(n16200), .B(n16199), .Z(n16201) );
  NAND U16383 ( .A(b[0]), .B(a[123]), .Z(n16074) );
  XNOR U16384 ( .A(b[1]), .B(n16074), .Z(n16076) );
  NANDN U16385 ( .A(b[0]), .B(a[122]), .Z(n16075) );
  NAND U16386 ( .A(n16076), .B(n16075), .Z(n16148) );
  NANDN U16387 ( .A(n19394), .B(n16077), .Z(n16079) );
  XOR U16388 ( .A(b[29]), .B(a[95]), .Z(n16223) );
  NANDN U16389 ( .A(n19395), .B(n16223), .Z(n16078) );
  AND U16390 ( .A(n16079), .B(n16078), .Z(n16146) );
  AND U16391 ( .A(b[31]), .B(a[91]), .Z(n16145) );
  XNOR U16392 ( .A(n16146), .B(n16145), .Z(n16147) );
  XNOR U16393 ( .A(n16148), .B(n16147), .Z(n16187) );
  NANDN U16394 ( .A(n19005), .B(n16080), .Z(n16082) );
  XOR U16395 ( .A(b[23]), .B(a[101]), .Z(n16229) );
  NANDN U16396 ( .A(n19055), .B(n16229), .Z(n16081) );
  AND U16397 ( .A(n16082), .B(n16081), .Z(n16220) );
  NANDN U16398 ( .A(n17362), .B(n16083), .Z(n16085) );
  XOR U16399 ( .A(a[117]), .B(b[7]), .Z(n16232) );
  NANDN U16400 ( .A(n17522), .B(n16232), .Z(n16084) );
  AND U16401 ( .A(n16085), .B(n16084), .Z(n16218) );
  NANDN U16402 ( .A(n19116), .B(n16086), .Z(n16088) );
  XOR U16403 ( .A(b[25]), .B(a[99]), .Z(n16235) );
  NANDN U16404 ( .A(n19179), .B(n16235), .Z(n16087) );
  NAND U16405 ( .A(n16088), .B(n16087), .Z(n16217) );
  XNOR U16406 ( .A(n16218), .B(n16217), .Z(n16219) );
  XOR U16407 ( .A(n16220), .B(n16219), .Z(n16188) );
  XNOR U16408 ( .A(n16187), .B(n16188), .Z(n16189) );
  NANDN U16409 ( .A(n18113), .B(n16089), .Z(n16091) );
  XOR U16410 ( .A(b[13]), .B(a[111]), .Z(n16238) );
  NANDN U16411 ( .A(n18229), .B(n16238), .Z(n16090) );
  AND U16412 ( .A(n16091), .B(n16090), .Z(n16182) );
  NANDN U16413 ( .A(n17888), .B(n16092), .Z(n16094) );
  XOR U16414 ( .A(a[113]), .B(b[11]), .Z(n16241) );
  NANDN U16415 ( .A(n18025), .B(n16241), .Z(n16093) );
  NAND U16416 ( .A(n16094), .B(n16093), .Z(n16181) );
  XNOR U16417 ( .A(n16182), .B(n16181), .Z(n16183) );
  NANDN U16418 ( .A(n18487), .B(n16095), .Z(n16097) );
  XOR U16419 ( .A(b[15]), .B(a[109]), .Z(n16244) );
  NANDN U16420 ( .A(n18311), .B(n16244), .Z(n16096) );
  AND U16421 ( .A(n16097), .B(n16096), .Z(n16178) );
  NANDN U16422 ( .A(n18853), .B(n16098), .Z(n16100) );
  XOR U16423 ( .A(b[21]), .B(a[103]), .Z(n16247) );
  NANDN U16424 ( .A(n18926), .B(n16247), .Z(n16099) );
  AND U16425 ( .A(n16100), .B(n16099), .Z(n16176) );
  NANDN U16426 ( .A(n17613), .B(n16101), .Z(n16103) );
  XOR U16427 ( .A(a[115]), .B(b[9]), .Z(n16250) );
  NANDN U16428 ( .A(n17739), .B(n16250), .Z(n16102) );
  NAND U16429 ( .A(n16103), .B(n16102), .Z(n16175) );
  XNOR U16430 ( .A(n16176), .B(n16175), .Z(n16177) );
  XOR U16431 ( .A(n16178), .B(n16177), .Z(n16184) );
  XOR U16432 ( .A(n16183), .B(n16184), .Z(n16190) );
  XOR U16433 ( .A(n16189), .B(n16190), .Z(n16202) );
  XNOR U16434 ( .A(n16201), .B(n16202), .Z(n16133) );
  XNOR U16435 ( .A(n16134), .B(n16133), .Z(n16135) );
  XOR U16436 ( .A(n16136), .B(n16135), .Z(n16254) );
  XNOR U16437 ( .A(n16253), .B(n16254), .Z(n16255) );
  XNOR U16438 ( .A(n16256), .B(n16255), .Z(n16129) );
  XOR U16439 ( .A(n16130), .B(n16129), .Z(n16122) );
  NANDN U16440 ( .A(n16105), .B(n16104), .Z(n16109) );
  NANDN U16441 ( .A(n16107), .B(n16106), .Z(n16108) );
  AND U16442 ( .A(n16109), .B(n16108), .Z(n16121) );
  XOR U16443 ( .A(n16122), .B(n16121), .Z(n16124) );
  XNOR U16444 ( .A(n16123), .B(n16124), .Z(n16115) );
  XNOR U16445 ( .A(n16116), .B(n16115), .Z(n16117) );
  XNOR U16446 ( .A(n16118), .B(n16117), .Z(n16259) );
  XNOR U16447 ( .A(sreg[219]), .B(n16259), .Z(n16261) );
  NANDN U16448 ( .A(sreg[218]), .B(n16110), .Z(n16114) );
  NAND U16449 ( .A(n16112), .B(n16111), .Z(n16113) );
  NAND U16450 ( .A(n16114), .B(n16113), .Z(n16260) );
  XNOR U16451 ( .A(n16261), .B(n16260), .Z(c[219]) );
  NANDN U16452 ( .A(n16116), .B(n16115), .Z(n16120) );
  NANDN U16453 ( .A(n16118), .B(n16117), .Z(n16119) );
  AND U16454 ( .A(n16120), .B(n16119), .Z(n16267) );
  NANDN U16455 ( .A(n16122), .B(n16121), .Z(n16126) );
  NANDN U16456 ( .A(n16124), .B(n16123), .Z(n16125) );
  AND U16457 ( .A(n16126), .B(n16125), .Z(n16265) );
  NANDN U16458 ( .A(n16128), .B(n16127), .Z(n16132) );
  NAND U16459 ( .A(n16130), .B(n16129), .Z(n16131) );
  AND U16460 ( .A(n16132), .B(n16131), .Z(n16402) );
  NANDN U16461 ( .A(n16134), .B(n16133), .Z(n16138) );
  NANDN U16462 ( .A(n16136), .B(n16135), .Z(n16137) );
  AND U16463 ( .A(n16138), .B(n16137), .Z(n16271) );
  NANDN U16464 ( .A(n16140), .B(n16139), .Z(n16144) );
  NAND U16465 ( .A(n16142), .B(n16141), .Z(n16143) );
  AND U16466 ( .A(n16144), .B(n16143), .Z(n16270) );
  XNOR U16467 ( .A(n16271), .B(n16270), .Z(n16273) );
  NANDN U16468 ( .A(n16146), .B(n16145), .Z(n16150) );
  NANDN U16469 ( .A(n16148), .B(n16147), .Z(n16149) );
  AND U16470 ( .A(n16150), .B(n16149), .Z(n16354) );
  NANDN U16471 ( .A(n19237), .B(n16151), .Z(n16153) );
  XOR U16472 ( .A(b[27]), .B(a[98]), .Z(n16300) );
  NANDN U16473 ( .A(n19277), .B(n16300), .Z(n16152) );
  AND U16474 ( .A(n16153), .B(n16152), .Z(n16397) );
  NANDN U16475 ( .A(n17072), .B(n16154), .Z(n16156) );
  XOR U16476 ( .A(a[120]), .B(b[5]), .Z(n16303) );
  NANDN U16477 ( .A(n17223), .B(n16303), .Z(n16155) );
  AND U16478 ( .A(n16156), .B(n16155), .Z(n16395) );
  NANDN U16479 ( .A(n18673), .B(n16157), .Z(n16159) );
  XOR U16480 ( .A(b[19]), .B(a[106]), .Z(n16306) );
  NANDN U16481 ( .A(n18758), .B(n16306), .Z(n16158) );
  NAND U16482 ( .A(n16159), .B(n16158), .Z(n16394) );
  XNOR U16483 ( .A(n16395), .B(n16394), .Z(n16396) );
  XNOR U16484 ( .A(n16397), .B(n16396), .Z(n16352) );
  NANDN U16485 ( .A(n19425), .B(n16160), .Z(n16162) );
  XOR U16486 ( .A(b[31]), .B(a[94]), .Z(n16309) );
  NANDN U16487 ( .A(n19426), .B(n16309), .Z(n16161) );
  AND U16488 ( .A(n16162), .B(n16161), .Z(n16321) );
  NANDN U16489 ( .A(n17067), .B(n16163), .Z(n16165) );
  XOR U16490 ( .A(a[122]), .B(b[3]), .Z(n16312) );
  NANDN U16491 ( .A(n17068), .B(n16312), .Z(n16164) );
  AND U16492 ( .A(n16165), .B(n16164), .Z(n16319) );
  NANDN U16493 ( .A(n18514), .B(n16166), .Z(n16168) );
  XOR U16494 ( .A(b[17]), .B(a[108]), .Z(n16315) );
  NANDN U16495 ( .A(n18585), .B(n16315), .Z(n16167) );
  NAND U16496 ( .A(n16168), .B(n16167), .Z(n16318) );
  XNOR U16497 ( .A(n16319), .B(n16318), .Z(n16320) );
  XOR U16498 ( .A(n16321), .B(n16320), .Z(n16353) );
  XOR U16499 ( .A(n16352), .B(n16353), .Z(n16355) );
  XOR U16500 ( .A(n16354), .B(n16355), .Z(n16289) );
  NANDN U16501 ( .A(n16170), .B(n16169), .Z(n16174) );
  NANDN U16502 ( .A(n16172), .B(n16171), .Z(n16173) );
  AND U16503 ( .A(n16174), .B(n16173), .Z(n16342) );
  NANDN U16504 ( .A(n16176), .B(n16175), .Z(n16180) );
  NANDN U16505 ( .A(n16178), .B(n16177), .Z(n16179) );
  NAND U16506 ( .A(n16180), .B(n16179), .Z(n16343) );
  XNOR U16507 ( .A(n16342), .B(n16343), .Z(n16344) );
  NANDN U16508 ( .A(n16182), .B(n16181), .Z(n16186) );
  NANDN U16509 ( .A(n16184), .B(n16183), .Z(n16185) );
  NAND U16510 ( .A(n16186), .B(n16185), .Z(n16345) );
  XNOR U16511 ( .A(n16344), .B(n16345), .Z(n16288) );
  XNOR U16512 ( .A(n16289), .B(n16288), .Z(n16291) );
  NANDN U16513 ( .A(n16188), .B(n16187), .Z(n16192) );
  NANDN U16514 ( .A(n16190), .B(n16189), .Z(n16191) );
  AND U16515 ( .A(n16192), .B(n16191), .Z(n16290) );
  XOR U16516 ( .A(n16291), .B(n16290), .Z(n16279) );
  NANDN U16517 ( .A(n16194), .B(n16193), .Z(n16198) );
  NANDN U16518 ( .A(n16196), .B(n16195), .Z(n16197) );
  AND U16519 ( .A(n16198), .B(n16197), .Z(n16276) );
  NANDN U16520 ( .A(n16200), .B(n16199), .Z(n16204) );
  NANDN U16521 ( .A(n16202), .B(n16201), .Z(n16203) );
  AND U16522 ( .A(n16204), .B(n16203), .Z(n16285) );
  NANDN U16523 ( .A(n16206), .B(n16205), .Z(n16210) );
  OR U16524 ( .A(n16208), .B(n16207), .Z(n16209) );
  AND U16525 ( .A(n16210), .B(n16209), .Z(n16283) );
  NANDN U16526 ( .A(n16212), .B(n16211), .Z(n16216) );
  NANDN U16527 ( .A(n16214), .B(n16213), .Z(n16215) );
  AND U16528 ( .A(n16216), .B(n16215), .Z(n16349) );
  NANDN U16529 ( .A(n16218), .B(n16217), .Z(n16222) );
  NANDN U16530 ( .A(n16220), .B(n16219), .Z(n16221) );
  NAND U16531 ( .A(n16222), .B(n16221), .Z(n16348) );
  XNOR U16532 ( .A(n16349), .B(n16348), .Z(n16351) );
  NANDN U16533 ( .A(n19394), .B(n16223), .Z(n16225) );
  XOR U16534 ( .A(b[29]), .B(a[96]), .Z(n16385) );
  NANDN U16535 ( .A(n19395), .B(n16385), .Z(n16224) );
  AND U16536 ( .A(n16225), .B(n16224), .Z(n16295) );
  AND U16537 ( .A(b[31]), .B(a[92]), .Z(n16294) );
  XNOR U16538 ( .A(n16295), .B(n16294), .Z(n16296) );
  NAND U16539 ( .A(b[0]), .B(a[124]), .Z(n16226) );
  XNOR U16540 ( .A(b[1]), .B(n16226), .Z(n16228) );
  NANDN U16541 ( .A(b[0]), .B(a[123]), .Z(n16227) );
  NAND U16542 ( .A(n16228), .B(n16227), .Z(n16297) );
  XNOR U16543 ( .A(n16296), .B(n16297), .Z(n16337) );
  NANDN U16544 ( .A(n19005), .B(n16229), .Z(n16231) );
  XOR U16545 ( .A(b[23]), .B(a[102]), .Z(n16373) );
  NANDN U16546 ( .A(n19055), .B(n16373), .Z(n16230) );
  AND U16547 ( .A(n16231), .B(n16230), .Z(n16390) );
  NANDN U16548 ( .A(n17362), .B(n16232), .Z(n16234) );
  XOR U16549 ( .A(a[118]), .B(b[7]), .Z(n16376) );
  NANDN U16550 ( .A(n17522), .B(n16376), .Z(n16233) );
  AND U16551 ( .A(n16234), .B(n16233), .Z(n16389) );
  NANDN U16552 ( .A(n19116), .B(n16235), .Z(n16237) );
  XOR U16553 ( .A(b[25]), .B(a[100]), .Z(n16379) );
  NANDN U16554 ( .A(n19179), .B(n16379), .Z(n16236) );
  NAND U16555 ( .A(n16237), .B(n16236), .Z(n16388) );
  XOR U16556 ( .A(n16389), .B(n16388), .Z(n16391) );
  XOR U16557 ( .A(n16390), .B(n16391), .Z(n16336) );
  XOR U16558 ( .A(n16337), .B(n16336), .Z(n16339) );
  NANDN U16559 ( .A(n18113), .B(n16238), .Z(n16240) );
  XOR U16560 ( .A(a[112]), .B(b[13]), .Z(n16358) );
  NANDN U16561 ( .A(n18229), .B(n16358), .Z(n16239) );
  AND U16562 ( .A(n16240), .B(n16239), .Z(n16331) );
  NANDN U16563 ( .A(n17888), .B(n16241), .Z(n16243) );
  XOR U16564 ( .A(a[114]), .B(b[11]), .Z(n16361) );
  NANDN U16565 ( .A(n18025), .B(n16361), .Z(n16242) );
  NAND U16566 ( .A(n16243), .B(n16242), .Z(n16330) );
  XNOR U16567 ( .A(n16331), .B(n16330), .Z(n16333) );
  NANDN U16568 ( .A(n18487), .B(n16244), .Z(n16246) );
  XOR U16569 ( .A(b[15]), .B(a[110]), .Z(n16364) );
  NANDN U16570 ( .A(n18311), .B(n16364), .Z(n16245) );
  AND U16571 ( .A(n16246), .B(n16245), .Z(n16327) );
  NANDN U16572 ( .A(n18853), .B(n16247), .Z(n16249) );
  XOR U16573 ( .A(b[21]), .B(a[104]), .Z(n16367) );
  NANDN U16574 ( .A(n18926), .B(n16367), .Z(n16248) );
  AND U16575 ( .A(n16249), .B(n16248), .Z(n16325) );
  NANDN U16576 ( .A(n17613), .B(n16250), .Z(n16252) );
  XOR U16577 ( .A(a[116]), .B(b[9]), .Z(n16370) );
  NANDN U16578 ( .A(n17739), .B(n16370), .Z(n16251) );
  NAND U16579 ( .A(n16252), .B(n16251), .Z(n16324) );
  XNOR U16580 ( .A(n16325), .B(n16324), .Z(n16326) );
  XNOR U16581 ( .A(n16327), .B(n16326), .Z(n16332) );
  XOR U16582 ( .A(n16333), .B(n16332), .Z(n16338) );
  XOR U16583 ( .A(n16339), .B(n16338), .Z(n16350) );
  XOR U16584 ( .A(n16351), .B(n16350), .Z(n16282) );
  XNOR U16585 ( .A(n16283), .B(n16282), .Z(n16284) );
  XOR U16586 ( .A(n16285), .B(n16284), .Z(n16277) );
  XNOR U16587 ( .A(n16276), .B(n16277), .Z(n16278) );
  XNOR U16588 ( .A(n16279), .B(n16278), .Z(n16272) );
  XOR U16589 ( .A(n16273), .B(n16272), .Z(n16401) );
  NANDN U16590 ( .A(n16254), .B(n16253), .Z(n16258) );
  NANDN U16591 ( .A(n16256), .B(n16255), .Z(n16257) );
  AND U16592 ( .A(n16258), .B(n16257), .Z(n16400) );
  XOR U16593 ( .A(n16401), .B(n16400), .Z(n16403) );
  XNOR U16594 ( .A(n16402), .B(n16403), .Z(n16264) );
  XNOR U16595 ( .A(n16265), .B(n16264), .Z(n16266) );
  XNOR U16596 ( .A(n16267), .B(n16266), .Z(n16406) );
  XNOR U16597 ( .A(sreg[220]), .B(n16406), .Z(n16408) );
  NANDN U16598 ( .A(sreg[219]), .B(n16259), .Z(n16263) );
  NAND U16599 ( .A(n16261), .B(n16260), .Z(n16262) );
  NAND U16600 ( .A(n16263), .B(n16262), .Z(n16407) );
  XNOR U16601 ( .A(n16408), .B(n16407), .Z(c[220]) );
  NANDN U16602 ( .A(n16265), .B(n16264), .Z(n16269) );
  NANDN U16603 ( .A(n16267), .B(n16266), .Z(n16268) );
  AND U16604 ( .A(n16269), .B(n16268), .Z(n16414) );
  NANDN U16605 ( .A(n16271), .B(n16270), .Z(n16275) );
  NAND U16606 ( .A(n16273), .B(n16272), .Z(n16274) );
  AND U16607 ( .A(n16275), .B(n16274), .Z(n16551) );
  NANDN U16608 ( .A(n16277), .B(n16276), .Z(n16281) );
  NANDN U16609 ( .A(n16279), .B(n16278), .Z(n16280) );
  AND U16610 ( .A(n16281), .B(n16280), .Z(n16550) );
  NANDN U16611 ( .A(n16283), .B(n16282), .Z(n16287) );
  NANDN U16612 ( .A(n16285), .B(n16284), .Z(n16286) );
  AND U16613 ( .A(n16287), .B(n16286), .Z(n16544) );
  NANDN U16614 ( .A(n16289), .B(n16288), .Z(n16293) );
  NAND U16615 ( .A(n16291), .B(n16290), .Z(n16292) );
  AND U16616 ( .A(n16293), .B(n16292), .Z(n16543) );
  XNOR U16617 ( .A(n16544), .B(n16543), .Z(n16545) );
  NANDN U16618 ( .A(n16295), .B(n16294), .Z(n16299) );
  NANDN U16619 ( .A(n16297), .B(n16296), .Z(n16298) );
  AND U16620 ( .A(n16299), .B(n16298), .Z(n16515) );
  NANDN U16621 ( .A(n19237), .B(n16300), .Z(n16302) );
  XOR U16622 ( .A(b[27]), .B(a[99]), .Z(n16429) );
  NANDN U16623 ( .A(n19277), .B(n16429), .Z(n16301) );
  AND U16624 ( .A(n16302), .B(n16301), .Z(n16504) );
  NANDN U16625 ( .A(n17072), .B(n16303), .Z(n16305) );
  XOR U16626 ( .A(a[121]), .B(b[5]), .Z(n16432) );
  NANDN U16627 ( .A(n17223), .B(n16432), .Z(n16304) );
  AND U16628 ( .A(n16305), .B(n16304), .Z(n16502) );
  NANDN U16629 ( .A(n18673), .B(n16306), .Z(n16308) );
  XOR U16630 ( .A(b[19]), .B(a[107]), .Z(n16435) );
  NANDN U16631 ( .A(n18758), .B(n16435), .Z(n16307) );
  NAND U16632 ( .A(n16308), .B(n16307), .Z(n16501) );
  XNOR U16633 ( .A(n16502), .B(n16501), .Z(n16503) );
  XNOR U16634 ( .A(n16504), .B(n16503), .Z(n16513) );
  NANDN U16635 ( .A(n19425), .B(n16309), .Z(n16311) );
  XOR U16636 ( .A(b[31]), .B(a[95]), .Z(n16438) );
  NANDN U16637 ( .A(n19426), .B(n16438), .Z(n16310) );
  AND U16638 ( .A(n16311), .B(n16310), .Z(n16456) );
  NANDN U16639 ( .A(n17067), .B(n16312), .Z(n16314) );
  XOR U16640 ( .A(a[123]), .B(b[3]), .Z(n16441) );
  NANDN U16641 ( .A(n17068), .B(n16441), .Z(n16313) );
  AND U16642 ( .A(n16314), .B(n16313), .Z(n16454) );
  NANDN U16643 ( .A(n18514), .B(n16315), .Z(n16317) );
  XOR U16644 ( .A(b[17]), .B(a[109]), .Z(n16444) );
  NANDN U16645 ( .A(n18585), .B(n16444), .Z(n16316) );
  NAND U16646 ( .A(n16317), .B(n16316), .Z(n16453) );
  XNOR U16647 ( .A(n16454), .B(n16453), .Z(n16455) );
  XOR U16648 ( .A(n16456), .B(n16455), .Z(n16514) );
  XOR U16649 ( .A(n16513), .B(n16514), .Z(n16516) );
  XOR U16650 ( .A(n16515), .B(n16516), .Z(n16526) );
  NANDN U16651 ( .A(n16319), .B(n16318), .Z(n16323) );
  NANDN U16652 ( .A(n16321), .B(n16320), .Z(n16322) );
  AND U16653 ( .A(n16323), .B(n16322), .Z(n16519) );
  NANDN U16654 ( .A(n16325), .B(n16324), .Z(n16329) );
  NANDN U16655 ( .A(n16327), .B(n16326), .Z(n16328) );
  NAND U16656 ( .A(n16329), .B(n16328), .Z(n16520) );
  XNOR U16657 ( .A(n16519), .B(n16520), .Z(n16521) );
  NANDN U16658 ( .A(n16331), .B(n16330), .Z(n16335) );
  NAND U16659 ( .A(n16333), .B(n16332), .Z(n16334) );
  NAND U16660 ( .A(n16335), .B(n16334), .Z(n16522) );
  XNOR U16661 ( .A(n16521), .B(n16522), .Z(n16525) );
  XNOR U16662 ( .A(n16526), .B(n16525), .Z(n16528) );
  NAND U16663 ( .A(n16337), .B(n16336), .Z(n16341) );
  NAND U16664 ( .A(n16339), .B(n16338), .Z(n16340) );
  AND U16665 ( .A(n16341), .B(n16340), .Z(n16527) );
  XOR U16666 ( .A(n16528), .B(n16527), .Z(n16540) );
  NANDN U16667 ( .A(n16343), .B(n16342), .Z(n16347) );
  NANDN U16668 ( .A(n16345), .B(n16344), .Z(n16346) );
  AND U16669 ( .A(n16347), .B(n16346), .Z(n16537) );
  NANDN U16670 ( .A(n16353), .B(n16352), .Z(n16357) );
  OR U16671 ( .A(n16355), .B(n16354), .Z(n16356) );
  AND U16672 ( .A(n16357), .B(n16356), .Z(n16532) );
  NANDN U16673 ( .A(n18113), .B(n16358), .Z(n16360) );
  XOR U16674 ( .A(a[113]), .B(b[13]), .Z(n16471) );
  NANDN U16675 ( .A(n18229), .B(n16471), .Z(n16359) );
  AND U16676 ( .A(n16360), .B(n16359), .Z(n16462) );
  NANDN U16677 ( .A(n17888), .B(n16361), .Z(n16363) );
  XOR U16678 ( .A(a[115]), .B(b[11]), .Z(n16474) );
  NANDN U16679 ( .A(n18025), .B(n16474), .Z(n16362) );
  AND U16680 ( .A(n16363), .B(n16362), .Z(n16460) );
  NANDN U16681 ( .A(n18487), .B(n16364), .Z(n16366) );
  XOR U16682 ( .A(b[15]), .B(a[111]), .Z(n16477) );
  NANDN U16683 ( .A(n18311), .B(n16477), .Z(n16365) );
  AND U16684 ( .A(n16366), .B(n16365), .Z(n16450) );
  NANDN U16685 ( .A(n18853), .B(n16367), .Z(n16369) );
  XOR U16686 ( .A(b[21]), .B(a[105]), .Z(n16480) );
  NANDN U16687 ( .A(n18926), .B(n16480), .Z(n16368) );
  AND U16688 ( .A(n16369), .B(n16368), .Z(n16448) );
  NANDN U16689 ( .A(n17613), .B(n16370), .Z(n16372) );
  XOR U16690 ( .A(a[117]), .B(b[9]), .Z(n16483) );
  NANDN U16691 ( .A(n17739), .B(n16483), .Z(n16371) );
  NAND U16692 ( .A(n16372), .B(n16371), .Z(n16447) );
  XNOR U16693 ( .A(n16448), .B(n16447), .Z(n16449) );
  XNOR U16694 ( .A(n16450), .B(n16449), .Z(n16459) );
  XNOR U16695 ( .A(n16460), .B(n16459), .Z(n16461) );
  XOR U16696 ( .A(n16462), .B(n16461), .Z(n16419) );
  NANDN U16697 ( .A(n19005), .B(n16373), .Z(n16375) );
  XOR U16698 ( .A(b[23]), .B(a[103]), .Z(n16486) );
  NANDN U16699 ( .A(n19055), .B(n16486), .Z(n16374) );
  AND U16700 ( .A(n16375), .B(n16374), .Z(n16510) );
  NANDN U16701 ( .A(n17362), .B(n16376), .Z(n16378) );
  XOR U16702 ( .A(a[119]), .B(b[7]), .Z(n16489) );
  NANDN U16703 ( .A(n17522), .B(n16489), .Z(n16377) );
  AND U16704 ( .A(n16378), .B(n16377), .Z(n16508) );
  NANDN U16705 ( .A(n19116), .B(n16379), .Z(n16381) );
  XOR U16706 ( .A(b[25]), .B(a[101]), .Z(n16492) );
  NANDN U16707 ( .A(n19179), .B(n16492), .Z(n16380) );
  NAND U16708 ( .A(n16381), .B(n16380), .Z(n16507) );
  XNOR U16709 ( .A(n16508), .B(n16507), .Z(n16509) );
  XOR U16710 ( .A(n16510), .B(n16509), .Z(n16418) );
  NAND U16711 ( .A(b[0]), .B(a[125]), .Z(n16382) );
  XNOR U16712 ( .A(b[1]), .B(n16382), .Z(n16384) );
  NANDN U16713 ( .A(b[0]), .B(a[124]), .Z(n16383) );
  NAND U16714 ( .A(n16384), .B(n16383), .Z(n16426) );
  NANDN U16715 ( .A(n19394), .B(n16385), .Z(n16387) );
  XOR U16716 ( .A(b[29]), .B(a[97]), .Z(n16498) );
  NANDN U16717 ( .A(n19395), .B(n16498), .Z(n16386) );
  AND U16718 ( .A(n16387), .B(n16386), .Z(n16424) );
  AND U16719 ( .A(b[31]), .B(a[93]), .Z(n16423) );
  XNOR U16720 ( .A(n16424), .B(n16423), .Z(n16425) );
  XOR U16721 ( .A(n16426), .B(n16425), .Z(n16417) );
  XNOR U16722 ( .A(n16418), .B(n16417), .Z(n16420) );
  NANDN U16723 ( .A(n16389), .B(n16388), .Z(n16393) );
  OR U16724 ( .A(n16391), .B(n16390), .Z(n16392) );
  AND U16725 ( .A(n16393), .B(n16392), .Z(n16466) );
  NANDN U16726 ( .A(n16395), .B(n16394), .Z(n16399) );
  NANDN U16727 ( .A(n16397), .B(n16396), .Z(n16398) );
  NAND U16728 ( .A(n16399), .B(n16398), .Z(n16465) );
  XNOR U16729 ( .A(n16466), .B(n16465), .Z(n16467) );
  XOR U16730 ( .A(n16468), .B(n16467), .Z(n16531) );
  XNOR U16731 ( .A(n16532), .B(n16531), .Z(n16533) );
  XOR U16732 ( .A(n16534), .B(n16533), .Z(n16538) );
  XNOR U16733 ( .A(n16537), .B(n16538), .Z(n16539) );
  XOR U16734 ( .A(n16540), .B(n16539), .Z(n16546) );
  XNOR U16735 ( .A(n16545), .B(n16546), .Z(n16549) );
  XOR U16736 ( .A(n16550), .B(n16549), .Z(n16552) );
  XOR U16737 ( .A(n16551), .B(n16552), .Z(n16412) );
  NANDN U16738 ( .A(n16401), .B(n16400), .Z(n16405) );
  NANDN U16739 ( .A(n16403), .B(n16402), .Z(n16404) );
  NAND U16740 ( .A(n16405), .B(n16404), .Z(n16411) );
  XNOR U16741 ( .A(n16412), .B(n16411), .Z(n16413) );
  XNOR U16742 ( .A(n16414), .B(n16413), .Z(n16555) );
  XNOR U16743 ( .A(sreg[221]), .B(n16555), .Z(n16557) );
  NANDN U16744 ( .A(sreg[220]), .B(n16406), .Z(n16410) );
  NAND U16745 ( .A(n16408), .B(n16407), .Z(n16409) );
  NAND U16746 ( .A(n16410), .B(n16409), .Z(n16556) );
  XNOR U16747 ( .A(n16557), .B(n16556), .Z(c[221]) );
  NANDN U16748 ( .A(n16412), .B(n16411), .Z(n16416) );
  NANDN U16749 ( .A(n16414), .B(n16413), .Z(n16415) );
  AND U16750 ( .A(n16416), .B(n16415), .Z(n16563) );
  NAND U16751 ( .A(n16418), .B(n16417), .Z(n16422) );
  NANDN U16752 ( .A(n16420), .B(n16419), .Z(n16421) );
  AND U16753 ( .A(n16422), .B(n16421), .Z(n16692) );
  NANDN U16754 ( .A(n16424), .B(n16423), .Z(n16428) );
  NANDN U16755 ( .A(n16426), .B(n16425), .Z(n16427) );
  AND U16756 ( .A(n16428), .B(n16427), .Z(n16592) );
  NANDN U16757 ( .A(n19237), .B(n16429), .Z(n16431) );
  XOR U16758 ( .A(b[27]), .B(a[100]), .Z(n16668) );
  NANDN U16759 ( .A(n19277), .B(n16668), .Z(n16430) );
  AND U16760 ( .A(n16431), .B(n16430), .Z(n16635) );
  NANDN U16761 ( .A(n17072), .B(n16432), .Z(n16434) );
  XOR U16762 ( .A(a[122]), .B(b[5]), .Z(n16671) );
  NANDN U16763 ( .A(n17223), .B(n16671), .Z(n16433) );
  AND U16764 ( .A(n16434), .B(n16433), .Z(n16633) );
  NANDN U16765 ( .A(n18673), .B(n16435), .Z(n16437) );
  XOR U16766 ( .A(b[19]), .B(a[108]), .Z(n16674) );
  NANDN U16767 ( .A(n18758), .B(n16674), .Z(n16436) );
  NAND U16768 ( .A(n16437), .B(n16436), .Z(n16632) );
  XNOR U16769 ( .A(n16633), .B(n16632), .Z(n16634) );
  XNOR U16770 ( .A(n16635), .B(n16634), .Z(n16590) );
  NANDN U16771 ( .A(n19425), .B(n16438), .Z(n16440) );
  XOR U16772 ( .A(b[31]), .B(a[96]), .Z(n16677) );
  NANDN U16773 ( .A(n19426), .B(n16677), .Z(n16439) );
  AND U16774 ( .A(n16440), .B(n16439), .Z(n16653) );
  NANDN U16775 ( .A(n17067), .B(n16441), .Z(n16443) );
  XOR U16776 ( .A(a[124]), .B(b[3]), .Z(n16680) );
  NANDN U16777 ( .A(n17068), .B(n16680), .Z(n16442) );
  AND U16778 ( .A(n16443), .B(n16442), .Z(n16651) );
  NANDN U16779 ( .A(n18514), .B(n16444), .Z(n16446) );
  XOR U16780 ( .A(b[17]), .B(a[110]), .Z(n16683) );
  NANDN U16781 ( .A(n18585), .B(n16683), .Z(n16445) );
  NAND U16782 ( .A(n16446), .B(n16445), .Z(n16650) );
  XNOR U16783 ( .A(n16651), .B(n16650), .Z(n16652) );
  XOR U16784 ( .A(n16653), .B(n16652), .Z(n16591) );
  XOR U16785 ( .A(n16590), .B(n16591), .Z(n16593) );
  XOR U16786 ( .A(n16592), .B(n16593), .Z(n16691) );
  NANDN U16787 ( .A(n16448), .B(n16447), .Z(n16452) );
  NANDN U16788 ( .A(n16450), .B(n16449), .Z(n16451) );
  AND U16789 ( .A(n16452), .B(n16451), .Z(n16578) );
  NANDN U16790 ( .A(n16454), .B(n16453), .Z(n16458) );
  NANDN U16791 ( .A(n16456), .B(n16455), .Z(n16457) );
  NAND U16792 ( .A(n16458), .B(n16457), .Z(n16579) );
  XNOR U16793 ( .A(n16578), .B(n16579), .Z(n16580) );
  NANDN U16794 ( .A(n16460), .B(n16459), .Z(n16464) );
  NANDN U16795 ( .A(n16462), .B(n16461), .Z(n16463) );
  NAND U16796 ( .A(n16464), .B(n16463), .Z(n16581) );
  XNOR U16797 ( .A(n16580), .B(n16581), .Z(n16690) );
  XOR U16798 ( .A(n16691), .B(n16690), .Z(n16693) );
  XOR U16799 ( .A(n16692), .B(n16693), .Z(n16574) );
  NANDN U16800 ( .A(n16466), .B(n16465), .Z(n16470) );
  NAND U16801 ( .A(n16468), .B(n16467), .Z(n16469) );
  AND U16802 ( .A(n16470), .B(n16469), .Z(n16689) );
  NANDN U16803 ( .A(n18113), .B(n16471), .Z(n16473) );
  XOR U16804 ( .A(a[114]), .B(b[13]), .Z(n16596) );
  NANDN U16805 ( .A(n18229), .B(n16596), .Z(n16472) );
  AND U16806 ( .A(n16473), .B(n16472), .Z(n16659) );
  NANDN U16807 ( .A(n17888), .B(n16474), .Z(n16476) );
  XOR U16808 ( .A(a[116]), .B(b[11]), .Z(n16599) );
  NANDN U16809 ( .A(n18025), .B(n16599), .Z(n16475) );
  AND U16810 ( .A(n16476), .B(n16475), .Z(n16657) );
  NANDN U16811 ( .A(n18487), .B(n16477), .Z(n16479) );
  XOR U16812 ( .A(b[15]), .B(a[112]), .Z(n16602) );
  NANDN U16813 ( .A(n18311), .B(n16602), .Z(n16478) );
  AND U16814 ( .A(n16479), .B(n16478), .Z(n16647) );
  NANDN U16815 ( .A(n18853), .B(n16480), .Z(n16482) );
  XOR U16816 ( .A(b[21]), .B(a[106]), .Z(n16605) );
  NANDN U16817 ( .A(n18926), .B(n16605), .Z(n16481) );
  AND U16818 ( .A(n16482), .B(n16481), .Z(n16645) );
  NANDN U16819 ( .A(n17613), .B(n16483), .Z(n16485) );
  XOR U16820 ( .A(a[118]), .B(b[9]), .Z(n16608) );
  NANDN U16821 ( .A(n17739), .B(n16608), .Z(n16484) );
  NAND U16822 ( .A(n16485), .B(n16484), .Z(n16644) );
  XNOR U16823 ( .A(n16645), .B(n16644), .Z(n16646) );
  XNOR U16824 ( .A(n16647), .B(n16646), .Z(n16656) );
  XNOR U16825 ( .A(n16657), .B(n16656), .Z(n16658) );
  XOR U16826 ( .A(n16659), .B(n16658), .Z(n16640) );
  NANDN U16827 ( .A(n19005), .B(n16486), .Z(n16488) );
  XOR U16828 ( .A(b[23]), .B(a[104]), .Z(n16611) );
  NANDN U16829 ( .A(n19055), .B(n16611), .Z(n16487) );
  AND U16830 ( .A(n16488), .B(n16487), .Z(n16629) );
  NANDN U16831 ( .A(n17362), .B(n16489), .Z(n16491) );
  XOR U16832 ( .A(a[120]), .B(b[7]), .Z(n16614) );
  NANDN U16833 ( .A(n17522), .B(n16614), .Z(n16490) );
  AND U16834 ( .A(n16491), .B(n16490), .Z(n16627) );
  NANDN U16835 ( .A(n19116), .B(n16492), .Z(n16494) );
  XOR U16836 ( .A(b[25]), .B(a[102]), .Z(n16617) );
  NANDN U16837 ( .A(n19179), .B(n16617), .Z(n16493) );
  NAND U16838 ( .A(n16494), .B(n16493), .Z(n16626) );
  XNOR U16839 ( .A(n16627), .B(n16626), .Z(n16628) );
  XOR U16840 ( .A(n16629), .B(n16628), .Z(n16639) );
  NAND U16841 ( .A(b[0]), .B(a[126]), .Z(n16495) );
  XNOR U16842 ( .A(b[1]), .B(n16495), .Z(n16497) );
  NANDN U16843 ( .A(b[0]), .B(a[125]), .Z(n16496) );
  NAND U16844 ( .A(n16497), .B(n16496), .Z(n16665) );
  NANDN U16845 ( .A(n19394), .B(n16498), .Z(n16500) );
  XOR U16846 ( .A(b[29]), .B(a[98]), .Z(n16620) );
  NANDN U16847 ( .A(n19395), .B(n16620), .Z(n16499) );
  AND U16848 ( .A(n16500), .B(n16499), .Z(n16663) );
  AND U16849 ( .A(b[31]), .B(a[94]), .Z(n16662) );
  XNOR U16850 ( .A(n16663), .B(n16662), .Z(n16664) );
  XOR U16851 ( .A(n16665), .B(n16664), .Z(n16638) );
  XOR U16852 ( .A(n16639), .B(n16638), .Z(n16641) );
  XNOR U16853 ( .A(n16640), .B(n16641), .Z(n16586) );
  NANDN U16854 ( .A(n16502), .B(n16501), .Z(n16506) );
  NANDN U16855 ( .A(n16504), .B(n16503), .Z(n16505) );
  AND U16856 ( .A(n16506), .B(n16505), .Z(n16585) );
  NANDN U16857 ( .A(n16508), .B(n16507), .Z(n16512) );
  NANDN U16858 ( .A(n16510), .B(n16509), .Z(n16511) );
  NAND U16859 ( .A(n16512), .B(n16511), .Z(n16584) );
  XOR U16860 ( .A(n16585), .B(n16584), .Z(n16587) );
  XOR U16861 ( .A(n16586), .B(n16587), .Z(n16686) );
  NANDN U16862 ( .A(n16514), .B(n16513), .Z(n16518) );
  OR U16863 ( .A(n16516), .B(n16515), .Z(n16517) );
  AND U16864 ( .A(n16518), .B(n16517), .Z(n16687) );
  XOR U16865 ( .A(n16686), .B(n16687), .Z(n16688) );
  XOR U16866 ( .A(n16689), .B(n16688), .Z(n16573) );
  NANDN U16867 ( .A(n16520), .B(n16519), .Z(n16524) );
  NANDN U16868 ( .A(n16522), .B(n16521), .Z(n16523) );
  AND U16869 ( .A(n16524), .B(n16523), .Z(n16572) );
  XOR U16870 ( .A(n16573), .B(n16572), .Z(n16575) );
  XOR U16871 ( .A(n16574), .B(n16575), .Z(n16569) );
  NANDN U16872 ( .A(n16526), .B(n16525), .Z(n16530) );
  NAND U16873 ( .A(n16528), .B(n16527), .Z(n16529) );
  AND U16874 ( .A(n16530), .B(n16529), .Z(n16567) );
  NANDN U16875 ( .A(n16532), .B(n16531), .Z(n16536) );
  NANDN U16876 ( .A(n16534), .B(n16533), .Z(n16535) );
  AND U16877 ( .A(n16536), .B(n16535), .Z(n16566) );
  XNOR U16878 ( .A(n16567), .B(n16566), .Z(n16568) );
  XNOR U16879 ( .A(n16569), .B(n16568), .Z(n16696) );
  NANDN U16880 ( .A(n16538), .B(n16537), .Z(n16542) );
  NANDN U16881 ( .A(n16540), .B(n16539), .Z(n16541) );
  NAND U16882 ( .A(n16542), .B(n16541), .Z(n16697) );
  XNOR U16883 ( .A(n16696), .B(n16697), .Z(n16698) );
  NANDN U16884 ( .A(n16544), .B(n16543), .Z(n16548) );
  NANDN U16885 ( .A(n16546), .B(n16545), .Z(n16547) );
  NAND U16886 ( .A(n16548), .B(n16547), .Z(n16699) );
  XNOR U16887 ( .A(n16698), .B(n16699), .Z(n16560) );
  NANDN U16888 ( .A(n16550), .B(n16549), .Z(n16554) );
  OR U16889 ( .A(n16552), .B(n16551), .Z(n16553) );
  NAND U16890 ( .A(n16554), .B(n16553), .Z(n16561) );
  XNOR U16891 ( .A(n16560), .B(n16561), .Z(n16562) );
  XNOR U16892 ( .A(n16563), .B(n16562), .Z(n16702) );
  XNOR U16893 ( .A(sreg[222]), .B(n16702), .Z(n16704) );
  NANDN U16894 ( .A(sreg[221]), .B(n16555), .Z(n16559) );
  NAND U16895 ( .A(n16557), .B(n16556), .Z(n16558) );
  NAND U16896 ( .A(n16559), .B(n16558), .Z(n16703) );
  XNOR U16897 ( .A(n16704), .B(n16703), .Z(c[222]) );
  NANDN U16898 ( .A(n16561), .B(n16560), .Z(n16565) );
  NANDN U16899 ( .A(n16563), .B(n16562), .Z(n16564) );
  AND U16900 ( .A(n16565), .B(n16564), .Z(n16715) );
  NANDN U16901 ( .A(n16567), .B(n16566), .Z(n16571) );
  NANDN U16902 ( .A(n16569), .B(n16568), .Z(n16570) );
  AND U16903 ( .A(n16571), .B(n16570), .Z(n16850) );
  NANDN U16904 ( .A(n16573), .B(n16572), .Z(n16577) );
  OR U16905 ( .A(n16575), .B(n16574), .Z(n16576) );
  AND U16906 ( .A(n16577), .B(n16576), .Z(n16848) );
  NANDN U16907 ( .A(n16579), .B(n16578), .Z(n16583) );
  NANDN U16908 ( .A(n16581), .B(n16580), .Z(n16582) );
  AND U16909 ( .A(n16583), .B(n16582), .Z(n16724) );
  NANDN U16910 ( .A(n16585), .B(n16584), .Z(n16589) );
  NANDN U16911 ( .A(n16587), .B(n16586), .Z(n16588) );
  AND U16912 ( .A(n16589), .B(n16588), .Z(n16838) );
  NANDN U16913 ( .A(n16591), .B(n16590), .Z(n16595) );
  OR U16914 ( .A(n16593), .B(n16592), .Z(n16594) );
  AND U16915 ( .A(n16595), .B(n16594), .Z(n16836) );
  NANDN U16916 ( .A(n18113), .B(n16596), .Z(n16598) );
  XOR U16917 ( .A(a[115]), .B(b[13]), .Z(n16793) );
  NANDN U16918 ( .A(n18229), .B(n16793), .Z(n16597) );
  AND U16919 ( .A(n16598), .B(n16597), .Z(n16774) );
  NANDN U16920 ( .A(n17888), .B(n16599), .Z(n16601) );
  XOR U16921 ( .A(a[117]), .B(b[11]), .Z(n16790) );
  NANDN U16922 ( .A(n18025), .B(n16790), .Z(n16600) );
  AND U16923 ( .A(n16601), .B(n16600), .Z(n16773) );
  NANDN U16924 ( .A(n18487), .B(n16602), .Z(n16604) );
  XOR U16925 ( .A(b[15]), .B(a[113]), .Z(n16796) );
  NANDN U16926 ( .A(n18311), .B(n16796), .Z(n16603) );
  AND U16927 ( .A(n16604), .B(n16603), .Z(n16763) );
  NANDN U16928 ( .A(n18853), .B(n16605), .Z(n16607) );
  XOR U16929 ( .A(b[21]), .B(a[107]), .Z(n16799) );
  NANDN U16930 ( .A(n18926), .B(n16799), .Z(n16606) );
  AND U16931 ( .A(n16607), .B(n16606), .Z(n16761) );
  NANDN U16932 ( .A(n17613), .B(n16608), .Z(n16610) );
  XOR U16933 ( .A(a[119]), .B(b[9]), .Z(n16802) );
  NANDN U16934 ( .A(n17739), .B(n16802), .Z(n16609) );
  NAND U16935 ( .A(n16610), .B(n16609), .Z(n16760) );
  XNOR U16936 ( .A(n16761), .B(n16760), .Z(n16762) );
  XNOR U16937 ( .A(n16763), .B(n16762), .Z(n16772) );
  XOR U16938 ( .A(n16773), .B(n16772), .Z(n16775) );
  XOR U16939 ( .A(n16774), .B(n16775), .Z(n16732) );
  NANDN U16940 ( .A(n19005), .B(n16611), .Z(n16613) );
  XOR U16941 ( .A(b[23]), .B(a[105]), .Z(n16805) );
  NANDN U16942 ( .A(n19055), .B(n16805), .Z(n16612) );
  AND U16943 ( .A(n16613), .B(n16612), .Z(n16825) );
  NANDN U16944 ( .A(n17362), .B(n16614), .Z(n16616) );
  XOR U16945 ( .A(a[121]), .B(b[7]), .Z(n16808) );
  NANDN U16946 ( .A(n17522), .B(n16808), .Z(n16615) );
  AND U16947 ( .A(n16616), .B(n16615), .Z(n16824) );
  NANDN U16948 ( .A(n19116), .B(n16617), .Z(n16619) );
  XOR U16949 ( .A(b[25]), .B(a[103]), .Z(n16811) );
  NANDN U16950 ( .A(n19179), .B(n16811), .Z(n16618) );
  NAND U16951 ( .A(n16619), .B(n16618), .Z(n16823) );
  XOR U16952 ( .A(n16824), .B(n16823), .Z(n16826) );
  XOR U16953 ( .A(n16825), .B(n16826), .Z(n16731) );
  NANDN U16954 ( .A(n19394), .B(n16620), .Z(n16622) );
  XOR U16955 ( .A(b[29]), .B(a[99]), .Z(n16814) );
  NANDN U16956 ( .A(n19395), .B(n16814), .Z(n16621) );
  AND U16957 ( .A(n16622), .B(n16621), .Z(n16737) );
  AND U16958 ( .A(b[31]), .B(a[95]), .Z(n16736) );
  XOR U16959 ( .A(n16737), .B(n16736), .Z(n16738) );
  NAND U16960 ( .A(b[0]), .B(a[127]), .Z(n16623) );
  XNOR U16961 ( .A(b[1]), .B(n16623), .Z(n16625) );
  NANDN U16962 ( .A(b[0]), .B(a[126]), .Z(n16624) );
  NAND U16963 ( .A(n16625), .B(n16624), .Z(n16739) );
  XNOR U16964 ( .A(n16738), .B(n16739), .Z(n16730) );
  XOR U16965 ( .A(n16731), .B(n16730), .Z(n16733) );
  XOR U16966 ( .A(n16732), .B(n16733), .Z(n16787) );
  NANDN U16967 ( .A(n16627), .B(n16626), .Z(n16631) );
  NANDN U16968 ( .A(n16629), .B(n16628), .Z(n16630) );
  AND U16969 ( .A(n16631), .B(n16630), .Z(n16785) );
  NANDN U16970 ( .A(n16633), .B(n16632), .Z(n16637) );
  NANDN U16971 ( .A(n16635), .B(n16634), .Z(n16636) );
  NAND U16972 ( .A(n16637), .B(n16636), .Z(n16784) );
  XNOR U16973 ( .A(n16785), .B(n16784), .Z(n16786) );
  XNOR U16974 ( .A(n16787), .B(n16786), .Z(n16835) );
  XNOR U16975 ( .A(n16836), .B(n16835), .Z(n16837) );
  XOR U16976 ( .A(n16838), .B(n16837), .Z(n16725) );
  XNOR U16977 ( .A(n16724), .B(n16725), .Z(n16727) );
  NAND U16978 ( .A(n16639), .B(n16638), .Z(n16643) );
  NAND U16979 ( .A(n16641), .B(n16640), .Z(n16642) );
  AND U16980 ( .A(n16643), .B(n16642), .Z(n16843) );
  NANDN U16981 ( .A(n16645), .B(n16644), .Z(n16649) );
  NANDN U16982 ( .A(n16647), .B(n16646), .Z(n16648) );
  AND U16983 ( .A(n16649), .B(n16648), .Z(n16778) );
  NANDN U16984 ( .A(n16651), .B(n16650), .Z(n16655) );
  NANDN U16985 ( .A(n16653), .B(n16652), .Z(n16654) );
  NAND U16986 ( .A(n16655), .B(n16654), .Z(n16779) );
  XNOR U16987 ( .A(n16778), .B(n16779), .Z(n16781) );
  NANDN U16988 ( .A(n16657), .B(n16656), .Z(n16661) );
  NANDN U16989 ( .A(n16659), .B(n16658), .Z(n16660) );
  AND U16990 ( .A(n16661), .B(n16660), .Z(n16780) );
  XOR U16991 ( .A(n16781), .B(n16780), .Z(n16842) );
  NANDN U16992 ( .A(n16663), .B(n16662), .Z(n16667) );
  NANDN U16993 ( .A(n16665), .B(n16664), .Z(n16666) );
  AND U16994 ( .A(n16667), .B(n16666), .Z(n16832) );
  NANDN U16995 ( .A(n19237), .B(n16668), .Z(n16670) );
  XOR U16996 ( .A(b[27]), .B(a[101]), .Z(n16742) );
  NANDN U16997 ( .A(n19277), .B(n16742), .Z(n16669) );
  AND U16998 ( .A(n16670), .B(n16669), .Z(n16820) );
  NANDN U16999 ( .A(n17072), .B(n16671), .Z(n16673) );
  XOR U17000 ( .A(a[123]), .B(b[5]), .Z(n16745) );
  NANDN U17001 ( .A(n17223), .B(n16745), .Z(n16672) );
  AND U17002 ( .A(n16673), .B(n16672), .Z(n16818) );
  NANDN U17003 ( .A(n18673), .B(n16674), .Z(n16676) );
  XOR U17004 ( .A(b[19]), .B(a[109]), .Z(n16748) );
  NANDN U17005 ( .A(n18758), .B(n16748), .Z(n16675) );
  NAND U17006 ( .A(n16676), .B(n16675), .Z(n16817) );
  XNOR U17007 ( .A(n16818), .B(n16817), .Z(n16819) );
  XNOR U17008 ( .A(n16820), .B(n16819), .Z(n16829) );
  NANDN U17009 ( .A(n19425), .B(n16677), .Z(n16679) );
  XOR U17010 ( .A(b[31]), .B(a[97]), .Z(n16751) );
  NANDN U17011 ( .A(n19426), .B(n16751), .Z(n16678) );
  AND U17012 ( .A(n16679), .B(n16678), .Z(n16769) );
  NANDN U17013 ( .A(n17067), .B(n16680), .Z(n16682) );
  XOR U17014 ( .A(a[125]), .B(b[3]), .Z(n16754) );
  NANDN U17015 ( .A(n17068), .B(n16754), .Z(n16681) );
  AND U17016 ( .A(n16682), .B(n16681), .Z(n16767) );
  NANDN U17017 ( .A(n18514), .B(n16683), .Z(n16685) );
  XOR U17018 ( .A(b[17]), .B(a[111]), .Z(n16757) );
  NANDN U17019 ( .A(n18585), .B(n16757), .Z(n16684) );
  NAND U17020 ( .A(n16685), .B(n16684), .Z(n16766) );
  XNOR U17021 ( .A(n16767), .B(n16766), .Z(n16768) );
  XOR U17022 ( .A(n16769), .B(n16768), .Z(n16830) );
  XNOR U17023 ( .A(n16829), .B(n16830), .Z(n16831) );
  XNOR U17024 ( .A(n16832), .B(n16831), .Z(n16841) );
  XOR U17025 ( .A(n16842), .B(n16841), .Z(n16844) );
  XNOR U17026 ( .A(n16843), .B(n16844), .Z(n16726) );
  XOR U17027 ( .A(n16727), .B(n16726), .Z(n16720) );
  NANDN U17028 ( .A(n16691), .B(n16690), .Z(n16695) );
  OR U17029 ( .A(n16693), .B(n16692), .Z(n16694) );
  NAND U17030 ( .A(n16695), .B(n16694), .Z(n16718) );
  XOR U17031 ( .A(n16719), .B(n16718), .Z(n16721) );
  XNOR U17032 ( .A(n16720), .B(n16721), .Z(n16847) );
  XNOR U17033 ( .A(n16848), .B(n16847), .Z(n16849) );
  XOR U17034 ( .A(n16850), .B(n16849), .Z(n16713) );
  NANDN U17035 ( .A(n16697), .B(n16696), .Z(n16701) );
  NANDN U17036 ( .A(n16699), .B(n16698), .Z(n16700) );
  NAND U17037 ( .A(n16701), .B(n16700), .Z(n16712) );
  XNOR U17038 ( .A(n16713), .B(n16712), .Z(n16714) );
  XNOR U17039 ( .A(n16715), .B(n16714), .Z(n16707) );
  XNOR U17040 ( .A(sreg[223]), .B(n16707), .Z(n16709) );
  NANDN U17041 ( .A(sreg[222]), .B(n16702), .Z(n16706) );
  NAND U17042 ( .A(n16704), .B(n16703), .Z(n16705) );
  NAND U17043 ( .A(n16706), .B(n16705), .Z(n16708) );
  XNOR U17044 ( .A(n16709), .B(n16708), .Z(c[223]) );
  NANDN U17045 ( .A(sreg[223]), .B(n16707), .Z(n16711) );
  NAND U17046 ( .A(n16709), .B(n16708), .Z(n16710) );
  AND U17047 ( .A(n16711), .B(n16710), .Z(n16854) );
  NANDN U17048 ( .A(n16713), .B(n16712), .Z(n16717) );
  NANDN U17049 ( .A(n16715), .B(n16714), .Z(n16716) );
  AND U17050 ( .A(n16717), .B(n16716), .Z(n16857) );
  NANDN U17051 ( .A(n16719), .B(n16718), .Z(n16723) );
  OR U17052 ( .A(n16721), .B(n16720), .Z(n16722) );
  AND U17053 ( .A(n16723), .B(n16722), .Z(n16993) );
  NANDN U17054 ( .A(n16725), .B(n16724), .Z(n16729) );
  NAND U17055 ( .A(n16727), .B(n16726), .Z(n16728) );
  AND U17056 ( .A(n16729), .B(n16728), .Z(n16991) );
  NANDN U17057 ( .A(n16731), .B(n16730), .Z(n16735) );
  OR U17058 ( .A(n16733), .B(n16732), .Z(n16734) );
  AND U17059 ( .A(n16735), .B(n16734), .Z(n16881) );
  NANDN U17060 ( .A(n16737), .B(n16736), .Z(n16741) );
  OR U17061 ( .A(n16739), .B(n16738), .Z(n16740) );
  AND U17062 ( .A(n16741), .B(n16740), .Z(n16938) );
  NANDN U17063 ( .A(n19237), .B(n16742), .Z(n16744) );
  XOR U17064 ( .A(b[27]), .B(a[102]), .Z(n16897) );
  NANDN U17065 ( .A(n19277), .B(n16897), .Z(n16743) );
  AND U17066 ( .A(n16744), .B(n16743), .Z(n16981) );
  NANDN U17067 ( .A(n17072), .B(n16745), .Z(n16747) );
  XOR U17068 ( .A(a[124]), .B(b[5]), .Z(n16960) );
  NANDN U17069 ( .A(n17223), .B(n16960), .Z(n16746) );
  AND U17070 ( .A(n16747), .B(n16746), .Z(n16979) );
  NANDN U17071 ( .A(n18673), .B(n16748), .Z(n16750) );
  XOR U17072 ( .A(b[19]), .B(a[110]), .Z(n16951) );
  NANDN U17073 ( .A(n18758), .B(n16951), .Z(n16749) );
  NAND U17074 ( .A(n16750), .B(n16749), .Z(n16978) );
  XNOR U17075 ( .A(n16979), .B(n16978), .Z(n16980) );
  XNOR U17076 ( .A(n16981), .B(n16980), .Z(n16936) );
  NANDN U17077 ( .A(n19425), .B(n16751), .Z(n16753) );
  XOR U17078 ( .A(b[31]), .B(a[98]), .Z(n16966) );
  NANDN U17079 ( .A(n19426), .B(n16966), .Z(n16752) );
  AND U17080 ( .A(n16753), .B(n16752), .Z(n16921) );
  NANDN U17081 ( .A(n17067), .B(n16754), .Z(n16756) );
  XOR U17082 ( .A(a[126]), .B(b[3]), .Z(n16906) );
  NANDN U17083 ( .A(n17068), .B(n16906), .Z(n16755) );
  AND U17084 ( .A(n16756), .B(n16755), .Z(n16919) );
  NANDN U17085 ( .A(n18514), .B(n16757), .Z(n16759) );
  XOR U17086 ( .A(b[17]), .B(a[112]), .Z(n16909) );
  NANDN U17087 ( .A(n18585), .B(n16909), .Z(n16758) );
  NAND U17088 ( .A(n16759), .B(n16758), .Z(n16918) );
  XNOR U17089 ( .A(n16919), .B(n16918), .Z(n16920) );
  XOR U17090 ( .A(n16921), .B(n16920), .Z(n16937) );
  XOR U17091 ( .A(n16936), .B(n16937), .Z(n16939) );
  XOR U17092 ( .A(n16938), .B(n16939), .Z(n16880) );
  NANDN U17093 ( .A(n16761), .B(n16760), .Z(n16765) );
  NANDN U17094 ( .A(n16763), .B(n16762), .Z(n16764) );
  AND U17095 ( .A(n16765), .B(n16764), .Z(n16930) );
  NANDN U17096 ( .A(n16767), .B(n16766), .Z(n16771) );
  NANDN U17097 ( .A(n16769), .B(n16768), .Z(n16770) );
  NAND U17098 ( .A(n16771), .B(n16770), .Z(n16931) );
  XNOR U17099 ( .A(n16930), .B(n16931), .Z(n16932) );
  NANDN U17100 ( .A(n16773), .B(n16772), .Z(n16777) );
  OR U17101 ( .A(n16775), .B(n16774), .Z(n16776) );
  NAND U17102 ( .A(n16777), .B(n16776), .Z(n16933) );
  XNOR U17103 ( .A(n16932), .B(n16933), .Z(n16879) );
  XOR U17104 ( .A(n16880), .B(n16879), .Z(n16882) );
  XOR U17105 ( .A(n16881), .B(n16882), .Z(n16869) );
  NANDN U17106 ( .A(n16779), .B(n16778), .Z(n16783) );
  NAND U17107 ( .A(n16781), .B(n16780), .Z(n16782) );
  AND U17108 ( .A(n16783), .B(n16782), .Z(n16867) );
  NANDN U17109 ( .A(n16785), .B(n16784), .Z(n16789) );
  NANDN U17110 ( .A(n16787), .B(n16786), .Z(n16788) );
  AND U17111 ( .A(n16789), .B(n16788), .Z(n16876) );
  NANDN U17112 ( .A(n17888), .B(n16790), .Z(n16792) );
  XOR U17113 ( .A(a[118]), .B(b[11]), .Z(n16945) );
  NANDN U17114 ( .A(n18025), .B(n16945), .Z(n16791) );
  AND U17115 ( .A(n16792), .B(n16791), .Z(n16926) );
  NANDN U17116 ( .A(n18113), .B(n16793), .Z(n16795) );
  XOR U17117 ( .A(a[116]), .B(b[13]), .Z(n16948) );
  NANDN U17118 ( .A(n18229), .B(n16948), .Z(n16794) );
  AND U17119 ( .A(n16795), .B(n16794), .Z(n16925) );
  NANDN U17120 ( .A(n18487), .B(n16796), .Z(n16798) );
  XOR U17121 ( .A(a[114]), .B(b[15]), .Z(n16900) );
  NANDN U17122 ( .A(n18311), .B(n16900), .Z(n16797) );
  AND U17123 ( .A(n16798), .B(n16797), .Z(n16915) );
  NANDN U17124 ( .A(n18853), .B(n16799), .Z(n16801) );
  XOR U17125 ( .A(b[21]), .B(a[108]), .Z(n16957) );
  NANDN U17126 ( .A(n18926), .B(n16957), .Z(n16800) );
  AND U17127 ( .A(n16801), .B(n16800), .Z(n16913) );
  NANDN U17128 ( .A(n17613), .B(n16802), .Z(n16804) );
  XOR U17129 ( .A(a[120]), .B(b[9]), .Z(n16942) );
  NANDN U17130 ( .A(n17739), .B(n16942), .Z(n16803) );
  NAND U17131 ( .A(n16804), .B(n16803), .Z(n16912) );
  XNOR U17132 ( .A(n16913), .B(n16912), .Z(n16914) );
  XNOR U17133 ( .A(n16915), .B(n16914), .Z(n16924) );
  XOR U17134 ( .A(n16925), .B(n16924), .Z(n16927) );
  XOR U17135 ( .A(n16926), .B(n16927), .Z(n16888) );
  NANDN U17136 ( .A(n19005), .B(n16805), .Z(n16807) );
  XOR U17137 ( .A(b[23]), .B(a[106]), .Z(n16963) );
  NANDN U17138 ( .A(n19055), .B(n16963), .Z(n16806) );
  AND U17139 ( .A(n16807), .B(n16806), .Z(n16974) );
  NANDN U17140 ( .A(n17362), .B(n16808), .Z(n16810) );
  XOR U17141 ( .A(a[122]), .B(b[7]), .Z(n16954) );
  NANDN U17142 ( .A(n17522), .B(n16954), .Z(n16809) );
  AND U17143 ( .A(n16810), .B(n16809), .Z(n16973) );
  NANDN U17144 ( .A(n19116), .B(n16811), .Z(n16813) );
  XOR U17145 ( .A(b[25]), .B(a[104]), .Z(n16903) );
  NANDN U17146 ( .A(n19179), .B(n16903), .Z(n16812) );
  NAND U17147 ( .A(n16813), .B(n16812), .Z(n16972) );
  XOR U17148 ( .A(n16973), .B(n16972), .Z(n16975) );
  XOR U17149 ( .A(n16974), .B(n16975), .Z(n16886) );
  NANDN U17150 ( .A(n19394), .B(n16814), .Z(n16816) );
  XOR U17151 ( .A(b[29]), .B(a[100]), .Z(n16969) );
  NANDN U17152 ( .A(n19395), .B(n16969), .Z(n16815) );
  AND U17153 ( .A(n16816), .B(n16815), .Z(n16892) );
  AND U17154 ( .A(b[31]), .B(a[96]), .Z(n16891) );
  XOR U17155 ( .A(n16892), .B(n16891), .Z(n16894) );
  XNOR U17156 ( .A(n16893), .B(n16894), .Z(n16885) );
  XNOR U17157 ( .A(n16886), .B(n16885), .Z(n16887) );
  XNOR U17158 ( .A(n16888), .B(n16887), .Z(n16987) );
  NANDN U17159 ( .A(n16818), .B(n16817), .Z(n16822) );
  NANDN U17160 ( .A(n16820), .B(n16819), .Z(n16821) );
  AND U17161 ( .A(n16822), .B(n16821), .Z(n16984) );
  NANDN U17162 ( .A(n16824), .B(n16823), .Z(n16828) );
  OR U17163 ( .A(n16826), .B(n16825), .Z(n16827) );
  NAND U17164 ( .A(n16828), .B(n16827), .Z(n16985) );
  XNOR U17165 ( .A(n16984), .B(n16985), .Z(n16986) );
  XOR U17166 ( .A(n16987), .B(n16986), .Z(n16874) );
  NANDN U17167 ( .A(n16830), .B(n16829), .Z(n16834) );
  NANDN U17168 ( .A(n16832), .B(n16831), .Z(n16833) );
  NAND U17169 ( .A(n16834), .B(n16833), .Z(n16873) );
  XNOR U17170 ( .A(n16874), .B(n16873), .Z(n16875) );
  XOR U17171 ( .A(n16876), .B(n16875), .Z(n16868) );
  XOR U17172 ( .A(n16867), .B(n16868), .Z(n16870) );
  XOR U17173 ( .A(n16869), .B(n16870), .Z(n16863) );
  NANDN U17174 ( .A(n16836), .B(n16835), .Z(n16840) );
  NANDN U17175 ( .A(n16838), .B(n16837), .Z(n16839) );
  AND U17176 ( .A(n16840), .B(n16839), .Z(n16861) );
  NANDN U17177 ( .A(n16842), .B(n16841), .Z(n16846) );
  NANDN U17178 ( .A(n16844), .B(n16843), .Z(n16845) );
  NAND U17179 ( .A(n16846), .B(n16845), .Z(n16862) );
  XOR U17180 ( .A(n16861), .B(n16862), .Z(n16864) );
  XNOR U17181 ( .A(n16863), .B(n16864), .Z(n16990) );
  XNOR U17182 ( .A(n16991), .B(n16990), .Z(n16992) );
  XOR U17183 ( .A(n16993), .B(n16992), .Z(n16856) );
  NANDN U17184 ( .A(n16848), .B(n16847), .Z(n16852) );
  NAND U17185 ( .A(n16850), .B(n16849), .Z(n16851) );
  AND U17186 ( .A(n16852), .B(n16851), .Z(n16855) );
  XOR U17187 ( .A(n16856), .B(n16855), .Z(n16858) );
  XNOR U17188 ( .A(n16857), .B(n16858), .Z(n16853) );
  XOR U17189 ( .A(n16854), .B(n16853), .Z(c[224]) );
  AND U17190 ( .A(n16854), .B(n16853), .Z(n16997) );
  NANDN U17191 ( .A(n16856), .B(n16855), .Z(n16860) );
  OR U17192 ( .A(n16858), .B(n16857), .Z(n16859) );
  AND U17193 ( .A(n16860), .B(n16859), .Z(n17000) );
  NANDN U17194 ( .A(n16862), .B(n16861), .Z(n16866) );
  OR U17195 ( .A(n16864), .B(n16863), .Z(n16865) );
  AND U17196 ( .A(n16866), .B(n16865), .Z(n17137) );
  NANDN U17197 ( .A(n16868), .B(n16867), .Z(n16872) );
  OR U17198 ( .A(n16870), .B(n16869), .Z(n16871) );
  AND U17199 ( .A(n16872), .B(n16871), .Z(n17135) );
  NANDN U17200 ( .A(n16874), .B(n16873), .Z(n16878) );
  NANDN U17201 ( .A(n16876), .B(n16875), .Z(n16877) );
  AND U17202 ( .A(n16878), .B(n16877), .Z(n17129) );
  NANDN U17203 ( .A(n16880), .B(n16879), .Z(n16884) );
  OR U17204 ( .A(n16882), .B(n16881), .Z(n16883) );
  AND U17205 ( .A(n16884), .B(n16883), .Z(n17128) );
  XNOR U17206 ( .A(n17129), .B(n17128), .Z(n17130) );
  NANDN U17207 ( .A(n16886), .B(n16885), .Z(n16890) );
  NANDN U17208 ( .A(n16888), .B(n16887), .Z(n16889) );
  AND U17209 ( .A(n16890), .B(n16889), .Z(n17006) );
  NANDN U17210 ( .A(n16892), .B(n16891), .Z(n16896) );
  OR U17211 ( .A(n16894), .B(n16893), .Z(n16895) );
  AND U17212 ( .A(n16896), .B(n16895), .Z(n17049) );
  NANDN U17213 ( .A(n19237), .B(n16897), .Z(n16899) );
  XOR U17214 ( .A(b[27]), .B(a[103]), .Z(n17060) );
  NANDN U17215 ( .A(n19277), .B(n17060), .Z(n16898) );
  AND U17216 ( .A(n16899), .B(n16898), .Z(n17053) );
  NANDN U17217 ( .A(n18487), .B(n16900), .Z(n16902) );
  XOR U17218 ( .A(a[115]), .B(b[15]), .Z(n17096) );
  NANDN U17219 ( .A(n18311), .B(n17096), .Z(n16901) );
  NAND U17220 ( .A(n16902), .B(n16901), .Z(n17052) );
  XOR U17221 ( .A(b[1]), .B(n17052), .Z(n17054) );
  XOR U17222 ( .A(n17053), .B(n17054), .Z(n17047) );
  NANDN U17223 ( .A(n19116), .B(n16903), .Z(n16905) );
  XOR U17224 ( .A(b[25]), .B(a[105]), .Z(n17025) );
  NANDN U17225 ( .A(n19179), .B(n17025), .Z(n16904) );
  AND U17226 ( .A(n16905), .B(n16904), .Z(n17036) );
  NANDN U17227 ( .A(n17067), .B(n16906), .Z(n16908) );
  XOR U17228 ( .A(a[127]), .B(b[3]), .Z(n17066) );
  NANDN U17229 ( .A(n17068), .B(n17066), .Z(n16907) );
  AND U17230 ( .A(n16908), .B(n16907), .Z(n17035) );
  NANDN U17231 ( .A(n18514), .B(n16909), .Z(n16911) );
  XOR U17232 ( .A(b[17]), .B(a[113]), .Z(n17063) );
  NANDN U17233 ( .A(n18585), .B(n17063), .Z(n16910) );
  NAND U17234 ( .A(n16911), .B(n16910), .Z(n17034) );
  XOR U17235 ( .A(n17035), .B(n17034), .Z(n17037) );
  XNOR U17236 ( .A(n17036), .B(n17037), .Z(n17046) );
  XNOR U17237 ( .A(n17047), .B(n17046), .Z(n17048) );
  XOR U17238 ( .A(n17049), .B(n17048), .Z(n17005) );
  NANDN U17239 ( .A(n16913), .B(n16912), .Z(n16917) );
  NANDN U17240 ( .A(n16915), .B(n16914), .Z(n16916) );
  AND U17241 ( .A(n16917), .B(n16916), .Z(n17116) );
  NANDN U17242 ( .A(n16919), .B(n16918), .Z(n16923) );
  NANDN U17243 ( .A(n16921), .B(n16920), .Z(n16922) );
  NAND U17244 ( .A(n16923), .B(n16922), .Z(n17117) );
  XNOR U17245 ( .A(n17116), .B(n17117), .Z(n17119) );
  NANDN U17246 ( .A(n16925), .B(n16924), .Z(n16929) );
  OR U17247 ( .A(n16927), .B(n16926), .Z(n16928) );
  AND U17248 ( .A(n16929), .B(n16928), .Z(n17118) );
  XNOR U17249 ( .A(n17119), .B(n17118), .Z(n17004) );
  XOR U17250 ( .A(n17005), .B(n17004), .Z(n17007) );
  XNOR U17251 ( .A(n17006), .B(n17007), .Z(n17124) );
  NANDN U17252 ( .A(n16931), .B(n16930), .Z(n16935) );
  NANDN U17253 ( .A(n16933), .B(n16932), .Z(n16934) );
  AND U17254 ( .A(n16935), .B(n16934), .Z(n17122) );
  NANDN U17255 ( .A(n16937), .B(n16936), .Z(n16941) );
  OR U17256 ( .A(n16939), .B(n16938), .Z(n16940) );
  AND U17257 ( .A(n16941), .B(n16940), .Z(n17085) );
  NANDN U17258 ( .A(n17613), .B(n16942), .Z(n16944) );
  XOR U17259 ( .A(a[121]), .B(b[9]), .Z(n17010) );
  NANDN U17260 ( .A(n17739), .B(n17010), .Z(n16943) );
  AND U17261 ( .A(n16944), .B(n16943), .Z(n17043) );
  NANDN U17262 ( .A(n17888), .B(n16945), .Z(n16947) );
  XOR U17263 ( .A(a[119]), .B(b[11]), .Z(n17022) );
  NANDN U17264 ( .A(n18025), .B(n17022), .Z(n16946) );
  AND U17265 ( .A(n16947), .B(n16946), .Z(n17041) );
  NANDN U17266 ( .A(n18113), .B(n16948), .Z(n16950) );
  XOR U17267 ( .A(a[117]), .B(b[13]), .Z(n17019) );
  NANDN U17268 ( .A(n18229), .B(n17019), .Z(n16949) );
  AND U17269 ( .A(n16950), .B(n16949), .Z(n17031) );
  NANDN U17270 ( .A(n18673), .B(n16951), .Z(n16953) );
  XOR U17271 ( .A(b[19]), .B(a[111]), .Z(n17075) );
  NANDN U17272 ( .A(n18758), .B(n17075), .Z(n16952) );
  AND U17273 ( .A(n16953), .B(n16952), .Z(n17029) );
  NANDN U17274 ( .A(n17362), .B(n16954), .Z(n16956) );
  XOR U17275 ( .A(a[123]), .B(b[7]), .Z(n17013) );
  NANDN U17276 ( .A(n17522), .B(n17013), .Z(n16955) );
  NAND U17277 ( .A(n16956), .B(n16955), .Z(n17028) );
  XNOR U17278 ( .A(n17029), .B(n17028), .Z(n17030) );
  XNOR U17279 ( .A(n17031), .B(n17030), .Z(n17040) );
  XNOR U17280 ( .A(n17041), .B(n17040), .Z(n17042) );
  XOR U17281 ( .A(n17043), .B(n17042), .Z(n17080) );
  NANDN U17282 ( .A(n18853), .B(n16957), .Z(n16959) );
  XOR U17283 ( .A(b[21]), .B(a[109]), .Z(n17016) );
  NANDN U17284 ( .A(n18926), .B(n17016), .Z(n16958) );
  AND U17285 ( .A(n16959), .B(n16958), .Z(n17113) );
  NANDN U17286 ( .A(n17072), .B(n16960), .Z(n16962) );
  XOR U17287 ( .A(a[125]), .B(b[5]), .Z(n17071) );
  NANDN U17288 ( .A(n17223), .B(n17071), .Z(n16961) );
  AND U17289 ( .A(n16962), .B(n16961), .Z(n17111) );
  NANDN U17290 ( .A(n19005), .B(n16963), .Z(n16965) );
  XOR U17291 ( .A(b[23]), .B(a[107]), .Z(n17057) );
  NANDN U17292 ( .A(n19055), .B(n17057), .Z(n16964) );
  NAND U17293 ( .A(n16965), .B(n16964), .Z(n17110) );
  XNOR U17294 ( .A(n17111), .B(n17110), .Z(n17112) );
  XOR U17295 ( .A(n17113), .B(n17112), .Z(n17079) );
  NANDN U17296 ( .A(n19425), .B(n16966), .Z(n16968) );
  XOR U17297 ( .A(b[31]), .B(a[99]), .Z(n17102) );
  NANDN U17298 ( .A(n19426), .B(n17102), .Z(n16967) );
  AND U17299 ( .A(n16968), .B(n16967), .Z(n17107) );
  NAND U17300 ( .A(b[31]), .B(a[97]), .Z(n17337) );
  NANDN U17301 ( .A(n19394), .B(n16969), .Z(n16971) );
  XOR U17302 ( .A(b[29]), .B(a[101]), .Z(n17099) );
  NANDN U17303 ( .A(n19395), .B(n17099), .Z(n16970) );
  NAND U17304 ( .A(n16971), .B(n16970), .Z(n17105) );
  XOR U17305 ( .A(n17337), .B(n17105), .Z(n17106) );
  XOR U17306 ( .A(n17107), .B(n17106), .Z(n17078) );
  XNOR U17307 ( .A(n17079), .B(n17078), .Z(n17081) );
  NANDN U17308 ( .A(n16973), .B(n16972), .Z(n16977) );
  OR U17309 ( .A(n16975), .B(n16974), .Z(n16976) );
  AND U17310 ( .A(n16977), .B(n16976), .Z(n17091) );
  NANDN U17311 ( .A(n16979), .B(n16978), .Z(n16983) );
  NANDN U17312 ( .A(n16981), .B(n16980), .Z(n16982) );
  NAND U17313 ( .A(n16983), .B(n16982), .Z(n17090) );
  XNOR U17314 ( .A(n17091), .B(n17090), .Z(n17092) );
  XOR U17315 ( .A(n17093), .B(n17092), .Z(n17084) );
  XNOR U17316 ( .A(n17085), .B(n17084), .Z(n17086) );
  NANDN U17317 ( .A(n16985), .B(n16984), .Z(n16989) );
  NAND U17318 ( .A(n16987), .B(n16986), .Z(n16988) );
  NAND U17319 ( .A(n16989), .B(n16988), .Z(n17087) );
  XOR U17320 ( .A(n17086), .B(n17087), .Z(n17123) );
  XOR U17321 ( .A(n17122), .B(n17123), .Z(n17125) );
  XOR U17322 ( .A(n17124), .B(n17125), .Z(n17131) );
  XNOR U17323 ( .A(n17130), .B(n17131), .Z(n17134) );
  XNOR U17324 ( .A(n17135), .B(n17134), .Z(n17136) );
  XOR U17325 ( .A(n17137), .B(n17136), .Z(n16999) );
  NANDN U17326 ( .A(n16991), .B(n16990), .Z(n16995) );
  NAND U17327 ( .A(n16993), .B(n16992), .Z(n16994) );
  AND U17328 ( .A(n16995), .B(n16994), .Z(n16998) );
  XOR U17329 ( .A(n16999), .B(n16998), .Z(n17001) );
  XNOR U17330 ( .A(n17000), .B(n17001), .Z(n16996) );
  XOR U17331 ( .A(n16997), .B(n16996), .Z(c[225]) );
  AND U17332 ( .A(n16997), .B(n16996), .Z(n17141) );
  NANDN U17333 ( .A(n16999), .B(n16998), .Z(n17003) );
  OR U17334 ( .A(n17001), .B(n17000), .Z(n17002) );
  AND U17335 ( .A(n17003), .B(n17002), .Z(n17144) );
  NANDN U17336 ( .A(n17005), .B(n17004), .Z(n17009) );
  NANDN U17337 ( .A(n17007), .B(n17006), .Z(n17008) );
  AND U17338 ( .A(n17009), .B(n17008), .Z(n17272) );
  NANDN U17339 ( .A(n17613), .B(n17010), .Z(n17012) );
  XOR U17340 ( .A(a[122]), .B(b[9]), .Z(n17236) );
  NANDN U17341 ( .A(n17739), .B(n17236), .Z(n17011) );
  AND U17342 ( .A(n17012), .B(n17011), .Z(n17195) );
  NANDN U17343 ( .A(n17362), .B(n17013), .Z(n17015) );
  XOR U17344 ( .A(a[124]), .B(b[7]), .Z(n17248) );
  NANDN U17345 ( .A(n17522), .B(n17248), .Z(n17014) );
  AND U17346 ( .A(n17015), .B(n17014), .Z(n17194) );
  NANDN U17347 ( .A(n18853), .B(n17016), .Z(n17018) );
  XOR U17348 ( .A(b[21]), .B(a[110]), .Z(n17254) );
  NANDN U17349 ( .A(n18926), .B(n17254), .Z(n17017) );
  NAND U17350 ( .A(n17018), .B(n17017), .Z(n17193) );
  XOR U17351 ( .A(n17194), .B(n17193), .Z(n17196) );
  XOR U17352 ( .A(n17195), .B(n17196), .Z(n17206) );
  NANDN U17353 ( .A(n18113), .B(n17019), .Z(n17021) );
  XOR U17354 ( .A(a[118]), .B(b[13]), .Z(n17178) );
  NANDN U17355 ( .A(n18229), .B(n17178), .Z(n17020) );
  AND U17356 ( .A(n17021), .B(n17020), .Z(n17219) );
  NANDN U17357 ( .A(n17888), .B(n17022), .Z(n17024) );
  XOR U17358 ( .A(a[120]), .B(b[11]), .Z(n17245) );
  NANDN U17359 ( .A(n18025), .B(n17245), .Z(n17023) );
  AND U17360 ( .A(n17024), .B(n17023), .Z(n17218) );
  NANDN U17361 ( .A(n19116), .B(n17025), .Z(n17027) );
  XOR U17362 ( .A(b[25]), .B(a[106]), .Z(n17239) );
  NANDN U17363 ( .A(n19179), .B(n17239), .Z(n17026) );
  NAND U17364 ( .A(n17027), .B(n17026), .Z(n17217) );
  XOR U17365 ( .A(n17218), .B(n17217), .Z(n17220) );
  XNOR U17366 ( .A(n17219), .B(n17220), .Z(n17205) );
  XNOR U17367 ( .A(n17206), .B(n17205), .Z(n17207) );
  NANDN U17368 ( .A(n17029), .B(n17028), .Z(n17033) );
  NANDN U17369 ( .A(n17031), .B(n17030), .Z(n17032) );
  NAND U17370 ( .A(n17033), .B(n17032), .Z(n17208) );
  XNOR U17371 ( .A(n17207), .B(n17208), .Z(n17263) );
  NANDN U17372 ( .A(n17035), .B(n17034), .Z(n17039) );
  OR U17373 ( .A(n17037), .B(n17036), .Z(n17038) );
  NAND U17374 ( .A(n17039), .B(n17038), .Z(n17264) );
  XNOR U17375 ( .A(n17263), .B(n17264), .Z(n17266) );
  NANDN U17376 ( .A(n17041), .B(n17040), .Z(n17045) );
  NANDN U17377 ( .A(n17043), .B(n17042), .Z(n17044) );
  AND U17378 ( .A(n17045), .B(n17044), .Z(n17265) );
  XOR U17379 ( .A(n17266), .B(n17265), .Z(n17270) );
  NANDN U17380 ( .A(n17047), .B(n17046), .Z(n17051) );
  NAND U17381 ( .A(n17049), .B(n17048), .Z(n17050) );
  AND U17382 ( .A(n17051), .B(n17050), .Z(n17162) );
  NANDN U17383 ( .A(b[1]), .B(n17052), .Z(n17056) );
  OR U17384 ( .A(n17054), .B(n17053), .Z(n17055) );
  AND U17385 ( .A(n17056), .B(n17055), .Z(n17214) );
  NANDN U17386 ( .A(n19005), .B(n17057), .Z(n17059) );
  XOR U17387 ( .A(b[23]), .B(a[108]), .Z(n17230) );
  NANDN U17388 ( .A(n19055), .B(n17230), .Z(n17058) );
  AND U17389 ( .A(n17059), .B(n17058), .Z(n17189) );
  NANDN U17390 ( .A(n19237), .B(n17060), .Z(n17062) );
  XOR U17391 ( .A(b[27]), .B(a[104]), .Z(n17242) );
  NANDN U17392 ( .A(n19277), .B(n17242), .Z(n17061) );
  AND U17393 ( .A(n17062), .B(n17061), .Z(n17188) );
  NANDN U17394 ( .A(n18514), .B(n17063), .Z(n17065) );
  XOR U17395 ( .A(b[17]), .B(a[114]), .Z(n17175) );
  NANDN U17396 ( .A(n18585), .B(n17175), .Z(n17064) );
  NAND U17397 ( .A(n17065), .B(n17064), .Z(n17187) );
  XOR U17398 ( .A(n17188), .B(n17187), .Z(n17190) );
  XOR U17399 ( .A(n17189), .B(n17190), .Z(n17212) );
  NANDN U17400 ( .A(n17067), .B(n17066), .Z(n17070) );
  NANDN U17401 ( .A(n17068), .B(b[3]), .Z(n17069) );
  AND U17402 ( .A(n17070), .B(n17069), .Z(n17182) );
  AND U17403 ( .A(b[31]), .B(a[98]), .Z(n17181) );
  XNOR U17404 ( .A(n17182), .B(n17181), .Z(n17183) );
  XOR U17405 ( .A(n17337), .B(n17183), .Z(n17202) );
  NANDN U17406 ( .A(n17072), .B(n17071), .Z(n17074) );
  XOR U17407 ( .A(a[126]), .B(b[5]), .Z(n17224) );
  NANDN U17408 ( .A(n17223), .B(n17224), .Z(n17073) );
  AND U17409 ( .A(n17074), .B(n17073), .Z(n17200) );
  NANDN U17410 ( .A(n18673), .B(n17075), .Z(n17077) );
  XOR U17411 ( .A(b[19]), .B(a[112]), .Z(n17227) );
  NANDN U17412 ( .A(n18758), .B(n17227), .Z(n17076) );
  NAND U17413 ( .A(n17077), .B(n17076), .Z(n17199) );
  XNOR U17414 ( .A(n17200), .B(n17199), .Z(n17201) );
  XNOR U17415 ( .A(n17202), .B(n17201), .Z(n17211) );
  XNOR U17416 ( .A(n17212), .B(n17211), .Z(n17213) );
  XOR U17417 ( .A(n17214), .B(n17213), .Z(n17161) );
  NAND U17418 ( .A(n17079), .B(n17078), .Z(n17083) );
  NANDN U17419 ( .A(n17081), .B(n17080), .Z(n17082) );
  AND U17420 ( .A(n17083), .B(n17082), .Z(n17160) );
  XOR U17421 ( .A(n17161), .B(n17160), .Z(n17163) );
  XNOR U17422 ( .A(n17162), .B(n17163), .Z(n17269) );
  XNOR U17423 ( .A(n17270), .B(n17269), .Z(n17271) );
  XNOR U17424 ( .A(n17272), .B(n17271), .Z(n17278) );
  NANDN U17425 ( .A(n17085), .B(n17084), .Z(n17089) );
  NANDN U17426 ( .A(n17087), .B(n17086), .Z(n17088) );
  AND U17427 ( .A(n17089), .B(n17088), .Z(n17276) );
  NANDN U17428 ( .A(n17091), .B(n17090), .Z(n17095) );
  NAND U17429 ( .A(n17093), .B(n17092), .Z(n17094) );
  AND U17430 ( .A(n17095), .B(n17094), .Z(n17157) );
  NANDN U17431 ( .A(n18487), .B(n17096), .Z(n17098) );
  XOR U17432 ( .A(a[116]), .B(b[15]), .Z(n17172) );
  NANDN U17433 ( .A(n18311), .B(n17172), .Z(n17097) );
  AND U17434 ( .A(n17098), .B(n17097), .Z(n17259) );
  NANDN U17435 ( .A(n19394), .B(n17099), .Z(n17101) );
  XOR U17436 ( .A(b[29]), .B(a[102]), .Z(n17233) );
  NANDN U17437 ( .A(n19395), .B(n17233), .Z(n17100) );
  AND U17438 ( .A(n17101), .B(n17100), .Z(n17258) );
  NANDN U17439 ( .A(n19425), .B(n17102), .Z(n17104) );
  XOR U17440 ( .A(b[31]), .B(a[100]), .Z(n17251) );
  NANDN U17441 ( .A(n19426), .B(n17251), .Z(n17103) );
  NAND U17442 ( .A(n17104), .B(n17103), .Z(n17257) );
  XOR U17443 ( .A(n17258), .B(n17257), .Z(n17260) );
  XOR U17444 ( .A(n17259), .B(n17260), .Z(n17167) );
  IV U17445 ( .A(n17337), .Z(n17184) );
  NANDN U17446 ( .A(n17184), .B(n17105), .Z(n17109) );
  NANDN U17447 ( .A(n17107), .B(n17106), .Z(n17108) );
  AND U17448 ( .A(n17109), .B(n17108), .Z(n17166) );
  XNOR U17449 ( .A(n17167), .B(n17166), .Z(n17169) );
  NANDN U17450 ( .A(n17111), .B(n17110), .Z(n17115) );
  NANDN U17451 ( .A(n17113), .B(n17112), .Z(n17114) );
  AND U17452 ( .A(n17115), .B(n17114), .Z(n17168) );
  XOR U17453 ( .A(n17169), .B(n17168), .Z(n17155) );
  NANDN U17454 ( .A(n17117), .B(n17116), .Z(n17121) );
  NAND U17455 ( .A(n17119), .B(n17118), .Z(n17120) );
  AND U17456 ( .A(n17121), .B(n17120), .Z(n17154) );
  XNOR U17457 ( .A(n17155), .B(n17154), .Z(n17156) );
  XNOR U17458 ( .A(n17157), .B(n17156), .Z(n17275) );
  XNOR U17459 ( .A(n17276), .B(n17275), .Z(n17277) );
  XOR U17460 ( .A(n17278), .B(n17277), .Z(n17149) );
  NANDN U17461 ( .A(n17123), .B(n17122), .Z(n17127) );
  NANDN U17462 ( .A(n17125), .B(n17124), .Z(n17126) );
  AND U17463 ( .A(n17127), .B(n17126), .Z(n17148) );
  XNOR U17464 ( .A(n17149), .B(n17148), .Z(n17150) );
  NANDN U17465 ( .A(n17129), .B(n17128), .Z(n17133) );
  NANDN U17466 ( .A(n17131), .B(n17130), .Z(n17132) );
  NAND U17467 ( .A(n17133), .B(n17132), .Z(n17151) );
  XNOR U17468 ( .A(n17150), .B(n17151), .Z(n17142) );
  NANDN U17469 ( .A(n17135), .B(n17134), .Z(n17139) );
  NAND U17470 ( .A(n17137), .B(n17136), .Z(n17138) );
  NAND U17471 ( .A(n17139), .B(n17138), .Z(n17143) );
  XOR U17472 ( .A(n17142), .B(n17143), .Z(n17145) );
  XNOR U17473 ( .A(n17144), .B(n17145), .Z(n17140) );
  XOR U17474 ( .A(n17141), .B(n17140), .Z(c[226]) );
  AND U17475 ( .A(n17141), .B(n17140), .Z(n17282) );
  NANDN U17476 ( .A(n17143), .B(n17142), .Z(n17147) );
  OR U17477 ( .A(n17145), .B(n17144), .Z(n17146) );
  AND U17478 ( .A(n17147), .B(n17146), .Z(n17285) );
  NANDN U17479 ( .A(n17149), .B(n17148), .Z(n17153) );
  NANDN U17480 ( .A(n17151), .B(n17150), .Z(n17152) );
  AND U17481 ( .A(n17153), .B(n17152), .Z(n17284) );
  NANDN U17482 ( .A(n17155), .B(n17154), .Z(n17159) );
  NANDN U17483 ( .A(n17157), .B(n17156), .Z(n17158) );
  AND U17484 ( .A(n17159), .B(n17158), .Z(n17296) );
  NANDN U17485 ( .A(n17161), .B(n17160), .Z(n17165) );
  NANDN U17486 ( .A(n17163), .B(n17162), .Z(n17164) );
  NAND U17487 ( .A(n17165), .B(n17164), .Z(n17295) );
  XNOR U17488 ( .A(n17296), .B(n17295), .Z(n17298) );
  NANDN U17489 ( .A(n17167), .B(n17166), .Z(n17171) );
  NAND U17490 ( .A(n17169), .B(n17168), .Z(n17170) );
  AND U17491 ( .A(n17171), .B(n17170), .Z(n17402) );
  NANDN U17492 ( .A(n18487), .B(n17172), .Z(n17174) );
  XOR U17493 ( .A(a[117]), .B(b[15]), .Z(n17325) );
  NANDN U17494 ( .A(n18311), .B(n17325), .Z(n17173) );
  AND U17495 ( .A(n17174), .B(n17173), .Z(n17342) );
  NANDN U17496 ( .A(n18514), .B(n17175), .Z(n17177) );
  XOR U17497 ( .A(b[17]), .B(a[115]), .Z(n17328) );
  NANDN U17498 ( .A(n18585), .B(n17328), .Z(n17176) );
  AND U17499 ( .A(n17177), .B(n17176), .Z(n17341) );
  NANDN U17500 ( .A(n18113), .B(n17178), .Z(n17180) );
  XOR U17501 ( .A(a[119]), .B(b[13]), .Z(n17331) );
  NANDN U17502 ( .A(n18229), .B(n17331), .Z(n17179) );
  NAND U17503 ( .A(n17180), .B(n17179), .Z(n17340) );
  XOR U17504 ( .A(n17341), .B(n17340), .Z(n17343) );
  XOR U17505 ( .A(n17342), .B(n17343), .Z(n17347) );
  NANDN U17506 ( .A(n17182), .B(n17181), .Z(n17186) );
  NANDN U17507 ( .A(n17184), .B(n17183), .Z(n17185) );
  AND U17508 ( .A(n17186), .B(n17185), .Z(n17346) );
  XNOR U17509 ( .A(n17347), .B(n17346), .Z(n17349) );
  NANDN U17510 ( .A(n17188), .B(n17187), .Z(n17192) );
  OR U17511 ( .A(n17190), .B(n17189), .Z(n17191) );
  AND U17512 ( .A(n17192), .B(n17191), .Z(n17348) );
  XOR U17513 ( .A(n17349), .B(n17348), .Z(n17408) );
  NANDN U17514 ( .A(n17194), .B(n17193), .Z(n17198) );
  OR U17515 ( .A(n17196), .B(n17195), .Z(n17197) );
  AND U17516 ( .A(n17198), .B(n17197), .Z(n17407) );
  NANDN U17517 ( .A(n17200), .B(n17199), .Z(n17204) );
  NAND U17518 ( .A(n17202), .B(n17201), .Z(n17203) );
  NAND U17519 ( .A(n17204), .B(n17203), .Z(n17406) );
  XOR U17520 ( .A(n17407), .B(n17406), .Z(n17409) );
  XOR U17521 ( .A(n17408), .B(n17409), .Z(n17401) );
  NANDN U17522 ( .A(n17206), .B(n17205), .Z(n17210) );
  NANDN U17523 ( .A(n17208), .B(n17207), .Z(n17209) );
  NAND U17524 ( .A(n17210), .B(n17209), .Z(n17400) );
  XOR U17525 ( .A(n17401), .B(n17400), .Z(n17403) );
  XOR U17526 ( .A(n17402), .B(n17403), .Z(n17304) );
  NANDN U17527 ( .A(n17212), .B(n17211), .Z(n17216) );
  NAND U17528 ( .A(n17214), .B(n17213), .Z(n17215) );
  AND U17529 ( .A(n17216), .B(n17215), .Z(n17309) );
  NANDN U17530 ( .A(n17218), .B(n17217), .Z(n17222) );
  OR U17531 ( .A(n17220), .B(n17219), .Z(n17221) );
  AND U17532 ( .A(n17222), .B(n17221), .Z(n17414) );
  XNOR U17533 ( .A(a[127]), .B(b[5]), .Z(n17389) );
  OR U17534 ( .A(n17389), .B(n17223), .Z(n17226) );
  NAND U17535 ( .A(n17390), .B(n17224), .Z(n17225) );
  AND U17536 ( .A(n17226), .B(n17225), .Z(n17320) );
  NANDN U17537 ( .A(n18673), .B(n17227), .Z(n17229) );
  XOR U17538 ( .A(b[19]), .B(a[113]), .Z(n17368) );
  NANDN U17539 ( .A(n18758), .B(n17368), .Z(n17228) );
  NAND U17540 ( .A(n17229), .B(n17228), .Z(n17319) );
  XNOR U17541 ( .A(n17320), .B(n17319), .Z(n17321) );
  AND U17542 ( .A(b[31]), .B(a[99]), .Z(n17334) );
  XNOR U17543 ( .A(n17334), .B(n17335), .Z(n17336) );
  XNOR U17544 ( .A(n17337), .B(n17336), .Z(n17322) );
  XOR U17545 ( .A(n17321), .B(n17322), .Z(n17412) );
  NANDN U17546 ( .A(n19005), .B(n17230), .Z(n17232) );
  XOR U17547 ( .A(b[23]), .B(a[109]), .Z(n17352) );
  NANDN U17548 ( .A(n19055), .B(n17352), .Z(n17231) );
  AND U17549 ( .A(n17232), .B(n17231), .Z(n17397) );
  NANDN U17550 ( .A(n19394), .B(n17233), .Z(n17235) );
  XOR U17551 ( .A(b[29]), .B(a[103]), .Z(n17365) );
  NANDN U17552 ( .A(n19395), .B(n17365), .Z(n17234) );
  AND U17553 ( .A(n17235), .B(n17234), .Z(n17395) );
  NANDN U17554 ( .A(n17613), .B(n17236), .Z(n17238) );
  XOR U17555 ( .A(a[123]), .B(b[9]), .Z(n17380) );
  NANDN U17556 ( .A(n17739), .B(n17380), .Z(n17237) );
  NAND U17557 ( .A(n17238), .B(n17237), .Z(n17394) );
  XNOR U17558 ( .A(n17395), .B(n17394), .Z(n17396) );
  XOR U17559 ( .A(n17397), .B(n17396), .Z(n17413) );
  XOR U17560 ( .A(n17412), .B(n17413), .Z(n17415) );
  XOR U17561 ( .A(n17414), .B(n17415), .Z(n17308) );
  NANDN U17562 ( .A(n19116), .B(n17239), .Z(n17241) );
  XOR U17563 ( .A(b[25]), .B(a[107]), .Z(n17355) );
  NANDN U17564 ( .A(n19179), .B(n17355), .Z(n17240) );
  AND U17565 ( .A(n17241), .B(n17240), .Z(n17373) );
  NANDN U17566 ( .A(n19237), .B(n17242), .Z(n17244) );
  XOR U17567 ( .A(b[27]), .B(a[105]), .Z(n17377) );
  NANDN U17568 ( .A(n19277), .B(n17377), .Z(n17243) );
  AND U17569 ( .A(n17244), .B(n17243), .Z(n17372) );
  NANDN U17570 ( .A(n17888), .B(n17245), .Z(n17247) );
  XOR U17571 ( .A(a[121]), .B(b[11]), .Z(n17358) );
  NANDN U17572 ( .A(n18025), .B(n17358), .Z(n17246) );
  NAND U17573 ( .A(n17247), .B(n17246), .Z(n17371) );
  XOR U17574 ( .A(n17372), .B(n17371), .Z(n17374) );
  XOR U17575 ( .A(n17373), .B(n17374), .Z(n17419) );
  NANDN U17576 ( .A(n17362), .B(n17248), .Z(n17250) );
  XOR U17577 ( .A(a[125]), .B(b[7]), .Z(n17361) );
  NANDN U17578 ( .A(n17522), .B(n17361), .Z(n17249) );
  AND U17579 ( .A(n17250), .B(n17249), .Z(n17315) );
  NANDN U17580 ( .A(n19425), .B(n17251), .Z(n17253) );
  XOR U17581 ( .A(b[31]), .B(a[101]), .Z(n17386) );
  NANDN U17582 ( .A(n19426), .B(n17386), .Z(n17252) );
  AND U17583 ( .A(n17253), .B(n17252), .Z(n17314) );
  NANDN U17584 ( .A(n18853), .B(n17254), .Z(n17256) );
  XOR U17585 ( .A(b[21]), .B(a[111]), .Z(n17383) );
  NANDN U17586 ( .A(n18926), .B(n17383), .Z(n17255) );
  NAND U17587 ( .A(n17256), .B(n17255), .Z(n17313) );
  XOR U17588 ( .A(n17314), .B(n17313), .Z(n17316) );
  XNOR U17589 ( .A(n17315), .B(n17316), .Z(n17418) );
  XNOR U17590 ( .A(n17419), .B(n17418), .Z(n17420) );
  NANDN U17591 ( .A(n17258), .B(n17257), .Z(n17262) );
  OR U17592 ( .A(n17260), .B(n17259), .Z(n17261) );
  NAND U17593 ( .A(n17262), .B(n17261), .Z(n17421) );
  XNOR U17594 ( .A(n17420), .B(n17421), .Z(n17307) );
  XOR U17595 ( .A(n17308), .B(n17307), .Z(n17310) );
  XOR U17596 ( .A(n17309), .B(n17310), .Z(n17302) );
  NANDN U17597 ( .A(n17264), .B(n17263), .Z(n17268) );
  NAND U17598 ( .A(n17266), .B(n17265), .Z(n17267) );
  AND U17599 ( .A(n17268), .B(n17267), .Z(n17301) );
  XNOR U17600 ( .A(n17302), .B(n17301), .Z(n17303) );
  XNOR U17601 ( .A(n17304), .B(n17303), .Z(n17297) );
  XOR U17602 ( .A(n17298), .B(n17297), .Z(n17292) );
  NANDN U17603 ( .A(n17270), .B(n17269), .Z(n17274) );
  NANDN U17604 ( .A(n17272), .B(n17271), .Z(n17273) );
  AND U17605 ( .A(n17274), .B(n17273), .Z(n17289) );
  NANDN U17606 ( .A(n17276), .B(n17275), .Z(n17280) );
  NAND U17607 ( .A(n17278), .B(n17277), .Z(n17279) );
  NAND U17608 ( .A(n17280), .B(n17279), .Z(n17290) );
  XNOR U17609 ( .A(n17289), .B(n17290), .Z(n17291) );
  XNOR U17610 ( .A(n17292), .B(n17291), .Z(n17283) );
  XOR U17611 ( .A(n17284), .B(n17283), .Z(n17286) );
  XNOR U17612 ( .A(n17285), .B(n17286), .Z(n17281) );
  XOR U17613 ( .A(n17282), .B(n17281), .Z(c[227]) );
  AND U17614 ( .A(n17282), .B(n17281), .Z(n17425) );
  NANDN U17615 ( .A(n17284), .B(n17283), .Z(n17288) );
  OR U17616 ( .A(n17286), .B(n17285), .Z(n17287) );
  AND U17617 ( .A(n17288), .B(n17287), .Z(n17428) );
  NANDN U17618 ( .A(n17290), .B(n17289), .Z(n17294) );
  NANDN U17619 ( .A(n17292), .B(n17291), .Z(n17293) );
  AND U17620 ( .A(n17294), .B(n17293), .Z(n17427) );
  NANDN U17621 ( .A(n17296), .B(n17295), .Z(n17300) );
  NAND U17622 ( .A(n17298), .B(n17297), .Z(n17299) );
  AND U17623 ( .A(n17300), .B(n17299), .Z(n17434) );
  NANDN U17624 ( .A(n17302), .B(n17301), .Z(n17306) );
  NANDN U17625 ( .A(n17304), .B(n17303), .Z(n17305) );
  AND U17626 ( .A(n17306), .B(n17305), .Z(n17432) );
  NANDN U17627 ( .A(n17308), .B(n17307), .Z(n17312) );
  OR U17628 ( .A(n17310), .B(n17309), .Z(n17311) );
  AND U17629 ( .A(n17312), .B(n17311), .Z(n17441) );
  NANDN U17630 ( .A(n17314), .B(n17313), .Z(n17318) );
  OR U17631 ( .A(n17316), .B(n17315), .Z(n17317) );
  AND U17632 ( .A(n17318), .B(n17317), .Z(n17445) );
  NANDN U17633 ( .A(n17320), .B(n17319), .Z(n17324) );
  NAND U17634 ( .A(n17322), .B(n17321), .Z(n17323) );
  NAND U17635 ( .A(n17324), .B(n17323), .Z(n17444) );
  XNOR U17636 ( .A(n17445), .B(n17444), .Z(n17447) );
  NANDN U17637 ( .A(n18487), .B(n17325), .Z(n17327) );
  XOR U17638 ( .A(a[118]), .B(b[15]), .Z(n17529) );
  NANDN U17639 ( .A(n18311), .B(n17529), .Z(n17326) );
  AND U17640 ( .A(n17327), .B(n17326), .Z(n17483) );
  NANDN U17641 ( .A(n18514), .B(n17328), .Z(n17330) );
  XOR U17642 ( .A(a[116]), .B(b[17]), .Z(n17535) );
  NANDN U17643 ( .A(n18585), .B(n17535), .Z(n17329) );
  AND U17644 ( .A(n17330), .B(n17329), .Z(n17481) );
  NANDN U17645 ( .A(n18113), .B(n17331), .Z(n17333) );
  XOR U17646 ( .A(a[120]), .B(b[13]), .Z(n17532) );
  NANDN U17647 ( .A(n18229), .B(n17532), .Z(n17332) );
  NAND U17648 ( .A(n17333), .B(n17332), .Z(n17480) );
  XNOR U17649 ( .A(n17481), .B(n17480), .Z(n17482) );
  XNOR U17650 ( .A(n17483), .B(n17482), .Z(n17475) );
  NANDN U17651 ( .A(n17335), .B(n17334), .Z(n17339) );
  NANDN U17652 ( .A(n17337), .B(n17336), .Z(n17338) );
  NAND U17653 ( .A(n17339), .B(n17338), .Z(n17474) );
  XOR U17654 ( .A(n17475), .B(n17474), .Z(n17477) );
  NANDN U17655 ( .A(n17341), .B(n17340), .Z(n17345) );
  OR U17656 ( .A(n17343), .B(n17342), .Z(n17344) );
  NAND U17657 ( .A(n17345), .B(n17344), .Z(n17476) );
  XOR U17658 ( .A(n17477), .B(n17476), .Z(n17446) );
  XOR U17659 ( .A(n17447), .B(n17446), .Z(n17439) );
  NANDN U17660 ( .A(n17347), .B(n17346), .Z(n17351) );
  NAND U17661 ( .A(n17349), .B(n17348), .Z(n17350) );
  AND U17662 ( .A(n17351), .B(n17350), .Z(n17471) );
  NANDN U17663 ( .A(n19005), .B(n17352), .Z(n17354) );
  XOR U17664 ( .A(b[23]), .B(a[110]), .Z(n17504) );
  NANDN U17665 ( .A(n19055), .B(n17504), .Z(n17353) );
  AND U17666 ( .A(n17354), .B(n17353), .Z(n17546) );
  NANDN U17667 ( .A(n19116), .B(n17355), .Z(n17357) );
  XOR U17668 ( .A(b[25]), .B(a[108]), .Z(n17538) );
  NANDN U17669 ( .A(n19179), .B(n17538), .Z(n17356) );
  AND U17670 ( .A(n17357), .B(n17356), .Z(n17545) );
  NANDN U17671 ( .A(n17888), .B(n17358), .Z(n17360) );
  XOR U17672 ( .A(a[122]), .B(b[11]), .Z(n17541) );
  NANDN U17673 ( .A(n18025), .B(n17541), .Z(n17359) );
  NAND U17674 ( .A(n17360), .B(n17359), .Z(n17544) );
  XOR U17675 ( .A(n17545), .B(n17544), .Z(n17547) );
  XOR U17676 ( .A(n17546), .B(n17547), .Z(n17457) );
  NANDN U17677 ( .A(n17362), .B(n17361), .Z(n17364) );
  XOR U17678 ( .A(a[126]), .B(b[7]), .Z(n17523) );
  NANDN U17679 ( .A(n17522), .B(n17523), .Z(n17363) );
  AND U17680 ( .A(n17364), .B(n17363), .Z(n17515) );
  NANDN U17681 ( .A(n19394), .B(n17365), .Z(n17367) );
  XOR U17682 ( .A(b[29]), .B(a[104]), .Z(n17519) );
  NANDN U17683 ( .A(n19395), .B(n17519), .Z(n17366) );
  AND U17684 ( .A(n17367), .B(n17366), .Z(n17514) );
  NANDN U17685 ( .A(n18673), .B(n17368), .Z(n17370) );
  XOR U17686 ( .A(b[19]), .B(a[114]), .Z(n17500) );
  NANDN U17687 ( .A(n18758), .B(n17500), .Z(n17369) );
  NAND U17688 ( .A(n17370), .B(n17369), .Z(n17513) );
  XOR U17689 ( .A(n17514), .B(n17513), .Z(n17516) );
  XNOR U17690 ( .A(n17515), .B(n17516), .Z(n17456) );
  XNOR U17691 ( .A(n17457), .B(n17456), .Z(n17458) );
  NANDN U17692 ( .A(n17372), .B(n17371), .Z(n17376) );
  OR U17693 ( .A(n17374), .B(n17373), .Z(n17375) );
  NAND U17694 ( .A(n17376), .B(n17375), .Z(n17459) );
  XNOR U17695 ( .A(n17458), .B(n17459), .Z(n17468) );
  NANDN U17696 ( .A(n19237), .B(n17377), .Z(n17379) );
  XOR U17697 ( .A(b[27]), .B(a[106]), .Z(n17510) );
  NANDN U17698 ( .A(n19277), .B(n17510), .Z(n17378) );
  AND U17699 ( .A(n17379), .B(n17378), .Z(n17488) );
  NANDN U17700 ( .A(n17613), .B(n17380), .Z(n17382) );
  XOR U17701 ( .A(a[124]), .B(b[9]), .Z(n17507) );
  NANDN U17702 ( .A(n17739), .B(n17507), .Z(n17381) );
  AND U17703 ( .A(n17382), .B(n17381), .Z(n17487) );
  NANDN U17704 ( .A(n18853), .B(n17383), .Z(n17385) );
  XOR U17705 ( .A(b[21]), .B(a[112]), .Z(n17526) );
  NANDN U17706 ( .A(n18926), .B(n17526), .Z(n17384) );
  NAND U17707 ( .A(n17385), .B(n17384), .Z(n17486) );
  XOR U17708 ( .A(n17487), .B(n17486), .Z(n17489) );
  XOR U17709 ( .A(n17488), .B(n17489), .Z(n17451) );
  NANDN U17710 ( .A(n19425), .B(n17386), .Z(n17388) );
  XOR U17711 ( .A(b[31]), .B(a[102]), .Z(n17497) );
  NANDN U17712 ( .A(n19426), .B(n17497), .Z(n17387) );
  AND U17713 ( .A(n17388), .B(n17387), .Z(n17494) );
  NAND U17714 ( .A(b[31]), .B(a[100]), .Z(n17503) );
  ANDN U17715 ( .B(n17390), .A(n17389), .Z(n17393) );
  NAND U17716 ( .A(b[5]), .B(n17391), .Z(n17392) );
  NANDN U17717 ( .A(n17393), .B(n17392), .Z(n17492) );
  XOR U17718 ( .A(n17503), .B(n17492), .Z(n17493) );
  XOR U17719 ( .A(n17494), .B(n17493), .Z(n17450) );
  XNOR U17720 ( .A(n17451), .B(n17450), .Z(n17452) );
  NANDN U17721 ( .A(n17395), .B(n17394), .Z(n17399) );
  NANDN U17722 ( .A(n17397), .B(n17396), .Z(n17398) );
  NAND U17723 ( .A(n17399), .B(n17398), .Z(n17453) );
  XOR U17724 ( .A(n17452), .B(n17453), .Z(n17469) );
  XNOR U17725 ( .A(n17468), .B(n17469), .Z(n17470) );
  XNOR U17726 ( .A(n17471), .B(n17470), .Z(n17438) );
  XNOR U17727 ( .A(n17439), .B(n17438), .Z(n17440) );
  XNOR U17728 ( .A(n17441), .B(n17440), .Z(n17552) );
  NANDN U17729 ( .A(n17401), .B(n17400), .Z(n17405) );
  OR U17730 ( .A(n17403), .B(n17402), .Z(n17404) );
  AND U17731 ( .A(n17405), .B(n17404), .Z(n17551) );
  NANDN U17732 ( .A(n17407), .B(n17406), .Z(n17411) );
  OR U17733 ( .A(n17409), .B(n17408), .Z(n17410) );
  AND U17734 ( .A(n17411), .B(n17410), .Z(n17464) );
  NANDN U17735 ( .A(n17413), .B(n17412), .Z(n17417) );
  OR U17736 ( .A(n17415), .B(n17414), .Z(n17416) );
  AND U17737 ( .A(n17417), .B(n17416), .Z(n17463) );
  NANDN U17738 ( .A(n17419), .B(n17418), .Z(n17423) );
  NANDN U17739 ( .A(n17421), .B(n17420), .Z(n17422) );
  AND U17740 ( .A(n17423), .B(n17422), .Z(n17462) );
  XOR U17741 ( .A(n17463), .B(n17462), .Z(n17465) );
  XNOR U17742 ( .A(n17464), .B(n17465), .Z(n17550) );
  XOR U17743 ( .A(n17551), .B(n17550), .Z(n17553) );
  XOR U17744 ( .A(n17552), .B(n17553), .Z(n17433) );
  XOR U17745 ( .A(n17432), .B(n17433), .Z(n17435) );
  XNOR U17746 ( .A(n17434), .B(n17435), .Z(n17426) );
  XOR U17747 ( .A(n17427), .B(n17426), .Z(n17429) );
  XNOR U17748 ( .A(n17428), .B(n17429), .Z(n17424) );
  XOR U17749 ( .A(n17425), .B(n17424), .Z(c[228]) );
  AND U17750 ( .A(n17425), .B(n17424), .Z(n17557) );
  NANDN U17751 ( .A(n17427), .B(n17426), .Z(n17431) );
  OR U17752 ( .A(n17429), .B(n17428), .Z(n17430) );
  AND U17753 ( .A(n17431), .B(n17430), .Z(n17560) );
  NANDN U17754 ( .A(n17433), .B(n17432), .Z(n17437) );
  NANDN U17755 ( .A(n17435), .B(n17434), .Z(n17436) );
  AND U17756 ( .A(n17437), .B(n17436), .Z(n17559) );
  NANDN U17757 ( .A(n17439), .B(n17438), .Z(n17443) );
  NANDN U17758 ( .A(n17441), .B(n17440), .Z(n17442) );
  AND U17759 ( .A(n17443), .B(n17442), .Z(n17566) );
  NANDN U17760 ( .A(n17445), .B(n17444), .Z(n17449) );
  NAND U17761 ( .A(n17447), .B(n17446), .Z(n17448) );
  AND U17762 ( .A(n17449), .B(n17448), .Z(n17573) );
  NANDN U17763 ( .A(n17451), .B(n17450), .Z(n17455) );
  NANDN U17764 ( .A(n17453), .B(n17452), .Z(n17454) );
  AND U17765 ( .A(n17455), .B(n17454), .Z(n17571) );
  NANDN U17766 ( .A(n17457), .B(n17456), .Z(n17461) );
  NANDN U17767 ( .A(n17459), .B(n17458), .Z(n17460) );
  NAND U17768 ( .A(n17461), .B(n17460), .Z(n17570) );
  XNOR U17769 ( .A(n17571), .B(n17570), .Z(n17572) );
  XOR U17770 ( .A(n17573), .B(n17572), .Z(n17565) );
  NANDN U17771 ( .A(n17463), .B(n17462), .Z(n17467) );
  OR U17772 ( .A(n17465), .B(n17464), .Z(n17466) );
  NAND U17773 ( .A(n17467), .B(n17466), .Z(n17564) );
  XOR U17774 ( .A(n17565), .B(n17564), .Z(n17567) );
  XNOR U17775 ( .A(n17566), .B(n17567), .Z(n17684) );
  NANDN U17776 ( .A(n17469), .B(n17468), .Z(n17473) );
  NANDN U17777 ( .A(n17471), .B(n17470), .Z(n17472) );
  AND U17778 ( .A(n17473), .B(n17472), .Z(n17680) );
  NAND U17779 ( .A(n17475), .B(n17474), .Z(n17479) );
  NAND U17780 ( .A(n17477), .B(n17476), .Z(n17478) );
  AND U17781 ( .A(n17479), .B(n17478), .Z(n17679) );
  NANDN U17782 ( .A(n17481), .B(n17480), .Z(n17485) );
  NANDN U17783 ( .A(n17483), .B(n17482), .Z(n17484) );
  AND U17784 ( .A(n17485), .B(n17484), .Z(n17640) );
  NANDN U17785 ( .A(n17487), .B(n17486), .Z(n17491) );
  OR U17786 ( .A(n17489), .B(n17488), .Z(n17490) );
  NAND U17787 ( .A(n17491), .B(n17490), .Z(n17639) );
  XNOR U17788 ( .A(n17640), .B(n17639), .Z(n17642) );
  IV U17789 ( .A(n17503), .Z(n17660) );
  NANDN U17790 ( .A(n17660), .B(n17492), .Z(n17496) );
  NANDN U17791 ( .A(n17494), .B(n17493), .Z(n17495) );
  AND U17792 ( .A(n17496), .B(n17495), .Z(n17591) );
  NANDN U17793 ( .A(n19425), .B(n17497), .Z(n17499) );
  XOR U17794 ( .A(b[31]), .B(a[103]), .Z(n17619) );
  NANDN U17795 ( .A(n19426), .B(n17619), .Z(n17498) );
  AND U17796 ( .A(n17499), .B(n17498), .Z(n17628) );
  NANDN U17797 ( .A(n18673), .B(n17500), .Z(n17502) );
  XOR U17798 ( .A(b[19]), .B(a[115]), .Z(n17597) );
  NANDN U17799 ( .A(n18758), .B(n17597), .Z(n17501) );
  NAND U17800 ( .A(n17502), .B(n17501), .Z(n17627) );
  XNOR U17801 ( .A(n17628), .B(n17627), .Z(n17629) );
  AND U17802 ( .A(b[31]), .B(a[101]), .Z(n17657) );
  XOR U17803 ( .A(n17658), .B(n17657), .Z(n17659) );
  XOR U17804 ( .A(n17503), .B(n17659), .Z(n17630) );
  XOR U17805 ( .A(n17629), .B(n17630), .Z(n17588) );
  NANDN U17806 ( .A(n19005), .B(n17504), .Z(n17506) );
  XOR U17807 ( .A(b[23]), .B(a[111]), .Z(n17594) );
  NANDN U17808 ( .A(n19055), .B(n17594), .Z(n17505) );
  AND U17809 ( .A(n17506), .B(n17505), .Z(n17654) );
  NANDN U17810 ( .A(n17613), .B(n17507), .Z(n17509) );
  XOR U17811 ( .A(a[125]), .B(b[9]), .Z(n17612) );
  NANDN U17812 ( .A(n17739), .B(n17612), .Z(n17508) );
  AND U17813 ( .A(n17509), .B(n17508), .Z(n17652) );
  NANDN U17814 ( .A(n19237), .B(n17510), .Z(n17512) );
  XOR U17815 ( .A(b[27]), .B(a[107]), .Z(n17600) );
  NANDN U17816 ( .A(n19277), .B(n17600), .Z(n17511) );
  NAND U17817 ( .A(n17512), .B(n17511), .Z(n17651) );
  XNOR U17818 ( .A(n17652), .B(n17651), .Z(n17653) );
  XOR U17819 ( .A(n17654), .B(n17653), .Z(n17589) );
  XNOR U17820 ( .A(n17588), .B(n17589), .Z(n17590) );
  XNOR U17821 ( .A(n17591), .B(n17590), .Z(n17641) );
  XOR U17822 ( .A(n17642), .B(n17641), .Z(n17578) );
  NANDN U17823 ( .A(n17514), .B(n17513), .Z(n17518) );
  OR U17824 ( .A(n17516), .B(n17515), .Z(n17517) );
  AND U17825 ( .A(n17518), .B(n17517), .Z(n17583) );
  NANDN U17826 ( .A(n19394), .B(n17519), .Z(n17521) );
  XOR U17827 ( .A(b[29]), .B(a[105]), .Z(n17603) );
  NANDN U17828 ( .A(n19395), .B(n17603), .Z(n17520) );
  AND U17829 ( .A(n17521), .B(n17520), .Z(n17675) );
  XNOR U17830 ( .A(a[127]), .B(b[7]), .Z(n17622) );
  OR U17831 ( .A(n17622), .B(n17522), .Z(n17525) );
  NAND U17832 ( .A(n17623), .B(n17523), .Z(n17524) );
  AND U17833 ( .A(n17525), .B(n17524), .Z(n17673) );
  NANDN U17834 ( .A(n18853), .B(n17526), .Z(n17528) );
  XOR U17835 ( .A(b[21]), .B(a[113]), .Z(n17616) );
  NANDN U17836 ( .A(n18926), .B(n17616), .Z(n17527) );
  NAND U17837 ( .A(n17528), .B(n17527), .Z(n17672) );
  XNOR U17838 ( .A(n17673), .B(n17672), .Z(n17674) );
  XNOR U17839 ( .A(n17675), .B(n17674), .Z(n17582) );
  XNOR U17840 ( .A(n17583), .B(n17582), .Z(n17585) );
  NANDN U17841 ( .A(n18487), .B(n17529), .Z(n17531) );
  XOR U17842 ( .A(a[119]), .B(b[15]), .Z(n17663) );
  NANDN U17843 ( .A(n18311), .B(n17663), .Z(n17530) );
  AND U17844 ( .A(n17531), .B(n17530), .Z(n17648) );
  NANDN U17845 ( .A(n18113), .B(n17532), .Z(n17534) );
  XOR U17846 ( .A(a[121]), .B(b[13]), .Z(n17666) );
  NANDN U17847 ( .A(n18229), .B(n17666), .Z(n17533) );
  AND U17848 ( .A(n17534), .B(n17533), .Z(n17646) );
  NANDN U17849 ( .A(n18514), .B(n17535), .Z(n17537) );
  XOR U17850 ( .A(a[117]), .B(b[17]), .Z(n17606) );
  NANDN U17851 ( .A(n18585), .B(n17606), .Z(n17536) );
  AND U17852 ( .A(n17537), .B(n17536), .Z(n17636) );
  NANDN U17853 ( .A(n19116), .B(n17538), .Z(n17540) );
  XOR U17854 ( .A(b[25]), .B(a[109]), .Z(n17669) );
  NANDN U17855 ( .A(n19179), .B(n17669), .Z(n17539) );
  AND U17856 ( .A(n17540), .B(n17539), .Z(n17634) );
  NANDN U17857 ( .A(n17888), .B(n17541), .Z(n17543) );
  XOR U17858 ( .A(a[123]), .B(b[11]), .Z(n17609) );
  NANDN U17859 ( .A(n18025), .B(n17609), .Z(n17542) );
  NAND U17860 ( .A(n17543), .B(n17542), .Z(n17633) );
  XNOR U17861 ( .A(n17634), .B(n17633), .Z(n17635) );
  XNOR U17862 ( .A(n17636), .B(n17635), .Z(n17645) );
  XNOR U17863 ( .A(n17646), .B(n17645), .Z(n17647) );
  XNOR U17864 ( .A(n17648), .B(n17647), .Z(n17584) );
  XOR U17865 ( .A(n17585), .B(n17584), .Z(n17577) );
  NANDN U17866 ( .A(n17545), .B(n17544), .Z(n17549) );
  OR U17867 ( .A(n17547), .B(n17546), .Z(n17548) );
  AND U17868 ( .A(n17549), .B(n17548), .Z(n17576) );
  XOR U17869 ( .A(n17577), .B(n17576), .Z(n17579) );
  XNOR U17870 ( .A(n17578), .B(n17579), .Z(n17678) );
  XOR U17871 ( .A(n17679), .B(n17678), .Z(n17681) );
  XOR U17872 ( .A(n17680), .B(n17681), .Z(n17685) );
  XNOR U17873 ( .A(n17684), .B(n17685), .Z(n17687) );
  NANDN U17874 ( .A(n17551), .B(n17550), .Z(n17555) );
  NANDN U17875 ( .A(n17553), .B(n17552), .Z(n17554) );
  AND U17876 ( .A(n17555), .B(n17554), .Z(n17686) );
  XNOR U17877 ( .A(n17687), .B(n17686), .Z(n17558) );
  XOR U17878 ( .A(n17559), .B(n17558), .Z(n17561) );
  XNOR U17879 ( .A(n17560), .B(n17561), .Z(n17556) );
  XOR U17880 ( .A(n17557), .B(n17556), .Z(c[229]) );
  AND U17881 ( .A(n17557), .B(n17556), .Z(n17691) );
  NANDN U17882 ( .A(n17559), .B(n17558), .Z(n17563) );
  OR U17883 ( .A(n17561), .B(n17560), .Z(n17562) );
  AND U17884 ( .A(n17563), .B(n17562), .Z(n17694) );
  NANDN U17885 ( .A(n17565), .B(n17564), .Z(n17569) );
  NANDN U17886 ( .A(n17567), .B(n17566), .Z(n17568) );
  AND U17887 ( .A(n17569), .B(n17568), .Z(n17700) );
  NANDN U17888 ( .A(n17571), .B(n17570), .Z(n17575) );
  NAND U17889 ( .A(n17573), .B(n17572), .Z(n17574) );
  AND U17890 ( .A(n17575), .B(n17574), .Z(n17706) );
  NANDN U17891 ( .A(n17577), .B(n17576), .Z(n17581) );
  OR U17892 ( .A(n17579), .B(n17578), .Z(n17580) );
  AND U17893 ( .A(n17581), .B(n17580), .Z(n17705) );
  NANDN U17894 ( .A(n17583), .B(n17582), .Z(n17587) );
  NAND U17895 ( .A(n17585), .B(n17584), .Z(n17586) );
  AND U17896 ( .A(n17587), .B(n17586), .Z(n17810) );
  NANDN U17897 ( .A(n17589), .B(n17588), .Z(n17593) );
  NANDN U17898 ( .A(n17591), .B(n17590), .Z(n17592) );
  AND U17899 ( .A(n17593), .B(n17592), .Z(n17809) );
  NANDN U17900 ( .A(n19005), .B(n17594), .Z(n17596) );
  XOR U17901 ( .A(b[23]), .B(a[112]), .Z(n17754) );
  NANDN U17902 ( .A(n19055), .B(n17754), .Z(n17595) );
  AND U17903 ( .A(n17596), .B(n17595), .Z(n17786) );
  NANDN U17904 ( .A(n18673), .B(n17597), .Z(n17599) );
  XOR U17905 ( .A(b[19]), .B(a[116]), .Z(n17775) );
  NANDN U17906 ( .A(n18758), .B(n17775), .Z(n17598) );
  AND U17907 ( .A(n17599), .B(n17598), .Z(n17785) );
  NANDN U17908 ( .A(n19237), .B(n17600), .Z(n17602) );
  XOR U17909 ( .A(b[27]), .B(a[108]), .Z(n17763) );
  NANDN U17910 ( .A(n19277), .B(n17763), .Z(n17601) );
  AND U17911 ( .A(n17602), .B(n17601), .Z(n17731) );
  NANDN U17912 ( .A(n19394), .B(n17603), .Z(n17605) );
  XOR U17913 ( .A(b[29]), .B(a[106]), .Z(n17748) );
  NANDN U17914 ( .A(n19395), .B(n17748), .Z(n17604) );
  AND U17915 ( .A(n17605), .B(n17604), .Z(n17729) );
  NANDN U17916 ( .A(n18514), .B(n17606), .Z(n17608) );
  XOR U17917 ( .A(a[118]), .B(b[17]), .Z(n17772) );
  NANDN U17918 ( .A(n18585), .B(n17772), .Z(n17607) );
  NAND U17919 ( .A(n17608), .B(n17607), .Z(n17728) );
  XNOR U17920 ( .A(n17729), .B(n17728), .Z(n17730) );
  XNOR U17921 ( .A(n17731), .B(n17730), .Z(n17784) );
  XOR U17922 ( .A(n17785), .B(n17784), .Z(n17787) );
  XOR U17923 ( .A(n17786), .B(n17787), .Z(n17804) );
  NANDN U17924 ( .A(n17888), .B(n17609), .Z(n17611) );
  XOR U17925 ( .A(a[124]), .B(b[11]), .Z(n17766) );
  NANDN U17926 ( .A(n18025), .B(n17766), .Z(n17610) );
  AND U17927 ( .A(n17611), .B(n17610), .Z(n17724) );
  NANDN U17928 ( .A(n17613), .B(n17612), .Z(n17615) );
  XOR U17929 ( .A(a[126]), .B(b[9]), .Z(n17740) );
  NANDN U17930 ( .A(n17739), .B(n17740), .Z(n17614) );
  AND U17931 ( .A(n17615), .B(n17614), .Z(n17723) );
  NANDN U17932 ( .A(n18853), .B(n17616), .Z(n17618) );
  XOR U17933 ( .A(b[21]), .B(a[114]), .Z(n17743) );
  NANDN U17934 ( .A(n18926), .B(n17743), .Z(n17617) );
  NAND U17935 ( .A(n17618), .B(n17617), .Z(n17722) );
  XOR U17936 ( .A(n17723), .B(n17722), .Z(n17725) );
  XOR U17937 ( .A(n17724), .B(n17725), .Z(n17803) );
  NANDN U17938 ( .A(n19425), .B(n17619), .Z(n17621) );
  XOR U17939 ( .A(b[31]), .B(a[104]), .Z(n17751) );
  NANDN U17940 ( .A(n19426), .B(n17751), .Z(n17620) );
  AND U17941 ( .A(n17621), .B(n17620), .Z(n17736) );
  NAND U17942 ( .A(b[31]), .B(a[102]), .Z(n17747) );
  ANDN U17943 ( .B(n17623), .A(n17622), .Z(n17626) );
  NAND U17944 ( .A(b[7]), .B(n17624), .Z(n17625) );
  NANDN U17945 ( .A(n17626), .B(n17625), .Z(n17734) );
  XOR U17946 ( .A(n17747), .B(n17734), .Z(n17735) );
  XOR U17947 ( .A(n17736), .B(n17735), .Z(n17802) );
  XOR U17948 ( .A(n17803), .B(n17802), .Z(n17805) );
  XOR U17949 ( .A(n17804), .B(n17805), .Z(n17793) );
  NANDN U17950 ( .A(n17628), .B(n17627), .Z(n17632) );
  NAND U17951 ( .A(n17630), .B(n17629), .Z(n17631) );
  AND U17952 ( .A(n17632), .B(n17631), .Z(n17791) );
  NANDN U17953 ( .A(n17634), .B(n17633), .Z(n17638) );
  NANDN U17954 ( .A(n17636), .B(n17635), .Z(n17637) );
  NAND U17955 ( .A(n17638), .B(n17637), .Z(n17790) );
  XNOR U17956 ( .A(n17791), .B(n17790), .Z(n17792) );
  XNOR U17957 ( .A(n17793), .B(n17792), .Z(n17808) );
  XOR U17958 ( .A(n17809), .B(n17808), .Z(n17811) );
  XOR U17959 ( .A(n17810), .B(n17811), .Z(n17713) );
  NANDN U17960 ( .A(n17640), .B(n17639), .Z(n17644) );
  NAND U17961 ( .A(n17642), .B(n17641), .Z(n17643) );
  AND U17962 ( .A(n17644), .B(n17643), .Z(n17710) );
  NANDN U17963 ( .A(n17646), .B(n17645), .Z(n17650) );
  NANDN U17964 ( .A(n17648), .B(n17647), .Z(n17649) );
  AND U17965 ( .A(n17650), .B(n17649), .Z(n17718) );
  NANDN U17966 ( .A(n17652), .B(n17651), .Z(n17656) );
  NANDN U17967 ( .A(n17654), .B(n17653), .Z(n17655) );
  AND U17968 ( .A(n17656), .B(n17655), .Z(n17798) );
  NANDN U17969 ( .A(n17658), .B(n17657), .Z(n17662) );
  ANDN U17970 ( .B(n17660), .A(n17659), .Z(n17661) );
  ANDN U17971 ( .B(n17662), .A(n17661), .Z(n17797) );
  NANDN U17972 ( .A(n18487), .B(n17663), .Z(n17665) );
  XOR U17973 ( .A(a[120]), .B(b[15]), .Z(n17781) );
  NANDN U17974 ( .A(n18311), .B(n17781), .Z(n17664) );
  AND U17975 ( .A(n17665), .B(n17664), .Z(n17760) );
  NANDN U17976 ( .A(n18113), .B(n17666), .Z(n17668) );
  XOR U17977 ( .A(a[122]), .B(b[13]), .Z(n17778) );
  NANDN U17978 ( .A(n18229), .B(n17778), .Z(n17667) );
  AND U17979 ( .A(n17668), .B(n17667), .Z(n17758) );
  NANDN U17980 ( .A(n19116), .B(n17669), .Z(n17671) );
  XOR U17981 ( .A(b[25]), .B(a[110]), .Z(n17769) );
  NANDN U17982 ( .A(n19179), .B(n17769), .Z(n17670) );
  NAND U17983 ( .A(n17671), .B(n17670), .Z(n17757) );
  XNOR U17984 ( .A(n17758), .B(n17757), .Z(n17759) );
  XNOR U17985 ( .A(n17760), .B(n17759), .Z(n17796) );
  XOR U17986 ( .A(n17797), .B(n17796), .Z(n17799) );
  XOR U17987 ( .A(n17798), .B(n17799), .Z(n17717) );
  NANDN U17988 ( .A(n17673), .B(n17672), .Z(n17677) );
  NANDN U17989 ( .A(n17675), .B(n17674), .Z(n17676) );
  AND U17990 ( .A(n17677), .B(n17676), .Z(n17716) );
  XOR U17991 ( .A(n17717), .B(n17716), .Z(n17719) );
  XOR U17992 ( .A(n17718), .B(n17719), .Z(n17711) );
  XNOR U17993 ( .A(n17710), .B(n17711), .Z(n17712) );
  XNOR U17994 ( .A(n17713), .B(n17712), .Z(n17704) );
  XOR U17995 ( .A(n17705), .B(n17704), .Z(n17707) );
  XOR U17996 ( .A(n17706), .B(n17707), .Z(n17699) );
  NANDN U17997 ( .A(n17679), .B(n17678), .Z(n17683) );
  NANDN U17998 ( .A(n17681), .B(n17680), .Z(n17682) );
  NAND U17999 ( .A(n17683), .B(n17682), .Z(n17698) );
  XOR U18000 ( .A(n17699), .B(n17698), .Z(n17701) );
  XOR U18001 ( .A(n17700), .B(n17701), .Z(n17693) );
  NANDN U18002 ( .A(n17685), .B(n17684), .Z(n17689) );
  NAND U18003 ( .A(n17687), .B(n17686), .Z(n17688) );
  AND U18004 ( .A(n17689), .B(n17688), .Z(n17692) );
  XOR U18005 ( .A(n17693), .B(n17692), .Z(n17695) );
  XNOR U18006 ( .A(n17694), .B(n17695), .Z(n17690) );
  XOR U18007 ( .A(n17691), .B(n17690), .Z(c[230]) );
  AND U18008 ( .A(n17691), .B(n17690), .Z(n17815) );
  NANDN U18009 ( .A(n17693), .B(n17692), .Z(n17697) );
  OR U18010 ( .A(n17695), .B(n17694), .Z(n17696) );
  AND U18011 ( .A(n17697), .B(n17696), .Z(n17818) );
  NANDN U18012 ( .A(n17699), .B(n17698), .Z(n17703) );
  OR U18013 ( .A(n17701), .B(n17700), .Z(n17702) );
  AND U18014 ( .A(n17703), .B(n17702), .Z(n17816) );
  NANDN U18015 ( .A(n17705), .B(n17704), .Z(n17709) );
  OR U18016 ( .A(n17707), .B(n17706), .Z(n17708) );
  AND U18017 ( .A(n17709), .B(n17708), .Z(n17825) );
  NANDN U18018 ( .A(n17711), .B(n17710), .Z(n17715) );
  NANDN U18019 ( .A(n17713), .B(n17712), .Z(n17714) );
  AND U18020 ( .A(n17715), .B(n17714), .Z(n17823) );
  NANDN U18021 ( .A(n17717), .B(n17716), .Z(n17721) );
  NANDN U18022 ( .A(n17719), .B(n17718), .Z(n17720) );
  AND U18023 ( .A(n17721), .B(n17720), .Z(n17936) );
  NANDN U18024 ( .A(n17723), .B(n17722), .Z(n17727) );
  OR U18025 ( .A(n17725), .B(n17724), .Z(n17726) );
  AND U18026 ( .A(n17727), .B(n17726), .Z(n17910) );
  NANDN U18027 ( .A(n17729), .B(n17728), .Z(n17733) );
  NANDN U18028 ( .A(n17731), .B(n17730), .Z(n17732) );
  NAND U18029 ( .A(n17733), .B(n17732), .Z(n17909) );
  XNOR U18030 ( .A(n17910), .B(n17909), .Z(n17912) );
  IV U18031 ( .A(n17747), .Z(n17876) );
  NANDN U18032 ( .A(n17876), .B(n17734), .Z(n17738) );
  NANDN U18033 ( .A(n17736), .B(n17735), .Z(n17737) );
  AND U18034 ( .A(n17738), .B(n17737), .Z(n17924) );
  XNOR U18035 ( .A(a[127]), .B(b[9]), .Z(n17880) );
  OR U18036 ( .A(n17880), .B(n17739), .Z(n17742) );
  NAND U18037 ( .A(n17881), .B(n17740), .Z(n17741) );
  AND U18038 ( .A(n17742), .B(n17741), .Z(n17898) );
  NANDN U18039 ( .A(n18853), .B(n17743), .Z(n17745) );
  XOR U18040 ( .A(b[21]), .B(a[115]), .Z(n17894) );
  NANDN U18041 ( .A(n18926), .B(n17894), .Z(n17744) );
  NAND U18042 ( .A(n17745), .B(n17744), .Z(n17897) );
  XNOR U18043 ( .A(n17898), .B(n17897), .Z(n17899) );
  IV U18044 ( .A(n17746), .Z(n17874) );
  AND U18045 ( .A(b[31]), .B(a[103]), .Z(n17873) );
  XOR U18046 ( .A(n17874), .B(n17873), .Z(n17875) );
  XOR U18047 ( .A(n17747), .B(n17875), .Z(n17900) );
  XOR U18048 ( .A(n17899), .B(n17900), .Z(n17921) );
  NANDN U18049 ( .A(n19394), .B(n17748), .Z(n17750) );
  XOR U18050 ( .A(b[29]), .B(a[107]), .Z(n17891) );
  NANDN U18051 ( .A(n19395), .B(n17891), .Z(n17749) );
  AND U18052 ( .A(n17750), .B(n17749), .Z(n17864) );
  NANDN U18053 ( .A(n19425), .B(n17751), .Z(n17753) );
  XOR U18054 ( .A(b[31]), .B(a[105]), .Z(n17884) );
  NANDN U18055 ( .A(n19426), .B(n17884), .Z(n17752) );
  AND U18056 ( .A(n17753), .B(n17752), .Z(n17862) );
  NANDN U18057 ( .A(n19005), .B(n17754), .Z(n17756) );
  XOR U18058 ( .A(b[23]), .B(a[113]), .Z(n17846) );
  NANDN U18059 ( .A(n19055), .B(n17846), .Z(n17755) );
  NAND U18060 ( .A(n17756), .B(n17755), .Z(n17861) );
  XNOR U18061 ( .A(n17862), .B(n17861), .Z(n17863) );
  XOR U18062 ( .A(n17864), .B(n17863), .Z(n17922) );
  XNOR U18063 ( .A(n17921), .B(n17922), .Z(n17923) );
  XNOR U18064 ( .A(n17924), .B(n17923), .Z(n17911) );
  XOR U18065 ( .A(n17912), .B(n17911), .Z(n17934) );
  NANDN U18066 ( .A(n17758), .B(n17757), .Z(n17762) );
  NANDN U18067 ( .A(n17760), .B(n17759), .Z(n17761) );
  AND U18068 ( .A(n17762), .B(n17761), .Z(n17834) );
  NANDN U18069 ( .A(n19237), .B(n17763), .Z(n17765) );
  XOR U18070 ( .A(b[27]), .B(a[109]), .Z(n17843) );
  NANDN U18071 ( .A(n19277), .B(n17843), .Z(n17764) );
  AND U18072 ( .A(n17765), .B(n17764), .Z(n17869) );
  NANDN U18073 ( .A(n17888), .B(n17766), .Z(n17768) );
  XOR U18074 ( .A(a[125]), .B(b[11]), .Z(n17887) );
  NANDN U18075 ( .A(n18025), .B(n17887), .Z(n17767) );
  AND U18076 ( .A(n17768), .B(n17767), .Z(n17868) );
  NANDN U18077 ( .A(n19116), .B(n17769), .Z(n17771) );
  XOR U18078 ( .A(b[25]), .B(a[111]), .Z(n17840) );
  NANDN U18079 ( .A(n19179), .B(n17840), .Z(n17770) );
  NAND U18080 ( .A(n17771), .B(n17770), .Z(n17867) );
  XOR U18081 ( .A(n17868), .B(n17867), .Z(n17870) );
  XOR U18082 ( .A(n17869), .B(n17870), .Z(n17918) );
  NANDN U18083 ( .A(n18514), .B(n17772), .Z(n17774) );
  XNOR U18084 ( .A(a[119]), .B(b[17]), .Z(n17858) );
  NANDN U18085 ( .A(n17858), .B(n18684), .Z(n17773) );
  AND U18086 ( .A(n17774), .B(n17773), .Z(n17905) );
  NANDN U18087 ( .A(n18673), .B(n17775), .Z(n17777) );
  XOR U18088 ( .A(b[19]), .B(a[117]), .Z(n17852) );
  NANDN U18089 ( .A(n18758), .B(n17852), .Z(n17776) );
  AND U18090 ( .A(n17777), .B(n17776), .Z(n17904) );
  NANDN U18091 ( .A(n18113), .B(n17778), .Z(n17780) );
  XOR U18092 ( .A(a[123]), .B(b[13]), .Z(n17855) );
  NANDN U18093 ( .A(n18229), .B(n17855), .Z(n17779) );
  NAND U18094 ( .A(n17780), .B(n17779), .Z(n17903) );
  XOR U18095 ( .A(n17904), .B(n17903), .Z(n17906) );
  XOR U18096 ( .A(n17905), .B(n17906), .Z(n17916) );
  NAND U18097 ( .A(n18439), .B(n17781), .Z(n17783) );
  XNOR U18098 ( .A(a[121]), .B(b[15]), .Z(n17849) );
  NANDN U18099 ( .A(n17849), .B(n18486), .Z(n17782) );
  AND U18100 ( .A(n17783), .B(n17782), .Z(n17915) );
  XNOR U18101 ( .A(n17916), .B(n17915), .Z(n17917) );
  XOR U18102 ( .A(n17918), .B(n17917), .Z(n17835) );
  XNOR U18103 ( .A(n17834), .B(n17835), .Z(n17836) );
  NANDN U18104 ( .A(n17785), .B(n17784), .Z(n17789) );
  OR U18105 ( .A(n17787), .B(n17786), .Z(n17788) );
  NAND U18106 ( .A(n17789), .B(n17788), .Z(n17837) );
  XNOR U18107 ( .A(n17836), .B(n17837), .Z(n17933) );
  XNOR U18108 ( .A(n17934), .B(n17933), .Z(n17935) );
  XNOR U18109 ( .A(n17936), .B(n17935), .Z(n17830) );
  NANDN U18110 ( .A(n17791), .B(n17790), .Z(n17795) );
  NANDN U18111 ( .A(n17793), .B(n17792), .Z(n17794) );
  AND U18112 ( .A(n17795), .B(n17794), .Z(n17929) );
  NANDN U18113 ( .A(n17797), .B(n17796), .Z(n17801) );
  OR U18114 ( .A(n17799), .B(n17798), .Z(n17800) );
  AND U18115 ( .A(n17801), .B(n17800), .Z(n17928) );
  NANDN U18116 ( .A(n17803), .B(n17802), .Z(n17807) );
  OR U18117 ( .A(n17805), .B(n17804), .Z(n17806) );
  AND U18118 ( .A(n17807), .B(n17806), .Z(n17927) );
  XOR U18119 ( .A(n17928), .B(n17927), .Z(n17930) );
  XOR U18120 ( .A(n17929), .B(n17930), .Z(n17829) );
  NANDN U18121 ( .A(n17809), .B(n17808), .Z(n17813) );
  OR U18122 ( .A(n17811), .B(n17810), .Z(n17812) );
  AND U18123 ( .A(n17813), .B(n17812), .Z(n17828) );
  XOR U18124 ( .A(n17829), .B(n17828), .Z(n17831) );
  XNOR U18125 ( .A(n17830), .B(n17831), .Z(n17822) );
  XNOR U18126 ( .A(n17823), .B(n17822), .Z(n17824) );
  XOR U18127 ( .A(n17825), .B(n17824), .Z(n17817) );
  XOR U18128 ( .A(n17816), .B(n17817), .Z(n17819) );
  XNOR U18129 ( .A(n17818), .B(n17819), .Z(n17814) );
  XOR U18130 ( .A(n17815), .B(n17814), .Z(c[231]) );
  AND U18131 ( .A(n17815), .B(n17814), .Z(n17940) );
  NANDN U18132 ( .A(n17817), .B(n17816), .Z(n17821) );
  OR U18133 ( .A(n17819), .B(n17818), .Z(n17820) );
  AND U18134 ( .A(n17821), .B(n17820), .Z(n17943) );
  NANDN U18135 ( .A(n17823), .B(n17822), .Z(n17827) );
  NANDN U18136 ( .A(n17825), .B(n17824), .Z(n17826) );
  AND U18137 ( .A(n17827), .B(n17826), .Z(n17942) );
  NANDN U18138 ( .A(n17829), .B(n17828), .Z(n17833) );
  NANDN U18139 ( .A(n17831), .B(n17830), .Z(n17832) );
  AND U18140 ( .A(n17833), .B(n17832), .Z(n17950) );
  NANDN U18141 ( .A(n17835), .B(n17834), .Z(n17839) );
  NANDN U18142 ( .A(n17837), .B(n17836), .Z(n17838) );
  AND U18143 ( .A(n17839), .B(n17838), .Z(n18046) );
  NANDN U18144 ( .A(n19116), .B(n17840), .Z(n17842) );
  XOR U18145 ( .A(b[25]), .B(a[112]), .Z(n18004) );
  NANDN U18146 ( .A(n19179), .B(n18004), .Z(n17841) );
  AND U18147 ( .A(n17842), .B(n17841), .Z(n17985) );
  NANDN U18148 ( .A(n19237), .B(n17843), .Z(n17845) );
  XOR U18149 ( .A(b[27]), .B(a[110]), .Z(n18007) );
  NANDN U18150 ( .A(n19277), .B(n18007), .Z(n17844) );
  AND U18151 ( .A(n17845), .B(n17844), .Z(n17984) );
  NANDN U18152 ( .A(n19005), .B(n17846), .Z(n17848) );
  XOR U18153 ( .A(b[23]), .B(a[114]), .Z(n18029) );
  NANDN U18154 ( .A(n19055), .B(n18029), .Z(n17847) );
  NAND U18155 ( .A(n17848), .B(n17847), .Z(n17983) );
  XOR U18156 ( .A(n17984), .B(n17983), .Z(n17986) );
  XOR U18157 ( .A(n17985), .B(n17986), .Z(n17973) );
  NANDN U18158 ( .A(n17849), .B(n18439), .Z(n17851) );
  XOR U18159 ( .A(a[122]), .B(b[15]), .Z(n18019) );
  NANDN U18160 ( .A(n18311), .B(n18019), .Z(n17850) );
  AND U18161 ( .A(n17851), .B(n17850), .Z(n18034) );
  NANDN U18162 ( .A(n18673), .B(n17852), .Z(n17854) );
  XOR U18163 ( .A(a[118]), .B(b[19]), .Z(n18010) );
  NANDN U18164 ( .A(n18758), .B(n18010), .Z(n17853) );
  AND U18165 ( .A(n17854), .B(n17853), .Z(n18033) );
  NANDN U18166 ( .A(n18113), .B(n17855), .Z(n17857) );
  XOR U18167 ( .A(a[124]), .B(b[13]), .Z(n18022) );
  NANDN U18168 ( .A(n18229), .B(n18022), .Z(n17856) );
  NAND U18169 ( .A(n17857), .B(n17856), .Z(n18032) );
  XOR U18170 ( .A(n18033), .B(n18032), .Z(n18035) );
  XOR U18171 ( .A(n18034), .B(n18035), .Z(n17972) );
  NANDN U18172 ( .A(n17858), .B(n18683), .Z(n17860) );
  XNOR U18173 ( .A(a[120]), .B(b[17]), .Z(n18016) );
  NANDN U18174 ( .A(n18016), .B(n18684), .Z(n17859) );
  AND U18175 ( .A(n17860), .B(n17859), .Z(n17971) );
  XOR U18176 ( .A(n17972), .B(n17971), .Z(n17974) );
  XOR U18177 ( .A(n17973), .B(n17974), .Z(n17961) );
  NANDN U18178 ( .A(n17862), .B(n17861), .Z(n17866) );
  NANDN U18179 ( .A(n17864), .B(n17863), .Z(n17865) );
  AND U18180 ( .A(n17866), .B(n17865), .Z(n17960) );
  NANDN U18181 ( .A(n17868), .B(n17867), .Z(n17872) );
  OR U18182 ( .A(n17870), .B(n17869), .Z(n17871) );
  AND U18183 ( .A(n17872), .B(n17871), .Z(n17980) );
  NANDN U18184 ( .A(n17874), .B(n17873), .Z(n17878) );
  ANDN U18185 ( .B(n17876), .A(n17875), .Z(n17877) );
  ANDN U18186 ( .B(n17878), .A(n17877), .Z(n17978) );
  NAND U18187 ( .A(b[9]), .B(n17879), .Z(n17883) );
  ANDN U18188 ( .B(n17881), .A(n17880), .Z(n17882) );
  ANDN U18189 ( .B(n17883), .A(n17882), .Z(n17991) );
  NAND U18190 ( .A(b[31]), .B(a[104]), .Z(n18135) );
  NANDN U18191 ( .A(n19425), .B(n17884), .Z(n17886) );
  XOR U18192 ( .A(b[31]), .B(a[106]), .Z(n17998) );
  NANDN U18193 ( .A(n19426), .B(n17998), .Z(n17885) );
  NAND U18194 ( .A(n17886), .B(n17885), .Z(n17989) );
  XOR U18195 ( .A(n18135), .B(n17989), .Z(n17990) );
  XNOR U18196 ( .A(n17991), .B(n17990), .Z(n17977) );
  XNOR U18197 ( .A(n17978), .B(n17977), .Z(n17979) );
  XNOR U18198 ( .A(n17980), .B(n17979), .Z(n17959) );
  XOR U18199 ( .A(n17960), .B(n17959), .Z(n17962) );
  XOR U18200 ( .A(n17961), .B(n17962), .Z(n18045) );
  NANDN U18201 ( .A(n17888), .B(n17887), .Z(n17890) );
  XOR U18202 ( .A(a[126]), .B(b[11]), .Z(n18026) );
  NANDN U18203 ( .A(n18025), .B(n18026), .Z(n17889) );
  AND U18204 ( .A(n17890), .B(n17889), .Z(n17994) );
  NANDN U18205 ( .A(n19394), .B(n17891), .Z(n17893) );
  XOR U18206 ( .A(b[29]), .B(a[108]), .Z(n18013) );
  NANDN U18207 ( .A(n19395), .B(n18013), .Z(n17892) );
  AND U18208 ( .A(n17893), .B(n17892), .Z(n17993) );
  NANDN U18209 ( .A(n18853), .B(n17894), .Z(n17896) );
  XOR U18210 ( .A(b[21]), .B(a[116]), .Z(n18001) );
  NANDN U18211 ( .A(n18926), .B(n18001), .Z(n17895) );
  NAND U18212 ( .A(n17896), .B(n17895), .Z(n17992) );
  XOR U18213 ( .A(n17993), .B(n17992), .Z(n17995) );
  XOR U18214 ( .A(n17994), .B(n17995), .Z(n17966) );
  NANDN U18215 ( .A(n17898), .B(n17897), .Z(n17902) );
  NAND U18216 ( .A(n17900), .B(n17899), .Z(n17901) );
  AND U18217 ( .A(n17902), .B(n17901), .Z(n17965) );
  XNOR U18218 ( .A(n17966), .B(n17965), .Z(n17967) );
  NANDN U18219 ( .A(n17904), .B(n17903), .Z(n17908) );
  OR U18220 ( .A(n17906), .B(n17905), .Z(n17907) );
  NAND U18221 ( .A(n17908), .B(n17907), .Z(n17968) );
  XNOR U18222 ( .A(n17967), .B(n17968), .Z(n18044) );
  XOR U18223 ( .A(n18045), .B(n18044), .Z(n18047) );
  XOR U18224 ( .A(n18046), .B(n18047), .Z(n17955) );
  NANDN U18225 ( .A(n17910), .B(n17909), .Z(n17914) );
  NAND U18226 ( .A(n17912), .B(n17911), .Z(n17913) );
  AND U18227 ( .A(n17914), .B(n17913), .Z(n18041) );
  NANDN U18228 ( .A(n17916), .B(n17915), .Z(n17920) );
  NANDN U18229 ( .A(n17918), .B(n17917), .Z(n17919) );
  AND U18230 ( .A(n17920), .B(n17919), .Z(n18039) );
  NANDN U18231 ( .A(n17922), .B(n17921), .Z(n17926) );
  NANDN U18232 ( .A(n17924), .B(n17923), .Z(n17925) );
  AND U18233 ( .A(n17926), .B(n17925), .Z(n18038) );
  XNOR U18234 ( .A(n18039), .B(n18038), .Z(n18040) );
  XOR U18235 ( .A(n18041), .B(n18040), .Z(n17954) );
  NANDN U18236 ( .A(n17928), .B(n17927), .Z(n17932) );
  OR U18237 ( .A(n17930), .B(n17929), .Z(n17931) );
  NAND U18238 ( .A(n17932), .B(n17931), .Z(n17953) );
  XOR U18239 ( .A(n17954), .B(n17953), .Z(n17956) );
  XOR U18240 ( .A(n17955), .B(n17956), .Z(n17948) );
  NANDN U18241 ( .A(n17934), .B(n17933), .Z(n17938) );
  NANDN U18242 ( .A(n17936), .B(n17935), .Z(n17937) );
  NAND U18243 ( .A(n17938), .B(n17937), .Z(n17947) );
  XNOR U18244 ( .A(n17948), .B(n17947), .Z(n17949) );
  XNOR U18245 ( .A(n17950), .B(n17949), .Z(n17941) );
  XOR U18246 ( .A(n17942), .B(n17941), .Z(n17944) );
  XNOR U18247 ( .A(n17943), .B(n17944), .Z(n17939) );
  XOR U18248 ( .A(n17940), .B(n17939), .Z(c[232]) );
  AND U18249 ( .A(n17940), .B(n17939), .Z(n18051) );
  NANDN U18250 ( .A(n17942), .B(n17941), .Z(n17946) );
  OR U18251 ( .A(n17944), .B(n17943), .Z(n17945) );
  AND U18252 ( .A(n17946), .B(n17945), .Z(n18054) );
  NANDN U18253 ( .A(n17948), .B(n17947), .Z(n17952) );
  NANDN U18254 ( .A(n17950), .B(n17949), .Z(n17951) );
  AND U18255 ( .A(n17952), .B(n17951), .Z(n18053) );
  NANDN U18256 ( .A(n17954), .B(n17953), .Z(n17958) );
  OR U18257 ( .A(n17956), .B(n17955), .Z(n17957) );
  AND U18258 ( .A(n17958), .B(n17957), .Z(n18060) );
  NANDN U18259 ( .A(n17960), .B(n17959), .Z(n17964) );
  OR U18260 ( .A(n17962), .B(n17961), .Z(n17963) );
  AND U18261 ( .A(n17964), .B(n17963), .Z(n18067) );
  NANDN U18262 ( .A(n17966), .B(n17965), .Z(n17970) );
  NANDN U18263 ( .A(n17968), .B(n17967), .Z(n17969) );
  AND U18264 ( .A(n17970), .B(n17969), .Z(n18065) );
  NANDN U18265 ( .A(n17972), .B(n17971), .Z(n17976) );
  OR U18266 ( .A(n17974), .B(n17973), .Z(n17975) );
  NAND U18267 ( .A(n17976), .B(n17975), .Z(n18064) );
  XNOR U18268 ( .A(n18065), .B(n18064), .Z(n18066) );
  XOR U18269 ( .A(n18067), .B(n18066), .Z(n18160) );
  NANDN U18270 ( .A(n17978), .B(n17977), .Z(n17982) );
  NANDN U18271 ( .A(n17980), .B(n17979), .Z(n17981) );
  AND U18272 ( .A(n17982), .B(n17981), .Z(n18073) );
  NANDN U18273 ( .A(n17984), .B(n17983), .Z(n17988) );
  OR U18274 ( .A(n17986), .B(n17985), .Z(n17987) );
  AND U18275 ( .A(n17988), .B(n17987), .Z(n18153) );
  XNOR U18276 ( .A(n18153), .B(n18152), .Z(n18155) );
  NANDN U18277 ( .A(n17993), .B(n17992), .Z(n17997) );
  OR U18278 ( .A(n17995), .B(n17994), .Z(n17996) );
  AND U18279 ( .A(n17997), .B(n17996), .Z(n18125) );
  NANDN U18280 ( .A(n19425), .B(n17998), .Z(n18000) );
  XOR U18281 ( .A(b[31]), .B(a[107]), .Z(n18080) );
  NANDN U18282 ( .A(n19426), .B(n18080), .Z(n17999) );
  AND U18283 ( .A(n18000), .B(n17999), .Z(n18077) );
  NANDN U18284 ( .A(n18853), .B(n18001), .Z(n18003) );
  XOR U18285 ( .A(b[21]), .B(a[117]), .Z(n18091) );
  NANDN U18286 ( .A(n18926), .B(n18091), .Z(n18002) );
  NAND U18287 ( .A(n18003), .B(n18002), .Z(n18076) );
  XNOR U18288 ( .A(n18077), .B(n18076), .Z(n18079) );
  AND U18289 ( .A(b[31]), .B(a[105]), .Z(n18136) );
  XOR U18290 ( .A(n18137), .B(n18136), .Z(n18078) );
  XOR U18291 ( .A(n18079), .B(n18078), .Z(n18122) );
  NANDN U18292 ( .A(n19116), .B(n18004), .Z(n18006) );
  XOR U18293 ( .A(b[25]), .B(a[113]), .Z(n18088) );
  NANDN U18294 ( .A(n19179), .B(n18088), .Z(n18005) );
  AND U18295 ( .A(n18006), .B(n18005), .Z(n18119) );
  NANDN U18296 ( .A(n19237), .B(n18007), .Z(n18009) );
  XOR U18297 ( .A(b[27]), .B(a[111]), .Z(n18103) );
  NANDN U18298 ( .A(n19277), .B(n18103), .Z(n18008) );
  AND U18299 ( .A(n18009), .B(n18008), .Z(n18117) );
  NANDN U18300 ( .A(n18673), .B(n18010), .Z(n18012) );
  XOR U18301 ( .A(a[119]), .B(b[19]), .Z(n18094) );
  NANDN U18302 ( .A(n18758), .B(n18094), .Z(n18011) );
  NAND U18303 ( .A(n18012), .B(n18011), .Z(n18116) );
  XNOR U18304 ( .A(n18117), .B(n18116), .Z(n18118) );
  XOR U18305 ( .A(n18119), .B(n18118), .Z(n18123) );
  XNOR U18306 ( .A(n18122), .B(n18123), .Z(n18124) );
  XNOR U18307 ( .A(n18125), .B(n18124), .Z(n18154) );
  XOR U18308 ( .A(n18155), .B(n18154), .Z(n18071) );
  NANDN U18309 ( .A(n19394), .B(n18013), .Z(n18015) );
  XOR U18310 ( .A(b[29]), .B(a[109]), .Z(n18097) );
  NANDN U18311 ( .A(n19395), .B(n18097), .Z(n18014) );
  AND U18312 ( .A(n18015), .B(n18014), .Z(n18130) );
  NANDN U18313 ( .A(n18016), .B(n18683), .Z(n18018) );
  XOR U18314 ( .A(a[121]), .B(b[17]), .Z(n18100) );
  NANDN U18315 ( .A(n18585), .B(n18100), .Z(n18017) );
  AND U18316 ( .A(n18018), .B(n18017), .Z(n18129) );
  NANDN U18317 ( .A(n18487), .B(n18019), .Z(n18021) );
  XOR U18318 ( .A(a[123]), .B(b[15]), .Z(n18109) );
  NANDN U18319 ( .A(n18311), .B(n18109), .Z(n18020) );
  NAND U18320 ( .A(n18021), .B(n18020), .Z(n18128) );
  XOR U18321 ( .A(n18129), .B(n18128), .Z(n18131) );
  XOR U18322 ( .A(n18130), .B(n18131), .Z(n18147) );
  NANDN U18323 ( .A(n18113), .B(n18022), .Z(n18024) );
  XOR U18324 ( .A(a[125]), .B(b[13]), .Z(n18112) );
  NANDN U18325 ( .A(n18229), .B(n18112), .Z(n18023) );
  AND U18326 ( .A(n18024), .B(n18023), .Z(n18142) );
  XNOR U18327 ( .A(a[127]), .B(b[11]), .Z(n18083) );
  OR U18328 ( .A(n18083), .B(n18025), .Z(n18028) );
  NAND U18329 ( .A(n18084), .B(n18026), .Z(n18027) );
  AND U18330 ( .A(n18028), .B(n18027), .Z(n18141) );
  NANDN U18331 ( .A(n19005), .B(n18029), .Z(n18031) );
  XOR U18332 ( .A(b[23]), .B(a[115]), .Z(n18106) );
  NANDN U18333 ( .A(n19055), .B(n18106), .Z(n18030) );
  NAND U18334 ( .A(n18031), .B(n18030), .Z(n18140) );
  XOR U18335 ( .A(n18141), .B(n18140), .Z(n18143) );
  XNOR U18336 ( .A(n18142), .B(n18143), .Z(n18146) );
  XNOR U18337 ( .A(n18147), .B(n18146), .Z(n18148) );
  NANDN U18338 ( .A(n18033), .B(n18032), .Z(n18037) );
  OR U18339 ( .A(n18035), .B(n18034), .Z(n18036) );
  NAND U18340 ( .A(n18037), .B(n18036), .Z(n18149) );
  XNOR U18341 ( .A(n18148), .B(n18149), .Z(n18070) );
  XNOR U18342 ( .A(n18071), .B(n18070), .Z(n18072) );
  XOR U18343 ( .A(n18073), .B(n18072), .Z(n18159) );
  NANDN U18344 ( .A(n18039), .B(n18038), .Z(n18043) );
  NAND U18345 ( .A(n18041), .B(n18040), .Z(n18042) );
  AND U18346 ( .A(n18043), .B(n18042), .Z(n18158) );
  XOR U18347 ( .A(n18159), .B(n18158), .Z(n18161) );
  XOR U18348 ( .A(n18160), .B(n18161), .Z(n18059) );
  NANDN U18349 ( .A(n18045), .B(n18044), .Z(n18049) );
  OR U18350 ( .A(n18047), .B(n18046), .Z(n18048) );
  NAND U18351 ( .A(n18049), .B(n18048), .Z(n18058) );
  XOR U18352 ( .A(n18059), .B(n18058), .Z(n18061) );
  XNOR U18353 ( .A(n18060), .B(n18061), .Z(n18052) );
  XOR U18354 ( .A(n18053), .B(n18052), .Z(n18055) );
  XNOR U18355 ( .A(n18054), .B(n18055), .Z(n18050) );
  XOR U18356 ( .A(n18051), .B(n18050), .Z(c[233]) );
  AND U18357 ( .A(n18051), .B(n18050), .Z(n18165) );
  NANDN U18358 ( .A(n18053), .B(n18052), .Z(n18057) );
  OR U18359 ( .A(n18055), .B(n18054), .Z(n18056) );
  AND U18360 ( .A(n18057), .B(n18056), .Z(n18168) );
  NANDN U18361 ( .A(n18059), .B(n18058), .Z(n18063) );
  NANDN U18362 ( .A(n18061), .B(n18060), .Z(n18062) );
  AND U18363 ( .A(n18063), .B(n18062), .Z(n18167) );
  NANDN U18364 ( .A(n18065), .B(n18064), .Z(n18069) );
  NAND U18365 ( .A(n18067), .B(n18066), .Z(n18068) );
  AND U18366 ( .A(n18069), .B(n18068), .Z(n18261) );
  NANDN U18367 ( .A(n18071), .B(n18070), .Z(n18075) );
  NAND U18368 ( .A(n18073), .B(n18072), .Z(n18074) );
  AND U18369 ( .A(n18075), .B(n18074), .Z(n18257) );
  NANDN U18370 ( .A(n19425), .B(n18080), .Z(n18082) );
  XOR U18371 ( .A(b[31]), .B(a[108]), .Z(n18236) );
  NANDN U18372 ( .A(n19426), .B(n18236), .Z(n18081) );
  AND U18373 ( .A(n18082), .B(n18081), .Z(n18225) );
  NAND U18374 ( .A(b[31]), .B(a[106]), .Z(n18318) );
  ANDN U18375 ( .B(n18084), .A(n18083), .Z(n18087) );
  NAND U18376 ( .A(b[11]), .B(n18085), .Z(n18086) );
  NANDN U18377 ( .A(n18087), .B(n18086), .Z(n18223) );
  XOR U18378 ( .A(n18318), .B(n18223), .Z(n18224) );
  XNOR U18379 ( .A(n18225), .B(n18224), .Z(n18184) );
  NANDN U18380 ( .A(n19116), .B(n18088), .Z(n18090) );
  XOR U18381 ( .A(b[25]), .B(a[114]), .Z(n18214) );
  NANDN U18382 ( .A(n19179), .B(n18214), .Z(n18089) );
  AND U18383 ( .A(n18090), .B(n18089), .Z(n18199) );
  NANDN U18384 ( .A(n18853), .B(n18091), .Z(n18093) );
  XOR U18385 ( .A(b[21]), .B(a[118]), .Z(n18233) );
  NANDN U18386 ( .A(n18926), .B(n18233), .Z(n18092) );
  AND U18387 ( .A(n18093), .B(n18092), .Z(n18197) );
  NANDN U18388 ( .A(n18673), .B(n18094), .Z(n18096) );
  XOR U18389 ( .A(a[120]), .B(b[19]), .Z(n18220) );
  NANDN U18390 ( .A(n18758), .B(n18220), .Z(n18095) );
  NAND U18391 ( .A(n18096), .B(n18095), .Z(n18196) );
  XNOR U18392 ( .A(n18197), .B(n18196), .Z(n18198) );
  XOR U18393 ( .A(n18199), .B(n18198), .Z(n18185) );
  XOR U18394 ( .A(n18184), .B(n18185), .Z(n18187) );
  XOR U18395 ( .A(n18186), .B(n18187), .Z(n18243) );
  NANDN U18396 ( .A(n19394), .B(n18097), .Z(n18099) );
  XOR U18397 ( .A(b[29]), .B(a[110]), .Z(n18226) );
  NANDN U18398 ( .A(n19395), .B(n18226), .Z(n18098) );
  AND U18399 ( .A(n18099), .B(n18098), .Z(n18192) );
  NANDN U18400 ( .A(n18514), .B(n18100), .Z(n18102) );
  XOR U18401 ( .A(a[122]), .B(b[17]), .Z(n18208) );
  NANDN U18402 ( .A(n18585), .B(n18208), .Z(n18101) );
  AND U18403 ( .A(n18102), .B(n18101), .Z(n18191) );
  NANDN U18404 ( .A(n19237), .B(n18103), .Z(n18105) );
  XOR U18405 ( .A(b[27]), .B(a[112]), .Z(n18217) );
  NANDN U18406 ( .A(n19277), .B(n18217), .Z(n18104) );
  NAND U18407 ( .A(n18105), .B(n18104), .Z(n18190) );
  XOR U18408 ( .A(n18191), .B(n18190), .Z(n18193) );
  XOR U18409 ( .A(n18192), .B(n18193), .Z(n18179) );
  NANDN U18410 ( .A(n19005), .B(n18106), .Z(n18108) );
  XOR U18411 ( .A(b[23]), .B(a[116]), .Z(n18239) );
  NANDN U18412 ( .A(n19055), .B(n18239), .Z(n18107) );
  AND U18413 ( .A(n18108), .B(n18107), .Z(n18204) );
  NANDN U18414 ( .A(n18487), .B(n18109), .Z(n18111) );
  XOR U18415 ( .A(a[124]), .B(b[15]), .Z(n18211) );
  NANDN U18416 ( .A(n18311), .B(n18211), .Z(n18110) );
  AND U18417 ( .A(n18111), .B(n18110), .Z(n18203) );
  NANDN U18418 ( .A(n18113), .B(n18112), .Z(n18115) );
  XOR U18419 ( .A(a[126]), .B(b[13]), .Z(n18230) );
  NANDN U18420 ( .A(n18229), .B(n18230), .Z(n18114) );
  NAND U18421 ( .A(n18115), .B(n18114), .Z(n18202) );
  XOR U18422 ( .A(n18203), .B(n18202), .Z(n18205) );
  XNOR U18423 ( .A(n18204), .B(n18205), .Z(n18178) );
  XNOR U18424 ( .A(n18179), .B(n18178), .Z(n18180) );
  NANDN U18425 ( .A(n18117), .B(n18116), .Z(n18121) );
  NANDN U18426 ( .A(n18119), .B(n18118), .Z(n18120) );
  NAND U18427 ( .A(n18121), .B(n18120), .Z(n18181) );
  XNOR U18428 ( .A(n18180), .B(n18181), .Z(n18242) );
  XNOR U18429 ( .A(n18243), .B(n18242), .Z(n18245) );
  NANDN U18430 ( .A(n18123), .B(n18122), .Z(n18127) );
  NANDN U18431 ( .A(n18125), .B(n18124), .Z(n18126) );
  AND U18432 ( .A(n18127), .B(n18126), .Z(n18244) );
  XOR U18433 ( .A(n18245), .B(n18244), .Z(n18174) );
  NANDN U18434 ( .A(n18129), .B(n18128), .Z(n18133) );
  OR U18435 ( .A(n18131), .B(n18130), .Z(n18132) );
  AND U18436 ( .A(n18133), .B(n18132), .Z(n18251) );
  NANDN U18437 ( .A(n18135), .B(n18134), .Z(n18139) );
  NAND U18438 ( .A(n18137), .B(n18136), .Z(n18138) );
  AND U18439 ( .A(n18139), .B(n18138), .Z(n18248) );
  NANDN U18440 ( .A(n18141), .B(n18140), .Z(n18145) );
  OR U18441 ( .A(n18143), .B(n18142), .Z(n18144) );
  NAND U18442 ( .A(n18145), .B(n18144), .Z(n18249) );
  XNOR U18443 ( .A(n18248), .B(n18249), .Z(n18250) );
  XOR U18444 ( .A(n18251), .B(n18250), .Z(n18173) );
  NANDN U18445 ( .A(n18147), .B(n18146), .Z(n18151) );
  NANDN U18446 ( .A(n18149), .B(n18148), .Z(n18150) );
  AND U18447 ( .A(n18151), .B(n18150), .Z(n18172) );
  XOR U18448 ( .A(n18173), .B(n18172), .Z(n18175) );
  XOR U18449 ( .A(n18174), .B(n18175), .Z(n18255) );
  NANDN U18450 ( .A(n18153), .B(n18152), .Z(n18157) );
  NAND U18451 ( .A(n18155), .B(n18154), .Z(n18156) );
  AND U18452 ( .A(n18157), .B(n18156), .Z(n18254) );
  XNOR U18453 ( .A(n18255), .B(n18254), .Z(n18256) );
  XNOR U18454 ( .A(n18257), .B(n18256), .Z(n18260) );
  XNOR U18455 ( .A(n18261), .B(n18260), .Z(n18262) );
  NANDN U18456 ( .A(n18159), .B(n18158), .Z(n18163) );
  OR U18457 ( .A(n18161), .B(n18160), .Z(n18162) );
  NAND U18458 ( .A(n18163), .B(n18162), .Z(n18263) );
  XNOR U18459 ( .A(n18262), .B(n18263), .Z(n18166) );
  XOR U18460 ( .A(n18167), .B(n18166), .Z(n18169) );
  XNOR U18461 ( .A(n18168), .B(n18169), .Z(n18164) );
  XOR U18462 ( .A(n18165), .B(n18164), .Z(c[234]) );
  AND U18463 ( .A(n18165), .B(n18164), .Z(n18267) );
  NANDN U18464 ( .A(n18167), .B(n18166), .Z(n18171) );
  OR U18465 ( .A(n18169), .B(n18168), .Z(n18170) );
  AND U18466 ( .A(n18171), .B(n18170), .Z(n18270) );
  NANDN U18467 ( .A(n18173), .B(n18172), .Z(n18177) );
  OR U18468 ( .A(n18175), .B(n18174), .Z(n18176) );
  AND U18469 ( .A(n18177), .B(n18176), .Z(n18275) );
  NANDN U18470 ( .A(n18179), .B(n18178), .Z(n18183) );
  NANDN U18471 ( .A(n18181), .B(n18180), .Z(n18182) );
  AND U18472 ( .A(n18183), .B(n18182), .Z(n18287) );
  NANDN U18473 ( .A(n18185), .B(n18184), .Z(n18189) );
  OR U18474 ( .A(n18187), .B(n18186), .Z(n18188) );
  AND U18475 ( .A(n18189), .B(n18188), .Z(n18286) );
  XNOR U18476 ( .A(n18287), .B(n18286), .Z(n18289) );
  NANDN U18477 ( .A(n18191), .B(n18190), .Z(n18195) );
  OR U18478 ( .A(n18193), .B(n18192), .Z(n18194) );
  AND U18479 ( .A(n18195), .B(n18194), .Z(n18362) );
  NANDN U18480 ( .A(n18197), .B(n18196), .Z(n18201) );
  NANDN U18481 ( .A(n18199), .B(n18198), .Z(n18200) );
  AND U18482 ( .A(n18201), .B(n18200), .Z(n18360) );
  NANDN U18483 ( .A(n18203), .B(n18202), .Z(n18207) );
  OR U18484 ( .A(n18205), .B(n18204), .Z(n18206) );
  AND U18485 ( .A(n18207), .B(n18206), .Z(n18364) );
  NANDN U18486 ( .A(n18514), .B(n18208), .Z(n18210) );
  XOR U18487 ( .A(a[123]), .B(b[17]), .Z(n18307) );
  NANDN U18488 ( .A(n18585), .B(n18307), .Z(n18209) );
  AND U18489 ( .A(n18210), .B(n18209), .Z(n18332) );
  NANDN U18490 ( .A(n18487), .B(n18211), .Z(n18213) );
  XOR U18491 ( .A(a[125]), .B(b[15]), .Z(n18310) );
  NANDN U18492 ( .A(n18311), .B(n18310), .Z(n18212) );
  AND U18493 ( .A(n18213), .B(n18212), .Z(n18330) );
  NAND U18494 ( .A(n19223), .B(n18214), .Z(n18216) );
  XNOR U18495 ( .A(b[25]), .B(a[115]), .Z(n18314) );
  NANDN U18496 ( .A(n18314), .B(n19224), .Z(n18215) );
  NAND U18497 ( .A(n18216), .B(n18215), .Z(n18355) );
  NAND U18498 ( .A(n19321), .B(n18217), .Z(n18219) );
  XNOR U18499 ( .A(b[27]), .B(a[113]), .Z(n18298) );
  NANDN U18500 ( .A(n18298), .B(n19322), .Z(n18218) );
  NAND U18501 ( .A(n18219), .B(n18218), .Z(n18354) );
  NANDN U18502 ( .A(n18673), .B(n18220), .Z(n18222) );
  XOR U18503 ( .A(a[121]), .B(b[19]), .Z(n18292) );
  NANDN U18504 ( .A(n18758), .B(n18292), .Z(n18221) );
  NAND U18505 ( .A(n18222), .B(n18221), .Z(n18353) );
  XOR U18506 ( .A(n18354), .B(n18353), .Z(n18356) );
  XOR U18507 ( .A(n18355), .B(n18356), .Z(n18329) );
  XNOR U18508 ( .A(n18330), .B(n18329), .Z(n18331) );
  XOR U18509 ( .A(n18332), .B(n18331), .Z(n18363) );
  XOR U18510 ( .A(n18364), .B(n18363), .Z(n18366) );
  NANDN U18511 ( .A(n19394), .B(n18226), .Z(n18228) );
  XOR U18512 ( .A(b[29]), .B(a[111]), .Z(n18301) );
  NANDN U18513 ( .A(n19395), .B(n18301), .Z(n18227) );
  AND U18514 ( .A(n18228), .B(n18227), .Z(n18325) );
  XNOR U18515 ( .A(a[127]), .B(b[13]), .Z(n18346) );
  OR U18516 ( .A(n18346), .B(n18229), .Z(n18232) );
  NAND U18517 ( .A(n18347), .B(n18230), .Z(n18231) );
  AND U18518 ( .A(n18232), .B(n18231), .Z(n18324) );
  NANDN U18519 ( .A(n18853), .B(n18233), .Z(n18235) );
  XOR U18520 ( .A(b[21]), .B(a[119]), .Z(n18295) );
  NANDN U18521 ( .A(n18926), .B(n18295), .Z(n18234) );
  NAND U18522 ( .A(n18235), .B(n18234), .Z(n18323) );
  XOR U18523 ( .A(n18324), .B(n18323), .Z(n18326) );
  XOR U18524 ( .A(n18325), .B(n18326), .Z(n18336) );
  AND U18525 ( .A(b[31]), .B(a[107]), .Z(n18320) );
  XNOR U18526 ( .A(n18319), .B(n18320), .Z(n18317) );
  XOR U18527 ( .A(n18318), .B(n18317), .Z(n18341) );
  NAND U18528 ( .A(n19409), .B(n18236), .Z(n18238) );
  XNOR U18529 ( .A(b[31]), .B(a[109]), .Z(n18350) );
  NANDN U18530 ( .A(n18350), .B(n19411), .Z(n18237) );
  AND U18531 ( .A(n18238), .B(n18237), .Z(n18342) );
  XOR U18532 ( .A(n18341), .B(n18342), .Z(n18343) );
  NAND U18533 ( .A(n19126), .B(n18239), .Z(n18241) );
  XNOR U18534 ( .A(b[23]), .B(a[117]), .Z(n18304) );
  NANDN U18535 ( .A(n18304), .B(n19127), .Z(n18240) );
  NAND U18536 ( .A(n18241), .B(n18240), .Z(n18344) );
  XNOR U18537 ( .A(n18343), .B(n18344), .Z(n18335) );
  XNOR U18538 ( .A(n18336), .B(n18335), .Z(n18337) );
  XOR U18539 ( .A(n18338), .B(n18337), .Z(n18365) );
  XOR U18540 ( .A(n18366), .B(n18365), .Z(n18359) );
  XOR U18541 ( .A(n18360), .B(n18359), .Z(n18361) );
  XOR U18542 ( .A(n18362), .B(n18361), .Z(n18288) );
  XOR U18543 ( .A(n18289), .B(n18288), .Z(n18283) );
  NANDN U18544 ( .A(n18243), .B(n18242), .Z(n18247) );
  NAND U18545 ( .A(n18245), .B(n18244), .Z(n18246) );
  AND U18546 ( .A(n18247), .B(n18246), .Z(n18280) );
  NANDN U18547 ( .A(n18249), .B(n18248), .Z(n18253) );
  NAND U18548 ( .A(n18251), .B(n18250), .Z(n18252) );
  NAND U18549 ( .A(n18253), .B(n18252), .Z(n18281) );
  XNOR U18550 ( .A(n18280), .B(n18281), .Z(n18282) );
  XNOR U18551 ( .A(n18283), .B(n18282), .Z(n18274) );
  XNOR U18552 ( .A(n18275), .B(n18274), .Z(n18277) );
  NANDN U18553 ( .A(n18255), .B(n18254), .Z(n18259) );
  NANDN U18554 ( .A(n18257), .B(n18256), .Z(n18258) );
  AND U18555 ( .A(n18259), .B(n18258), .Z(n18276) );
  XOR U18556 ( .A(n18277), .B(n18276), .Z(n18269) );
  NANDN U18557 ( .A(n18261), .B(n18260), .Z(n18265) );
  NANDN U18558 ( .A(n18263), .B(n18262), .Z(n18264) );
  NAND U18559 ( .A(n18265), .B(n18264), .Z(n18268) );
  XOR U18560 ( .A(n18269), .B(n18268), .Z(n18271) );
  XNOR U18561 ( .A(n18270), .B(n18271), .Z(n18266) );
  XOR U18562 ( .A(n18267), .B(n18266), .Z(c[235]) );
  AND U18563 ( .A(n18267), .B(n18266), .Z(n18370) );
  NANDN U18564 ( .A(n18269), .B(n18268), .Z(n18273) );
  OR U18565 ( .A(n18271), .B(n18270), .Z(n18272) );
  AND U18566 ( .A(n18273), .B(n18272), .Z(n18373) );
  NANDN U18567 ( .A(n18275), .B(n18274), .Z(n18279) );
  NAND U18568 ( .A(n18277), .B(n18276), .Z(n18278) );
  AND U18569 ( .A(n18279), .B(n18278), .Z(n18371) );
  NANDN U18570 ( .A(n18281), .B(n18280), .Z(n18285) );
  NANDN U18571 ( .A(n18283), .B(n18282), .Z(n18284) );
  AND U18572 ( .A(n18285), .B(n18284), .Z(n18379) );
  NANDN U18573 ( .A(n18287), .B(n18286), .Z(n18291) );
  NAND U18574 ( .A(n18289), .B(n18288), .Z(n18290) );
  AND U18575 ( .A(n18291), .B(n18290), .Z(n18378) );
  NANDN U18576 ( .A(n18673), .B(n18292), .Z(n18294) );
  XOR U18577 ( .A(a[122]), .B(b[19]), .Z(n18414) );
  NANDN U18578 ( .A(n18758), .B(n18414), .Z(n18293) );
  AND U18579 ( .A(n18294), .B(n18293), .Z(n18428) );
  NANDN U18580 ( .A(n18853), .B(n18295), .Z(n18297) );
  XOR U18581 ( .A(a[120]), .B(b[21]), .Z(n18417) );
  NANDN U18582 ( .A(n18926), .B(n18417), .Z(n18296) );
  AND U18583 ( .A(n18297), .B(n18296), .Z(n18427) );
  NANDN U18584 ( .A(n18298), .B(n19321), .Z(n18300) );
  XOR U18585 ( .A(b[27]), .B(a[114]), .Z(n18408) );
  NANDN U18586 ( .A(n19277), .B(n18408), .Z(n18299) );
  AND U18587 ( .A(n18300), .B(n18299), .Z(n18435) );
  NANDN U18588 ( .A(n19394), .B(n18301), .Z(n18303) );
  XOR U18589 ( .A(b[29]), .B(a[112]), .Z(n18411) );
  NANDN U18590 ( .A(n19395), .B(n18411), .Z(n18302) );
  AND U18591 ( .A(n18303), .B(n18302), .Z(n18433) );
  NANDN U18592 ( .A(n18304), .B(n19126), .Z(n18306) );
  XOR U18593 ( .A(b[23]), .B(a[118]), .Z(n18405) );
  NANDN U18594 ( .A(n19055), .B(n18405), .Z(n18305) );
  NAND U18595 ( .A(n18306), .B(n18305), .Z(n18432) );
  XNOR U18596 ( .A(n18433), .B(n18432), .Z(n18434) );
  XNOR U18597 ( .A(n18435), .B(n18434), .Z(n18426) );
  XOR U18598 ( .A(n18427), .B(n18426), .Z(n18429) );
  XOR U18599 ( .A(n18428), .B(n18429), .Z(n18451) );
  NANDN U18600 ( .A(n18514), .B(n18307), .Z(n18309) );
  XOR U18601 ( .A(a[124]), .B(b[17]), .Z(n18399) );
  NANDN U18602 ( .A(n18585), .B(n18399), .Z(n18308) );
  AND U18603 ( .A(n18309), .B(n18308), .Z(n18422) );
  NANDN U18604 ( .A(n18487), .B(n18310), .Z(n18313) );
  XOR U18605 ( .A(a[126]), .B(b[15]), .Z(n18438) );
  NANDN U18606 ( .A(n18311), .B(n18438), .Z(n18312) );
  AND U18607 ( .A(n18313), .B(n18312), .Z(n18421) );
  NANDN U18608 ( .A(n18314), .B(n19223), .Z(n18316) );
  XOR U18609 ( .A(b[25]), .B(a[116]), .Z(n18442) );
  NANDN U18610 ( .A(n19179), .B(n18442), .Z(n18315) );
  NAND U18611 ( .A(n18316), .B(n18315), .Z(n18420) );
  XOR U18612 ( .A(n18421), .B(n18420), .Z(n18423) );
  XOR U18613 ( .A(n18422), .B(n18423), .Z(n18449) );
  NANDN U18614 ( .A(n18318), .B(n18317), .Z(n18322) );
  ANDN U18615 ( .B(n18320), .A(n18319), .Z(n18321) );
  ANDN U18616 ( .B(n18322), .A(n18321), .Z(n18448) );
  XNOR U18617 ( .A(n18449), .B(n18448), .Z(n18450) );
  XNOR U18618 ( .A(n18451), .B(n18450), .Z(n18389) );
  NANDN U18619 ( .A(n18324), .B(n18323), .Z(n18328) );
  OR U18620 ( .A(n18326), .B(n18325), .Z(n18327) );
  NAND U18621 ( .A(n18328), .B(n18327), .Z(n18390) );
  XNOR U18622 ( .A(n18389), .B(n18390), .Z(n18391) );
  NANDN U18623 ( .A(n18330), .B(n18329), .Z(n18334) );
  NANDN U18624 ( .A(n18332), .B(n18331), .Z(n18333) );
  NAND U18625 ( .A(n18334), .B(n18333), .Z(n18392) );
  XNOR U18626 ( .A(n18391), .B(n18392), .Z(n18385) );
  NANDN U18627 ( .A(n18336), .B(n18335), .Z(n18340) );
  NAND U18628 ( .A(n18338), .B(n18337), .Z(n18339) );
  AND U18629 ( .A(n18340), .B(n18339), .Z(n18384) );
  NAND U18630 ( .A(b[13]), .B(n18345), .Z(n18349) );
  ANDN U18631 ( .B(n18347), .A(n18346), .Z(n18348) );
  ANDN U18632 ( .B(n18349), .A(n18348), .Z(n18447) );
  NAND U18633 ( .A(b[31]), .B(a[108]), .Z(n18482) );
  NANDN U18634 ( .A(n18350), .B(n19409), .Z(n18352) );
  XOR U18635 ( .A(b[31]), .B(a[110]), .Z(n18402) );
  NANDN U18636 ( .A(n19426), .B(n18402), .Z(n18351) );
  NAND U18637 ( .A(n18352), .B(n18351), .Z(n18445) );
  XOR U18638 ( .A(n18482), .B(n18445), .Z(n18446) );
  XOR U18639 ( .A(n18447), .B(n18446), .Z(n18395) );
  NAND U18640 ( .A(n18354), .B(n18353), .Z(n18358) );
  NAND U18641 ( .A(n18356), .B(n18355), .Z(n18357) );
  AND U18642 ( .A(n18358), .B(n18357), .Z(n18396) );
  XOR U18643 ( .A(n18395), .B(n18396), .Z(n18397) );
  XNOR U18644 ( .A(n18398), .B(n18397), .Z(n18383) );
  XOR U18645 ( .A(n18384), .B(n18383), .Z(n18386) );
  XNOR U18646 ( .A(n18385), .B(n18386), .Z(n18456) );
  NAND U18647 ( .A(n18364), .B(n18363), .Z(n18368) );
  NAND U18648 ( .A(n18366), .B(n18365), .Z(n18367) );
  NAND U18649 ( .A(n18368), .B(n18367), .Z(n18454) );
  XOR U18650 ( .A(n18455), .B(n18454), .Z(n18457) );
  XNOR U18651 ( .A(n18456), .B(n18457), .Z(n18377) );
  XOR U18652 ( .A(n18378), .B(n18377), .Z(n18380) );
  XOR U18653 ( .A(n18379), .B(n18380), .Z(n18372) );
  XOR U18654 ( .A(n18371), .B(n18372), .Z(n18374) );
  XNOR U18655 ( .A(n18373), .B(n18374), .Z(n18369) );
  XOR U18656 ( .A(n18370), .B(n18369), .Z(c[236]) );
  AND U18657 ( .A(n18370), .B(n18369), .Z(n18461) );
  NANDN U18658 ( .A(n18372), .B(n18371), .Z(n18376) );
  OR U18659 ( .A(n18374), .B(n18373), .Z(n18375) );
  AND U18660 ( .A(n18376), .B(n18375), .Z(n18464) );
  NANDN U18661 ( .A(n18378), .B(n18377), .Z(n18382) );
  NANDN U18662 ( .A(n18380), .B(n18379), .Z(n18381) );
  AND U18663 ( .A(n18382), .B(n18381), .Z(n18463) );
  NANDN U18664 ( .A(n18384), .B(n18383), .Z(n18388) );
  NANDN U18665 ( .A(n18386), .B(n18385), .Z(n18387) );
  AND U18666 ( .A(n18388), .B(n18387), .Z(n18550) );
  NANDN U18667 ( .A(n18390), .B(n18389), .Z(n18394) );
  NANDN U18668 ( .A(n18392), .B(n18391), .Z(n18393) );
  AND U18669 ( .A(n18394), .B(n18393), .Z(n18468) );
  XNOR U18670 ( .A(n18468), .B(n18469), .Z(n18470) );
  NANDN U18671 ( .A(n18514), .B(n18399), .Z(n18401) );
  XOR U18672 ( .A(a[125]), .B(b[17]), .Z(n18513) );
  NANDN U18673 ( .A(n18585), .B(n18513), .Z(n18400) );
  AND U18674 ( .A(n18401), .B(n18400), .Z(n18528) );
  NANDN U18675 ( .A(n19425), .B(n18402), .Z(n18404) );
  XOR U18676 ( .A(b[31]), .B(a[111]), .Z(n18491) );
  NANDN U18677 ( .A(n19426), .B(n18491), .Z(n18403) );
  AND U18678 ( .A(n18404), .B(n18403), .Z(n18527) );
  NANDN U18679 ( .A(n19005), .B(n18405), .Z(n18407) );
  XOR U18680 ( .A(b[23]), .B(a[119]), .Z(n18510) );
  NANDN U18681 ( .A(n19055), .B(n18510), .Z(n18406) );
  NAND U18682 ( .A(n18407), .B(n18406), .Z(n18526) );
  XOR U18683 ( .A(n18527), .B(n18526), .Z(n18529) );
  XOR U18684 ( .A(n18528), .B(n18529), .Z(n18477) );
  NANDN U18685 ( .A(n19237), .B(n18408), .Z(n18410) );
  XOR U18686 ( .A(b[27]), .B(a[115]), .Z(n18498) );
  NANDN U18687 ( .A(n19277), .B(n18498), .Z(n18409) );
  AND U18688 ( .A(n18410), .B(n18409), .Z(n18522) );
  NANDN U18689 ( .A(n19394), .B(n18411), .Z(n18413) );
  XOR U18690 ( .A(b[29]), .B(a[113]), .Z(n18501) );
  NANDN U18691 ( .A(n19395), .B(n18501), .Z(n18412) );
  AND U18692 ( .A(n18413), .B(n18412), .Z(n18521) );
  NANDN U18693 ( .A(n18673), .B(n18414), .Z(n18416) );
  XOR U18694 ( .A(a[123]), .B(b[19]), .Z(n18517) );
  NANDN U18695 ( .A(n18758), .B(n18517), .Z(n18415) );
  NAND U18696 ( .A(n18416), .B(n18415), .Z(n18520) );
  XOR U18697 ( .A(n18521), .B(n18520), .Z(n18523) );
  XOR U18698 ( .A(n18522), .B(n18523), .Z(n18475) );
  NAND U18699 ( .A(n18997), .B(n18417), .Z(n18419) );
  XNOR U18700 ( .A(a[121]), .B(b[21]), .Z(n18507) );
  NANDN U18701 ( .A(n18507), .B(n18998), .Z(n18418) );
  AND U18702 ( .A(n18419), .B(n18418), .Z(n18474) );
  XNOR U18703 ( .A(n18475), .B(n18474), .Z(n18476) );
  XNOR U18704 ( .A(n18477), .B(n18476), .Z(n18538) );
  NANDN U18705 ( .A(n18421), .B(n18420), .Z(n18425) );
  OR U18706 ( .A(n18423), .B(n18422), .Z(n18424) );
  NAND U18707 ( .A(n18425), .B(n18424), .Z(n18539) );
  XNOR U18708 ( .A(n18538), .B(n18539), .Z(n18541) );
  NANDN U18709 ( .A(n18427), .B(n18426), .Z(n18431) );
  OR U18710 ( .A(n18429), .B(n18428), .Z(n18430) );
  AND U18711 ( .A(n18431), .B(n18430), .Z(n18540) );
  XOR U18712 ( .A(n18541), .B(n18540), .Z(n18547) );
  NANDN U18713 ( .A(n18433), .B(n18432), .Z(n18437) );
  NANDN U18714 ( .A(n18435), .B(n18434), .Z(n18436) );
  AND U18715 ( .A(n18437), .B(n18436), .Z(n18532) );
  AND U18716 ( .A(b[31]), .B(a[109]), .Z(n18480) );
  XNOR U18717 ( .A(n18481), .B(n18480), .Z(n18483) );
  XOR U18718 ( .A(n18482), .B(n18483), .Z(n18494) );
  NAND U18719 ( .A(n18439), .B(n18438), .Z(n18441) );
  XOR U18720 ( .A(a[127]), .B(b[15]), .Z(n18488) );
  NAND U18721 ( .A(n18486), .B(n18488), .Z(n18440) );
  AND U18722 ( .A(n18441), .B(n18440), .Z(n18495) );
  XOR U18723 ( .A(n18494), .B(n18495), .Z(n18496) );
  NAND U18724 ( .A(n19223), .B(n18442), .Z(n18444) );
  XNOR U18725 ( .A(b[25]), .B(a[117]), .Z(n18504) );
  NANDN U18726 ( .A(n18504), .B(n19224), .Z(n18443) );
  NAND U18727 ( .A(n18444), .B(n18443), .Z(n18497) );
  XOR U18728 ( .A(n18496), .B(n18497), .Z(n18533) );
  XNOR U18729 ( .A(n18532), .B(n18533), .Z(n18535) );
  XOR U18730 ( .A(n18535), .B(n18534), .Z(n18545) );
  NANDN U18731 ( .A(n18449), .B(n18448), .Z(n18453) );
  NANDN U18732 ( .A(n18451), .B(n18450), .Z(n18452) );
  AND U18733 ( .A(n18453), .B(n18452), .Z(n18544) );
  XNOR U18734 ( .A(n18545), .B(n18544), .Z(n18546) );
  XOR U18735 ( .A(n18547), .B(n18546), .Z(n18471) );
  XOR U18736 ( .A(n18470), .B(n18471), .Z(n18551) );
  XNOR U18737 ( .A(n18550), .B(n18551), .Z(n18553) );
  NANDN U18738 ( .A(n18455), .B(n18454), .Z(n18459) );
  NANDN U18739 ( .A(n18457), .B(n18456), .Z(n18458) );
  AND U18740 ( .A(n18459), .B(n18458), .Z(n18552) );
  XNOR U18741 ( .A(n18553), .B(n18552), .Z(n18462) );
  XOR U18742 ( .A(n18463), .B(n18462), .Z(n18465) );
  XNOR U18743 ( .A(n18464), .B(n18465), .Z(n18460) );
  XOR U18744 ( .A(n18461), .B(n18460), .Z(c[237]) );
  AND U18745 ( .A(n18461), .B(n18460), .Z(n18557) );
  NANDN U18746 ( .A(n18463), .B(n18462), .Z(n18467) );
  OR U18747 ( .A(n18465), .B(n18464), .Z(n18466) );
  AND U18748 ( .A(n18467), .B(n18466), .Z(n18560) );
  NANDN U18749 ( .A(n18469), .B(n18468), .Z(n18473) );
  NANDN U18750 ( .A(n18471), .B(n18470), .Z(n18472) );
  AND U18751 ( .A(n18473), .B(n18472), .Z(n18566) );
  NANDN U18752 ( .A(n18475), .B(n18474), .Z(n18479) );
  NANDN U18753 ( .A(n18477), .B(n18476), .Z(n18478) );
  AND U18754 ( .A(n18479), .B(n18478), .Z(n18576) );
  NANDN U18755 ( .A(n18481), .B(n18480), .Z(n18485) );
  ANDN U18756 ( .B(n18483), .A(n18482), .Z(n18484) );
  ANDN U18757 ( .B(n18485), .A(n18484), .Z(n18632) );
  NAND U18758 ( .A(b[15]), .B(n18486), .Z(n18490) );
  ANDN U18759 ( .B(n18488), .A(n18487), .Z(n18489) );
  ANDN U18760 ( .B(n18490), .A(n18489), .Z(n18612) );
  NAND U18761 ( .A(b[31]), .B(a[110]), .Z(n18621) );
  NANDN U18762 ( .A(n19425), .B(n18491), .Z(n18493) );
  XOR U18763 ( .A(b[31]), .B(a[112]), .Z(n18615) );
  NANDN U18764 ( .A(n19426), .B(n18615), .Z(n18492) );
  NAND U18765 ( .A(n18493), .B(n18492), .Z(n18610) );
  XOR U18766 ( .A(n18621), .B(n18610), .Z(n18611) );
  XNOR U18767 ( .A(n18612), .B(n18611), .Z(n18631) );
  XNOR U18768 ( .A(n18632), .B(n18631), .Z(n18633) );
  XOR U18769 ( .A(n18633), .B(n18634), .Z(n18577) );
  XNOR U18770 ( .A(n18576), .B(n18577), .Z(n18579) );
  NANDN U18771 ( .A(n19237), .B(n18498), .Z(n18500) );
  XOR U18772 ( .A(b[27]), .B(a[116]), .Z(n18622) );
  NANDN U18773 ( .A(n19277), .B(n18622), .Z(n18499) );
  AND U18774 ( .A(n18500), .B(n18499), .Z(n18594) );
  NANDN U18775 ( .A(n19394), .B(n18501), .Z(n18503) );
  XOR U18776 ( .A(b[29]), .B(a[114]), .Z(n18625) );
  NANDN U18777 ( .A(n19395), .B(n18625), .Z(n18502) );
  AND U18778 ( .A(n18503), .B(n18502), .Z(n18593) );
  NANDN U18779 ( .A(n18504), .B(n19223), .Z(n18506) );
  XOR U18780 ( .A(b[25]), .B(a[118]), .Z(n18618) );
  NANDN U18781 ( .A(n19179), .B(n18618), .Z(n18505) );
  NAND U18782 ( .A(n18506), .B(n18505), .Z(n18592) );
  XOR U18783 ( .A(n18593), .B(n18592), .Z(n18595) );
  XOR U18784 ( .A(n18594), .B(n18595), .Z(n18606) );
  NANDN U18785 ( .A(n18507), .B(n18997), .Z(n18509) );
  XOR U18786 ( .A(a[122]), .B(b[21]), .Z(n18628) );
  NANDN U18787 ( .A(n18926), .B(n18628), .Z(n18508) );
  AND U18788 ( .A(n18509), .B(n18508), .Z(n18600) );
  NANDN U18789 ( .A(n19005), .B(n18510), .Z(n18512) );
  XOR U18790 ( .A(b[23]), .B(a[120]), .Z(n18589) );
  NANDN U18791 ( .A(n19055), .B(n18589), .Z(n18511) );
  AND U18792 ( .A(n18512), .B(n18511), .Z(n18599) );
  NANDN U18793 ( .A(n18514), .B(n18513), .Z(n18516) );
  XOR U18794 ( .A(a[126]), .B(b[17]), .Z(n18586) );
  NANDN U18795 ( .A(n18585), .B(n18586), .Z(n18515) );
  NAND U18796 ( .A(n18516), .B(n18515), .Z(n18598) );
  XOR U18797 ( .A(n18599), .B(n18598), .Z(n18601) );
  XOR U18798 ( .A(n18600), .B(n18601), .Z(n18605) );
  NAND U18799 ( .A(n18881), .B(n18517), .Z(n18519) );
  XNOR U18800 ( .A(a[124]), .B(b[19]), .Z(n18582) );
  NANDN U18801 ( .A(n18582), .B(n18882), .Z(n18518) );
  AND U18802 ( .A(n18519), .B(n18518), .Z(n18604) );
  XOR U18803 ( .A(n18605), .B(n18604), .Z(n18607) );
  XOR U18804 ( .A(n18606), .B(n18607), .Z(n18640) );
  NANDN U18805 ( .A(n18521), .B(n18520), .Z(n18525) );
  OR U18806 ( .A(n18523), .B(n18522), .Z(n18524) );
  AND U18807 ( .A(n18525), .B(n18524), .Z(n18638) );
  NANDN U18808 ( .A(n18527), .B(n18526), .Z(n18531) );
  OR U18809 ( .A(n18529), .B(n18528), .Z(n18530) );
  NAND U18810 ( .A(n18531), .B(n18530), .Z(n18637) );
  XNOR U18811 ( .A(n18638), .B(n18637), .Z(n18639) );
  XNOR U18812 ( .A(n18640), .B(n18639), .Z(n18578) );
  XOR U18813 ( .A(n18579), .B(n18578), .Z(n18572) );
  NANDN U18814 ( .A(n18533), .B(n18532), .Z(n18537) );
  NAND U18815 ( .A(n18535), .B(n18534), .Z(n18536) );
  AND U18816 ( .A(n18537), .B(n18536), .Z(n18571) );
  NANDN U18817 ( .A(n18539), .B(n18538), .Z(n18543) );
  NAND U18818 ( .A(n18541), .B(n18540), .Z(n18542) );
  NAND U18819 ( .A(n18543), .B(n18542), .Z(n18570) );
  XOR U18820 ( .A(n18571), .B(n18570), .Z(n18573) );
  XOR U18821 ( .A(n18572), .B(n18573), .Z(n18565) );
  NANDN U18822 ( .A(n18545), .B(n18544), .Z(n18549) );
  NANDN U18823 ( .A(n18547), .B(n18546), .Z(n18548) );
  NAND U18824 ( .A(n18549), .B(n18548), .Z(n18564) );
  XOR U18825 ( .A(n18565), .B(n18564), .Z(n18567) );
  XOR U18826 ( .A(n18566), .B(n18567), .Z(n18559) );
  NANDN U18827 ( .A(n18551), .B(n18550), .Z(n18555) );
  NAND U18828 ( .A(n18553), .B(n18552), .Z(n18554) );
  AND U18829 ( .A(n18555), .B(n18554), .Z(n18558) );
  XOR U18830 ( .A(n18559), .B(n18558), .Z(n18561) );
  XNOR U18831 ( .A(n18560), .B(n18561), .Z(n18556) );
  XOR U18832 ( .A(n18557), .B(n18556), .Z(c[238]) );
  AND U18833 ( .A(n18557), .B(n18556), .Z(n18644) );
  NANDN U18834 ( .A(n18559), .B(n18558), .Z(n18563) );
  OR U18835 ( .A(n18561), .B(n18560), .Z(n18562) );
  AND U18836 ( .A(n18563), .B(n18562), .Z(n18647) );
  NANDN U18837 ( .A(n18565), .B(n18564), .Z(n18569) );
  OR U18838 ( .A(n18567), .B(n18566), .Z(n18568) );
  AND U18839 ( .A(n18569), .B(n18568), .Z(n18645) );
  NANDN U18840 ( .A(n18571), .B(n18570), .Z(n18575) );
  OR U18841 ( .A(n18573), .B(n18572), .Z(n18574) );
  AND U18842 ( .A(n18575), .B(n18574), .Z(n18654) );
  NANDN U18843 ( .A(n18577), .B(n18576), .Z(n18581) );
  NAND U18844 ( .A(n18579), .B(n18578), .Z(n18580) );
  AND U18845 ( .A(n18581), .B(n18580), .Z(n18651) );
  NANDN U18846 ( .A(n18582), .B(n18881), .Z(n18584) );
  XOR U18847 ( .A(a[125]), .B(b[19]), .Z(n18672) );
  NANDN U18848 ( .A(n18758), .B(n18672), .Z(n18583) );
  AND U18849 ( .A(n18584), .B(n18583), .Z(n18689) );
  XNOR U18850 ( .A(a[127]), .B(b[17]), .Z(n18682) );
  OR U18851 ( .A(n18682), .B(n18585), .Z(n18588) );
  NAND U18852 ( .A(n18683), .B(n18586), .Z(n18587) );
  AND U18853 ( .A(n18588), .B(n18587), .Z(n18688) );
  NANDN U18854 ( .A(n19005), .B(n18589), .Z(n18591) );
  XOR U18855 ( .A(b[23]), .B(a[121]), .Z(n18711) );
  NANDN U18856 ( .A(n19055), .B(n18711), .Z(n18590) );
  NAND U18857 ( .A(n18591), .B(n18590), .Z(n18687) );
  XOR U18858 ( .A(n18688), .B(n18687), .Z(n18690) );
  XOR U18859 ( .A(n18689), .B(n18690), .Z(n18715) );
  NANDN U18860 ( .A(n18593), .B(n18592), .Z(n18597) );
  OR U18861 ( .A(n18595), .B(n18594), .Z(n18596) );
  AND U18862 ( .A(n18597), .B(n18596), .Z(n18714) );
  XNOR U18863 ( .A(n18715), .B(n18714), .Z(n18717) );
  NANDN U18864 ( .A(n18599), .B(n18598), .Z(n18603) );
  OR U18865 ( .A(n18601), .B(n18600), .Z(n18602) );
  AND U18866 ( .A(n18603), .B(n18602), .Z(n18716) );
  XOR U18867 ( .A(n18717), .B(n18716), .Z(n18728) );
  NANDN U18868 ( .A(n18605), .B(n18604), .Z(n18609) );
  OR U18869 ( .A(n18607), .B(n18606), .Z(n18608) );
  AND U18870 ( .A(n18609), .B(n18608), .Z(n18726) );
  IV U18871 ( .A(n18621), .Z(n18702) );
  NANDN U18872 ( .A(n18702), .B(n18610), .Z(n18614) );
  NANDN U18873 ( .A(n18612), .B(n18611), .Z(n18613) );
  AND U18874 ( .A(n18614), .B(n18613), .Z(n18723) );
  NANDN U18875 ( .A(n19425), .B(n18615), .Z(n18617) );
  XOR U18876 ( .A(b[31]), .B(a[113]), .Z(n18679) );
  NANDN U18877 ( .A(n19426), .B(n18679), .Z(n18616) );
  AND U18878 ( .A(n18617), .B(n18616), .Z(n18664) );
  NANDN U18879 ( .A(n19116), .B(n18618), .Z(n18620) );
  XOR U18880 ( .A(b[25]), .B(a[119]), .Z(n18705) );
  NANDN U18881 ( .A(n19179), .B(n18705), .Z(n18619) );
  NAND U18882 ( .A(n18620), .B(n18619), .Z(n18663) );
  XNOR U18883 ( .A(n18664), .B(n18663), .Z(n18665) );
  AND U18884 ( .A(b[31]), .B(a[111]), .Z(n18699) );
  XOR U18885 ( .A(n18700), .B(n18699), .Z(n18701) );
  XOR U18886 ( .A(n18621), .B(n18701), .Z(n18666) );
  XOR U18887 ( .A(n18665), .B(n18666), .Z(n18720) );
  NANDN U18888 ( .A(n19237), .B(n18622), .Z(n18624) );
  XOR U18889 ( .A(b[27]), .B(a[117]), .Z(n18676) );
  NANDN U18890 ( .A(n19277), .B(n18676), .Z(n18623) );
  AND U18891 ( .A(n18624), .B(n18623), .Z(n18696) );
  NANDN U18892 ( .A(n19394), .B(n18625), .Z(n18627) );
  XOR U18893 ( .A(b[29]), .B(a[115]), .Z(n18708) );
  NANDN U18894 ( .A(n19395), .B(n18708), .Z(n18626) );
  AND U18895 ( .A(n18627), .B(n18626), .Z(n18694) );
  NANDN U18896 ( .A(n18853), .B(n18628), .Z(n18630) );
  XOR U18897 ( .A(a[123]), .B(b[21]), .Z(n18669) );
  NANDN U18898 ( .A(n18926), .B(n18669), .Z(n18629) );
  NAND U18899 ( .A(n18630), .B(n18629), .Z(n18693) );
  XNOR U18900 ( .A(n18694), .B(n18693), .Z(n18695) );
  XOR U18901 ( .A(n18696), .B(n18695), .Z(n18721) );
  XNOR U18902 ( .A(n18720), .B(n18721), .Z(n18722) );
  XOR U18903 ( .A(n18723), .B(n18722), .Z(n18727) );
  XOR U18904 ( .A(n18726), .B(n18727), .Z(n18729) );
  XOR U18905 ( .A(n18728), .B(n18729), .Z(n18660) );
  NANDN U18906 ( .A(n18632), .B(n18631), .Z(n18636) );
  NANDN U18907 ( .A(n18634), .B(n18633), .Z(n18635) );
  AND U18908 ( .A(n18636), .B(n18635), .Z(n18657) );
  NANDN U18909 ( .A(n18638), .B(n18637), .Z(n18642) );
  NANDN U18910 ( .A(n18640), .B(n18639), .Z(n18641) );
  NAND U18911 ( .A(n18642), .B(n18641), .Z(n18658) );
  XNOR U18912 ( .A(n18657), .B(n18658), .Z(n18659) );
  XOR U18913 ( .A(n18660), .B(n18659), .Z(n18652) );
  XNOR U18914 ( .A(n18651), .B(n18652), .Z(n18653) );
  XOR U18915 ( .A(n18654), .B(n18653), .Z(n18646) );
  XOR U18916 ( .A(n18645), .B(n18646), .Z(n18648) );
  XNOR U18917 ( .A(n18647), .B(n18648), .Z(n18643) );
  XOR U18918 ( .A(n18644), .B(n18643), .Z(c[239]) );
  AND U18919 ( .A(n18644), .B(n18643), .Z(n18733) );
  NANDN U18920 ( .A(n18646), .B(n18645), .Z(n18650) );
  OR U18921 ( .A(n18648), .B(n18647), .Z(n18649) );
  AND U18922 ( .A(n18650), .B(n18649), .Z(n18736) );
  NANDN U18923 ( .A(n18652), .B(n18651), .Z(n18656) );
  NANDN U18924 ( .A(n18654), .B(n18653), .Z(n18655) );
  AND U18925 ( .A(n18656), .B(n18655), .Z(n18735) );
  NANDN U18926 ( .A(n18658), .B(n18657), .Z(n18662) );
  NANDN U18927 ( .A(n18660), .B(n18659), .Z(n18661) );
  AND U18928 ( .A(n18662), .B(n18661), .Z(n18743) );
  NANDN U18929 ( .A(n18664), .B(n18663), .Z(n18668) );
  NAND U18930 ( .A(n18666), .B(n18665), .Z(n18667) );
  AND U18931 ( .A(n18668), .B(n18667), .Z(n18753) );
  NANDN U18932 ( .A(n18853), .B(n18669), .Z(n18671) );
  XOR U18933 ( .A(a[124]), .B(b[21]), .Z(n18772) );
  NANDN U18934 ( .A(n18926), .B(n18772), .Z(n18670) );
  AND U18935 ( .A(n18671), .B(n18670), .Z(n18801) );
  NANDN U18936 ( .A(n18673), .B(n18672), .Z(n18675) );
  XOR U18937 ( .A(a[126]), .B(b[19]), .Z(n18759) );
  NANDN U18938 ( .A(n18758), .B(n18759), .Z(n18674) );
  AND U18939 ( .A(n18675), .B(n18674), .Z(n18800) );
  NANDN U18940 ( .A(n19237), .B(n18676), .Z(n18678) );
  XOR U18941 ( .A(b[27]), .B(a[118]), .Z(n18762) );
  NANDN U18942 ( .A(n19277), .B(n18762), .Z(n18677) );
  NAND U18943 ( .A(n18678), .B(n18677), .Z(n18799) );
  XOR U18944 ( .A(n18800), .B(n18799), .Z(n18802) );
  XOR U18945 ( .A(n18801), .B(n18802), .Z(n18788) );
  NANDN U18946 ( .A(n19425), .B(n18679), .Z(n18681) );
  XOR U18947 ( .A(b[31]), .B(a[114]), .Z(n18775) );
  NANDN U18948 ( .A(n19426), .B(n18775), .Z(n18680) );
  AND U18949 ( .A(n18681), .B(n18680), .Z(n18808) );
  NAND U18950 ( .A(b[31]), .B(a[112]), .Z(n18805) );
  ANDN U18951 ( .B(n18683), .A(n18682), .Z(n18686) );
  NAND U18952 ( .A(b[17]), .B(n18684), .Z(n18685) );
  NANDN U18953 ( .A(n18686), .B(n18685), .Z(n18806) );
  XOR U18954 ( .A(n18805), .B(n18806), .Z(n18807) );
  XOR U18955 ( .A(n18808), .B(n18807), .Z(n18787) );
  XNOR U18956 ( .A(n18788), .B(n18787), .Z(n18790) );
  NANDN U18957 ( .A(n18688), .B(n18687), .Z(n18692) );
  OR U18958 ( .A(n18690), .B(n18689), .Z(n18691) );
  AND U18959 ( .A(n18692), .B(n18691), .Z(n18789) );
  XNOR U18960 ( .A(n18790), .B(n18789), .Z(n18752) );
  XNOR U18961 ( .A(n18753), .B(n18752), .Z(n18755) );
  NANDN U18962 ( .A(n18694), .B(n18693), .Z(n18698) );
  NANDN U18963 ( .A(n18696), .B(n18695), .Z(n18697) );
  AND U18964 ( .A(n18698), .B(n18697), .Z(n18796) );
  NANDN U18965 ( .A(n18700), .B(n18699), .Z(n18704) );
  ANDN U18966 ( .B(n18702), .A(n18701), .Z(n18703) );
  ANDN U18967 ( .B(n18704), .A(n18703), .Z(n18794) );
  NANDN U18968 ( .A(n19116), .B(n18705), .Z(n18707) );
  XOR U18969 ( .A(b[25]), .B(a[120]), .Z(n18778) );
  NANDN U18970 ( .A(n19179), .B(n18778), .Z(n18706) );
  AND U18971 ( .A(n18707), .B(n18706), .Z(n18784) );
  NANDN U18972 ( .A(n19394), .B(n18708), .Z(n18710) );
  XOR U18973 ( .A(b[29]), .B(a[116]), .Z(n18766) );
  NANDN U18974 ( .A(n19395), .B(n18766), .Z(n18709) );
  AND U18975 ( .A(n18710), .B(n18709), .Z(n18782) );
  NANDN U18976 ( .A(n19005), .B(n18711), .Z(n18713) );
  XOR U18977 ( .A(a[122]), .B(b[23]), .Z(n18769) );
  NANDN U18978 ( .A(n19055), .B(n18769), .Z(n18712) );
  NAND U18979 ( .A(n18713), .B(n18712), .Z(n18781) );
  XNOR U18980 ( .A(n18782), .B(n18781), .Z(n18783) );
  XNOR U18981 ( .A(n18784), .B(n18783), .Z(n18793) );
  XNOR U18982 ( .A(n18794), .B(n18793), .Z(n18795) );
  XNOR U18983 ( .A(n18796), .B(n18795), .Z(n18754) );
  XOR U18984 ( .A(n18755), .B(n18754), .Z(n18749) );
  NANDN U18985 ( .A(n18715), .B(n18714), .Z(n18719) );
  NAND U18986 ( .A(n18717), .B(n18716), .Z(n18718) );
  AND U18987 ( .A(n18719), .B(n18718), .Z(n18747) );
  NANDN U18988 ( .A(n18721), .B(n18720), .Z(n18725) );
  NANDN U18989 ( .A(n18723), .B(n18722), .Z(n18724) );
  AND U18990 ( .A(n18725), .B(n18724), .Z(n18746) );
  XNOR U18991 ( .A(n18747), .B(n18746), .Z(n18748) );
  XNOR U18992 ( .A(n18749), .B(n18748), .Z(n18740) );
  NANDN U18993 ( .A(n18727), .B(n18726), .Z(n18731) );
  OR U18994 ( .A(n18729), .B(n18728), .Z(n18730) );
  NAND U18995 ( .A(n18731), .B(n18730), .Z(n18741) );
  XNOR U18996 ( .A(n18740), .B(n18741), .Z(n18742) );
  XNOR U18997 ( .A(n18743), .B(n18742), .Z(n18734) );
  XOR U18998 ( .A(n18735), .B(n18734), .Z(n18737) );
  XNOR U18999 ( .A(n18736), .B(n18737), .Z(n18732) );
  XOR U19000 ( .A(n18733), .B(n18732), .Z(c[240]) );
  AND U19001 ( .A(n18733), .B(n18732), .Z(n18812) );
  NANDN U19002 ( .A(n18735), .B(n18734), .Z(n18739) );
  OR U19003 ( .A(n18737), .B(n18736), .Z(n18738) );
  AND U19004 ( .A(n18739), .B(n18738), .Z(n18815) );
  NANDN U19005 ( .A(n18741), .B(n18740), .Z(n18745) );
  NANDN U19006 ( .A(n18743), .B(n18742), .Z(n18744) );
  AND U19007 ( .A(n18745), .B(n18744), .Z(n18814) );
  NANDN U19008 ( .A(n18747), .B(n18746), .Z(n18751) );
  NANDN U19009 ( .A(n18749), .B(n18748), .Z(n18750) );
  AND U19010 ( .A(n18751), .B(n18750), .Z(n18822) );
  NANDN U19011 ( .A(n18753), .B(n18752), .Z(n18757) );
  NAND U19012 ( .A(n18755), .B(n18754), .Z(n18756) );
  AND U19013 ( .A(n18757), .B(n18756), .Z(n18820) );
  XNOR U19014 ( .A(a[127]), .B(b[19]), .Z(n18880) );
  OR U19015 ( .A(n18880), .B(n18758), .Z(n18761) );
  NAND U19016 ( .A(n18881), .B(n18759), .Z(n18760) );
  AND U19017 ( .A(n18761), .B(n18760), .Z(n18866) );
  NANDN U19018 ( .A(n19237), .B(n18762), .Z(n18764) );
  XOR U19019 ( .A(b[27]), .B(a[119]), .Z(n18862) );
  NANDN U19020 ( .A(n19277), .B(n18862), .Z(n18763) );
  NAND U19021 ( .A(n18764), .B(n18763), .Z(n18865) );
  XNOR U19022 ( .A(n18866), .B(n18865), .Z(n18868) );
  IV U19023 ( .A(n18765), .Z(n18872) );
  AND U19024 ( .A(b[31]), .B(a[113]), .Z(n18871) );
  XOR U19025 ( .A(n18872), .B(n18871), .Z(n18873) );
  XOR U19026 ( .A(n18805), .B(n18873), .Z(n18867) );
  XOR U19027 ( .A(n18868), .B(n18867), .Z(n18838) );
  NANDN U19028 ( .A(n19394), .B(n18766), .Z(n18768) );
  XOR U19029 ( .A(b[29]), .B(a[117]), .Z(n18859) );
  NANDN U19030 ( .A(n19395), .B(n18859), .Z(n18767) );
  AND U19031 ( .A(n18768), .B(n18767), .Z(n18887) );
  NANDN U19032 ( .A(n19005), .B(n18769), .Z(n18771) );
  XOR U19033 ( .A(a[123]), .B(b[23]), .Z(n18849) );
  NANDN U19034 ( .A(n19055), .B(n18849), .Z(n18770) );
  AND U19035 ( .A(n18771), .B(n18770), .Z(n18886) );
  NANDN U19036 ( .A(n18853), .B(n18772), .Z(n18774) );
  XOR U19037 ( .A(a[125]), .B(b[21]), .Z(n18852) );
  NANDN U19038 ( .A(n18926), .B(n18852), .Z(n18773) );
  AND U19039 ( .A(n18774), .B(n18773), .Z(n18846) );
  NANDN U19040 ( .A(n19425), .B(n18775), .Z(n18777) );
  XOR U19041 ( .A(b[31]), .B(a[115]), .Z(n18877) );
  NANDN U19042 ( .A(n19426), .B(n18877), .Z(n18776) );
  AND U19043 ( .A(n18777), .B(n18776), .Z(n18844) );
  NANDN U19044 ( .A(n19116), .B(n18778), .Z(n18780) );
  XOR U19045 ( .A(b[25]), .B(a[121]), .Z(n18856) );
  NANDN U19046 ( .A(n19179), .B(n18856), .Z(n18779) );
  NAND U19047 ( .A(n18780), .B(n18779), .Z(n18843) );
  XNOR U19048 ( .A(n18844), .B(n18843), .Z(n18845) );
  XNOR U19049 ( .A(n18846), .B(n18845), .Z(n18885) );
  XOR U19050 ( .A(n18886), .B(n18885), .Z(n18888) );
  XNOR U19051 ( .A(n18887), .B(n18888), .Z(n18837) );
  XNOR U19052 ( .A(n18838), .B(n18837), .Z(n18840) );
  NANDN U19053 ( .A(n18782), .B(n18781), .Z(n18786) );
  NANDN U19054 ( .A(n18784), .B(n18783), .Z(n18785) );
  AND U19055 ( .A(n18786), .B(n18785), .Z(n18839) );
  XOR U19056 ( .A(n18840), .B(n18839), .Z(n18826) );
  NANDN U19057 ( .A(n18788), .B(n18787), .Z(n18792) );
  NAND U19058 ( .A(n18790), .B(n18789), .Z(n18791) );
  AND U19059 ( .A(n18792), .B(n18791), .Z(n18825) );
  XNOR U19060 ( .A(n18826), .B(n18825), .Z(n18827) );
  NANDN U19061 ( .A(n18794), .B(n18793), .Z(n18798) );
  NANDN U19062 ( .A(n18796), .B(n18795), .Z(n18797) );
  AND U19063 ( .A(n18798), .B(n18797), .Z(n18834) );
  NANDN U19064 ( .A(n18800), .B(n18799), .Z(n18804) );
  OR U19065 ( .A(n18802), .B(n18801), .Z(n18803) );
  AND U19066 ( .A(n18804), .B(n18803), .Z(n18832) );
  IV U19067 ( .A(n18805), .Z(n18874) );
  NANDN U19068 ( .A(n18874), .B(n18806), .Z(n18810) );
  NANDN U19069 ( .A(n18808), .B(n18807), .Z(n18809) );
  NAND U19070 ( .A(n18810), .B(n18809), .Z(n18831) );
  XNOR U19071 ( .A(n18832), .B(n18831), .Z(n18833) );
  XOR U19072 ( .A(n18834), .B(n18833), .Z(n18828) );
  XNOR U19073 ( .A(n18827), .B(n18828), .Z(n18819) );
  XNOR U19074 ( .A(n18820), .B(n18819), .Z(n18821) );
  XNOR U19075 ( .A(n18822), .B(n18821), .Z(n18813) );
  XOR U19076 ( .A(n18814), .B(n18813), .Z(n18816) );
  XNOR U19077 ( .A(n18815), .B(n18816), .Z(n18811) );
  XOR U19078 ( .A(n18812), .B(n18811), .Z(c[241]) );
  AND U19079 ( .A(n18812), .B(n18811), .Z(n18892) );
  NANDN U19080 ( .A(n18814), .B(n18813), .Z(n18818) );
  OR U19081 ( .A(n18816), .B(n18815), .Z(n18817) );
  AND U19082 ( .A(n18818), .B(n18817), .Z(n18895) );
  NANDN U19083 ( .A(n18820), .B(n18819), .Z(n18824) );
  NAND U19084 ( .A(n18822), .B(n18821), .Z(n18823) );
  AND U19085 ( .A(n18824), .B(n18823), .Z(n18893) );
  NANDN U19086 ( .A(n18826), .B(n18825), .Z(n18830) );
  NANDN U19087 ( .A(n18828), .B(n18827), .Z(n18829) );
  AND U19088 ( .A(n18830), .B(n18829), .Z(n18901) );
  NANDN U19089 ( .A(n18832), .B(n18831), .Z(n18836) );
  NANDN U19090 ( .A(n18834), .B(n18833), .Z(n18835) );
  AND U19091 ( .A(n18836), .B(n18835), .Z(n18899) );
  NANDN U19092 ( .A(n18838), .B(n18837), .Z(n18842) );
  NAND U19093 ( .A(n18840), .B(n18839), .Z(n18841) );
  AND U19094 ( .A(n18842), .B(n18841), .Z(n18954) );
  NANDN U19095 ( .A(n18844), .B(n18843), .Z(n18848) );
  NANDN U19096 ( .A(n18846), .B(n18845), .Z(n18847) );
  AND U19097 ( .A(n18848), .B(n18847), .Z(n18946) );
  NANDN U19098 ( .A(n19005), .B(n18849), .Z(n18851) );
  XOR U19099 ( .A(a[124]), .B(b[23]), .Z(n18920) );
  NANDN U19100 ( .A(n19055), .B(n18920), .Z(n18850) );
  AND U19101 ( .A(n18851), .B(n18850), .Z(n18936) );
  NANDN U19102 ( .A(n18853), .B(n18852), .Z(n18855) );
  XOR U19103 ( .A(a[126]), .B(b[21]), .Z(n18927) );
  NANDN U19104 ( .A(n18926), .B(n18927), .Z(n18854) );
  AND U19105 ( .A(n18855), .B(n18854), .Z(n18934) );
  NANDN U19106 ( .A(n19116), .B(n18856), .Z(n18858) );
  XOR U19107 ( .A(b[25]), .B(a[122]), .Z(n18917) );
  NANDN U19108 ( .A(n19179), .B(n18917), .Z(n18857) );
  AND U19109 ( .A(n18858), .B(n18857), .Z(n18908) );
  NANDN U19110 ( .A(n19394), .B(n18859), .Z(n18861) );
  XOR U19111 ( .A(b[29]), .B(a[118]), .Z(n18914) );
  NANDN U19112 ( .A(n19395), .B(n18914), .Z(n18860) );
  AND U19113 ( .A(n18861), .B(n18860), .Z(n18906) );
  NANDN U19114 ( .A(n19237), .B(n18862), .Z(n18864) );
  XOR U19115 ( .A(b[27]), .B(a[120]), .Z(n18930) );
  NANDN U19116 ( .A(n19277), .B(n18930), .Z(n18863) );
  NAND U19117 ( .A(n18864), .B(n18863), .Z(n18905) );
  XNOR U19118 ( .A(n18906), .B(n18905), .Z(n18907) );
  XNOR U19119 ( .A(n18908), .B(n18907), .Z(n18933) );
  XNOR U19120 ( .A(n18934), .B(n18933), .Z(n18935) );
  XNOR U19121 ( .A(n18936), .B(n18935), .Z(n18945) );
  XNOR U19122 ( .A(n18946), .B(n18945), .Z(n18948) );
  NANDN U19123 ( .A(n18866), .B(n18865), .Z(n18870) );
  NAND U19124 ( .A(n18868), .B(n18867), .Z(n18869) );
  AND U19125 ( .A(n18870), .B(n18869), .Z(n18942) );
  NANDN U19126 ( .A(n18872), .B(n18871), .Z(n18876) );
  ANDN U19127 ( .B(n18874), .A(n18873), .Z(n18875) );
  ANDN U19128 ( .B(n18876), .A(n18875), .Z(n18940) );
  NANDN U19129 ( .A(n19425), .B(n18877), .Z(n18879) );
  XOR U19130 ( .A(b[31]), .B(a[116]), .Z(n18923) );
  NANDN U19131 ( .A(n19426), .B(n18923), .Z(n18878) );
  AND U19132 ( .A(n18879), .B(n18878), .Z(n18913) );
  NAND U19133 ( .A(b[31]), .B(a[114]), .Z(n18978) );
  ANDN U19134 ( .B(n18881), .A(n18880), .Z(n18884) );
  NAND U19135 ( .A(b[19]), .B(n18882), .Z(n18883) );
  NANDN U19136 ( .A(n18884), .B(n18883), .Z(n18911) );
  XOR U19137 ( .A(n18978), .B(n18911), .Z(n18912) );
  XNOR U19138 ( .A(n18913), .B(n18912), .Z(n18939) );
  XNOR U19139 ( .A(n18940), .B(n18939), .Z(n18941) );
  XNOR U19140 ( .A(n18942), .B(n18941), .Z(n18947) );
  XOR U19141 ( .A(n18948), .B(n18947), .Z(n18952) );
  NANDN U19142 ( .A(n18886), .B(n18885), .Z(n18890) );
  OR U19143 ( .A(n18888), .B(n18887), .Z(n18889) );
  AND U19144 ( .A(n18890), .B(n18889), .Z(n18951) );
  XNOR U19145 ( .A(n18952), .B(n18951), .Z(n18953) );
  XOR U19146 ( .A(n18954), .B(n18953), .Z(n18900) );
  XOR U19147 ( .A(n18899), .B(n18900), .Z(n18902) );
  XOR U19148 ( .A(n18901), .B(n18902), .Z(n18894) );
  XOR U19149 ( .A(n18893), .B(n18894), .Z(n18896) );
  XNOR U19150 ( .A(n18895), .B(n18896), .Z(n18891) );
  XOR U19151 ( .A(n18892), .B(n18891), .Z(c[242]) );
  AND U19152 ( .A(n18892), .B(n18891), .Z(n18958) );
  NANDN U19153 ( .A(n18894), .B(n18893), .Z(n18898) );
  OR U19154 ( .A(n18896), .B(n18895), .Z(n18897) );
  AND U19155 ( .A(n18898), .B(n18897), .Z(n18961) );
  NANDN U19156 ( .A(n18900), .B(n18899), .Z(n18904) );
  NANDN U19157 ( .A(n18902), .B(n18901), .Z(n18903) );
  AND U19158 ( .A(n18904), .B(n18903), .Z(n18960) );
  NANDN U19159 ( .A(n18906), .B(n18905), .Z(n18910) );
  NANDN U19160 ( .A(n18908), .B(n18907), .Z(n18909) );
  AND U19161 ( .A(n18910), .B(n18909), .Z(n19020) );
  XNOR U19162 ( .A(n19020), .B(n19019), .Z(n19022) );
  NANDN U19163 ( .A(n19394), .B(n18914), .Z(n18916) );
  XOR U19164 ( .A(b[29]), .B(a[119]), .Z(n19011) );
  NANDN U19165 ( .A(n19395), .B(n19011), .Z(n18915) );
  AND U19166 ( .A(n18916), .B(n18915), .Z(n19016) );
  NANDN U19167 ( .A(n19116), .B(n18917), .Z(n18919) );
  XOR U19168 ( .A(b[25]), .B(a[123]), .Z(n19001) );
  NANDN U19169 ( .A(n19179), .B(n19001), .Z(n18918) );
  AND U19170 ( .A(n18919), .B(n18918), .Z(n18990) );
  NANDN U19171 ( .A(n19005), .B(n18920), .Z(n18922) );
  XOR U19172 ( .A(a[125]), .B(b[23]), .Z(n19004) );
  NANDN U19173 ( .A(n19055), .B(n19004), .Z(n18921) );
  AND U19174 ( .A(n18922), .B(n18921), .Z(n18988) );
  NANDN U19175 ( .A(n19425), .B(n18923), .Z(n18925) );
  XOR U19176 ( .A(b[31]), .B(a[117]), .Z(n18993) );
  NANDN U19177 ( .A(n19426), .B(n18993), .Z(n18924) );
  NAND U19178 ( .A(n18925), .B(n18924), .Z(n18987) );
  XNOR U19179 ( .A(n18988), .B(n18987), .Z(n18989) );
  XNOR U19180 ( .A(n18990), .B(n18989), .Z(n19015) );
  XNOR U19181 ( .A(n19016), .B(n19015), .Z(n19018) );
  XNOR U19182 ( .A(a[127]), .B(b[21]), .Z(n18996) );
  OR U19183 ( .A(n18996), .B(n18926), .Z(n18929) );
  NAND U19184 ( .A(n18997), .B(n18927), .Z(n18928) );
  AND U19185 ( .A(n18929), .B(n18928), .Z(n18982) );
  NANDN U19186 ( .A(n19237), .B(n18930), .Z(n18932) );
  XOR U19187 ( .A(b[27]), .B(a[121]), .Z(n19008) );
  NANDN U19188 ( .A(n19277), .B(n19008), .Z(n18931) );
  NAND U19189 ( .A(n18932), .B(n18931), .Z(n18981) );
  XNOR U19190 ( .A(n18982), .B(n18981), .Z(n18983) );
  AND U19191 ( .A(b[31]), .B(a[115]), .Z(n18980) );
  XOR U19192 ( .A(n18979), .B(n18980), .Z(n18977) );
  XNOR U19193 ( .A(n18978), .B(n18977), .Z(n18984) );
  XOR U19194 ( .A(n18983), .B(n18984), .Z(n19017) );
  XOR U19195 ( .A(n19018), .B(n19017), .Z(n19021) );
  XOR U19196 ( .A(n19022), .B(n19021), .Z(n18973) );
  NANDN U19197 ( .A(n18934), .B(n18933), .Z(n18938) );
  NANDN U19198 ( .A(n18936), .B(n18935), .Z(n18937) );
  AND U19199 ( .A(n18938), .B(n18937), .Z(n18971) );
  NANDN U19200 ( .A(n18940), .B(n18939), .Z(n18944) );
  NANDN U19201 ( .A(n18942), .B(n18941), .Z(n18943) );
  NAND U19202 ( .A(n18944), .B(n18943), .Z(n18972) );
  XOR U19203 ( .A(n18971), .B(n18972), .Z(n18974) );
  XOR U19204 ( .A(n18973), .B(n18974), .Z(n18966) );
  NANDN U19205 ( .A(n18946), .B(n18945), .Z(n18950) );
  NAND U19206 ( .A(n18948), .B(n18947), .Z(n18949) );
  NAND U19207 ( .A(n18950), .B(n18949), .Z(n18965) );
  XNOR U19208 ( .A(n18966), .B(n18965), .Z(n18968) );
  NANDN U19209 ( .A(n18952), .B(n18951), .Z(n18956) );
  NANDN U19210 ( .A(n18954), .B(n18953), .Z(n18955) );
  AND U19211 ( .A(n18956), .B(n18955), .Z(n18967) );
  XNOR U19212 ( .A(n18968), .B(n18967), .Z(n18959) );
  XOR U19213 ( .A(n18960), .B(n18959), .Z(n18962) );
  XNOR U19214 ( .A(n18961), .B(n18962), .Z(n18957) );
  XOR U19215 ( .A(n18958), .B(n18957), .Z(c[243]) );
  AND U19216 ( .A(n18958), .B(n18957), .Z(n19026) );
  NANDN U19217 ( .A(n18960), .B(n18959), .Z(n18964) );
  OR U19218 ( .A(n18962), .B(n18961), .Z(n18963) );
  AND U19219 ( .A(n18964), .B(n18963), .Z(n19029) );
  NANDN U19220 ( .A(n18966), .B(n18965), .Z(n18970) );
  NAND U19221 ( .A(n18968), .B(n18967), .Z(n18969) );
  AND U19222 ( .A(n18970), .B(n18969), .Z(n19027) );
  NANDN U19223 ( .A(n18972), .B(n18971), .Z(n18976) );
  OR U19224 ( .A(n18974), .B(n18973), .Z(n18975) );
  AND U19225 ( .A(n18976), .B(n18975), .Z(n19036) );
  NANDN U19226 ( .A(n18982), .B(n18981), .Z(n18986) );
  NAND U19227 ( .A(n18984), .B(n18983), .Z(n18985) );
  NAND U19228 ( .A(n18986), .B(n18985), .Z(n19038) );
  XNOR U19229 ( .A(n19037), .B(n19038), .Z(n19040) );
  NANDN U19230 ( .A(n18988), .B(n18987), .Z(n18992) );
  NANDN U19231 ( .A(n18990), .B(n18989), .Z(n18991) );
  AND U19232 ( .A(n18992), .B(n18991), .Z(n19039) );
  XOR U19233 ( .A(n19040), .B(n19039), .Z(n19081) );
  NANDN U19234 ( .A(n19425), .B(n18993), .Z(n18995) );
  XOR U19235 ( .A(b[31]), .B(a[118]), .Z(n19069) );
  NANDN U19236 ( .A(n19426), .B(n19069), .Z(n18994) );
  AND U19237 ( .A(n18995), .B(n18994), .Z(n19075) );
  NAND U19238 ( .A(b[31]), .B(a[116]), .Z(n19107) );
  ANDN U19239 ( .B(n18997), .A(n18996), .Z(n19000) );
  NAND U19240 ( .A(b[21]), .B(n18998), .Z(n18999) );
  NANDN U19241 ( .A(n19000), .B(n18999), .Z(n19072) );
  XOR U19242 ( .A(n19107), .B(n19072), .Z(n19074) );
  XOR U19243 ( .A(n19075), .B(n19074), .Z(n19045) );
  NANDN U19244 ( .A(n19116), .B(n19001), .Z(n19003) );
  XOR U19245 ( .A(a[124]), .B(b[25]), .Z(n19062) );
  NANDN U19246 ( .A(n19179), .B(n19062), .Z(n19002) );
  AND U19247 ( .A(n19003), .B(n19002), .Z(n19051) );
  NANDN U19248 ( .A(n19005), .B(n19004), .Z(n19007) );
  XOR U19249 ( .A(a[126]), .B(b[23]), .Z(n19056) );
  NANDN U19250 ( .A(n19055), .B(n19056), .Z(n19006) );
  AND U19251 ( .A(n19007), .B(n19006), .Z(n19050) );
  NANDN U19252 ( .A(n19237), .B(n19008), .Z(n19010) );
  XOR U19253 ( .A(b[27]), .B(a[122]), .Z(n19059) );
  NANDN U19254 ( .A(n19277), .B(n19059), .Z(n19009) );
  NAND U19255 ( .A(n19010), .B(n19009), .Z(n19049) );
  XOR U19256 ( .A(n19050), .B(n19049), .Z(n19052) );
  XOR U19257 ( .A(n19051), .B(n19052), .Z(n19044) );
  NAND U19258 ( .A(n19065), .B(n19011), .Z(n19014) );
  XNOR U19259 ( .A(b[29]), .B(a[120]), .Z(n19066) );
  NANDN U19260 ( .A(n19066), .B(n19012), .Z(n19013) );
  AND U19261 ( .A(n19014), .B(n19013), .Z(n19043) );
  XOR U19262 ( .A(n19044), .B(n19043), .Z(n19046) );
  XOR U19263 ( .A(n19045), .B(n19046), .Z(n19078) );
  XOR U19264 ( .A(n19078), .B(n19079), .Z(n19080) );
  XOR U19265 ( .A(n19081), .B(n19080), .Z(n19033) );
  NANDN U19266 ( .A(n19020), .B(n19019), .Z(n19024) );
  NAND U19267 ( .A(n19022), .B(n19021), .Z(n19023) );
  AND U19268 ( .A(n19024), .B(n19023), .Z(n19034) );
  XOR U19269 ( .A(n19033), .B(n19034), .Z(n19035) );
  XOR U19270 ( .A(n19036), .B(n19035), .Z(n19028) );
  XOR U19271 ( .A(n19027), .B(n19028), .Z(n19030) );
  XNOR U19272 ( .A(n19029), .B(n19030), .Z(n19025) );
  XOR U19273 ( .A(n19026), .B(n19025), .Z(c[244]) );
  AND U19274 ( .A(n19026), .B(n19025), .Z(n19083) );
  NANDN U19275 ( .A(n19028), .B(n19027), .Z(n19032) );
  OR U19276 ( .A(n19030), .B(n19029), .Z(n19031) );
  AND U19277 ( .A(n19032), .B(n19031), .Z(n19086) );
  NANDN U19278 ( .A(n19038), .B(n19037), .Z(n19042) );
  NAND U19279 ( .A(n19040), .B(n19039), .Z(n19041) );
  AND U19280 ( .A(n19042), .B(n19041), .Z(n19091) );
  NANDN U19281 ( .A(n19044), .B(n19043), .Z(n19048) );
  NANDN U19282 ( .A(n19046), .B(n19045), .Z(n19047) );
  AND U19283 ( .A(n19048), .B(n19047), .Z(n19099) );
  NANDN U19284 ( .A(n19050), .B(n19049), .Z(n19054) );
  OR U19285 ( .A(n19052), .B(n19051), .Z(n19053) );
  AND U19286 ( .A(n19054), .B(n19053), .Z(n19138) );
  XNOR U19287 ( .A(a[127]), .B(b[23]), .Z(n19125) );
  OR U19288 ( .A(n19125), .B(n19055), .Z(n19058) );
  NAND U19289 ( .A(n19126), .B(n19056), .Z(n19057) );
  AND U19290 ( .A(n19058), .B(n19057), .Z(n19103) );
  NANDN U19291 ( .A(n19237), .B(n19059), .Z(n19061) );
  XOR U19292 ( .A(b[27]), .B(a[123]), .Z(n19112) );
  NANDN U19293 ( .A(n19277), .B(n19112), .Z(n19060) );
  NAND U19294 ( .A(n19061), .B(n19060), .Z(n19102) );
  XNOR U19295 ( .A(n19103), .B(n19102), .Z(n19105) );
  IV U19296 ( .A(n19107), .Z(n19073) );
  XOR U19297 ( .A(n19106), .B(n19073), .Z(n19109) );
  AND U19298 ( .A(b[31]), .B(a[117]), .Z(n19108) );
  XOR U19299 ( .A(n19109), .B(n19108), .Z(n19104) );
  XOR U19300 ( .A(n19105), .B(n19104), .Z(n19136) );
  NANDN U19301 ( .A(n19116), .B(n19062), .Z(n19064) );
  XOR U19302 ( .A(a[125]), .B(b[25]), .Z(n19115) );
  NANDN U19303 ( .A(n19179), .B(n19115), .Z(n19063) );
  AND U19304 ( .A(n19064), .B(n19063), .Z(n19133) );
  NANDN U19305 ( .A(n19066), .B(n19065), .Z(n19068) );
  XOR U19306 ( .A(b[29]), .B(a[121]), .Z(n19119) );
  NANDN U19307 ( .A(n19395), .B(n19119), .Z(n19067) );
  AND U19308 ( .A(n19068), .B(n19067), .Z(n19131) );
  NANDN U19309 ( .A(n19425), .B(n19069), .Z(n19071) );
  XOR U19310 ( .A(b[31]), .B(a[119]), .Z(n19122) );
  NANDN U19311 ( .A(n19426), .B(n19122), .Z(n19070) );
  NAND U19312 ( .A(n19071), .B(n19070), .Z(n19130) );
  XNOR U19313 ( .A(n19131), .B(n19130), .Z(n19132) );
  XOR U19314 ( .A(n19133), .B(n19132), .Z(n19137) );
  XOR U19315 ( .A(n19136), .B(n19137), .Z(n19139) );
  XOR U19316 ( .A(n19138), .B(n19139), .Z(n19097) );
  NANDN U19317 ( .A(n19073), .B(n19072), .Z(n19077) );
  NANDN U19318 ( .A(n19075), .B(n19074), .Z(n19076) );
  AND U19319 ( .A(n19077), .B(n19076), .Z(n19096) );
  XNOR U19320 ( .A(n19097), .B(n19096), .Z(n19098) );
  XNOR U19321 ( .A(n19099), .B(n19098), .Z(n19090) );
  XNOR U19322 ( .A(n19091), .B(n19090), .Z(n19092) );
  XNOR U19323 ( .A(n19092), .B(n19093), .Z(n19084) );
  XOR U19324 ( .A(n19085), .B(n19084), .Z(n19087) );
  XNOR U19325 ( .A(n19086), .B(n19087), .Z(n19082) );
  XOR U19326 ( .A(n19083), .B(n19082), .Z(c[245]) );
  AND U19327 ( .A(n19083), .B(n19082), .Z(n19143) );
  NANDN U19328 ( .A(n19085), .B(n19084), .Z(n19089) );
  OR U19329 ( .A(n19087), .B(n19086), .Z(n19088) );
  AND U19330 ( .A(n19089), .B(n19088), .Z(n19146) );
  NANDN U19331 ( .A(n19091), .B(n19090), .Z(n19095) );
  NANDN U19332 ( .A(n19093), .B(n19092), .Z(n19094) );
  AND U19333 ( .A(n19095), .B(n19094), .Z(n19145) );
  NANDN U19334 ( .A(n19097), .B(n19096), .Z(n19101) );
  NANDN U19335 ( .A(n19099), .B(n19098), .Z(n19100) );
  AND U19336 ( .A(n19101), .B(n19100), .Z(n19153) );
  NANDN U19337 ( .A(n19107), .B(n19106), .Z(n19111) );
  NAND U19338 ( .A(n19109), .B(n19108), .Z(n19110) );
  NAND U19339 ( .A(n19111), .B(n19110), .Z(n19157) );
  XNOR U19340 ( .A(n19156), .B(n19157), .Z(n19158) );
  NANDN U19341 ( .A(n19237), .B(n19112), .Z(n19114) );
  XOR U19342 ( .A(b[27]), .B(a[124]), .Z(n19176) );
  NANDN U19343 ( .A(n19277), .B(n19176), .Z(n19113) );
  AND U19344 ( .A(n19114), .B(n19113), .Z(n19164) );
  NANDN U19345 ( .A(n19116), .B(n19115), .Z(n19118) );
  XOR U19346 ( .A(a[126]), .B(b[25]), .Z(n19180) );
  NANDN U19347 ( .A(n19179), .B(n19180), .Z(n19117) );
  AND U19348 ( .A(n19118), .B(n19117), .Z(n19163) );
  NANDN U19349 ( .A(n19394), .B(n19119), .Z(n19121) );
  XOR U19350 ( .A(b[29]), .B(a[122]), .Z(n19183) );
  NANDN U19351 ( .A(n19395), .B(n19183), .Z(n19120) );
  NAND U19352 ( .A(n19121), .B(n19120), .Z(n19162) );
  XOR U19353 ( .A(n19163), .B(n19162), .Z(n19165) );
  XOR U19354 ( .A(n19164), .B(n19165), .Z(n19188) );
  NANDN U19355 ( .A(n19425), .B(n19122), .Z(n19124) );
  XOR U19356 ( .A(b[31]), .B(a[120]), .Z(n19173) );
  NANDN U19357 ( .A(n19426), .B(n19173), .Z(n19123) );
  AND U19358 ( .A(n19124), .B(n19123), .Z(n19170) );
  NAND U19359 ( .A(b[31]), .B(a[118]), .Z(n19186) );
  ANDN U19360 ( .B(n19126), .A(n19125), .Z(n19129) );
  NAND U19361 ( .A(b[23]), .B(n19127), .Z(n19128) );
  NANDN U19362 ( .A(n19129), .B(n19128), .Z(n19168) );
  XOR U19363 ( .A(n19186), .B(n19168), .Z(n19169) );
  XOR U19364 ( .A(n19170), .B(n19169), .Z(n19187) );
  XNOR U19365 ( .A(n19188), .B(n19187), .Z(n19189) );
  NANDN U19366 ( .A(n19131), .B(n19130), .Z(n19135) );
  NANDN U19367 ( .A(n19133), .B(n19132), .Z(n19134) );
  NAND U19368 ( .A(n19135), .B(n19134), .Z(n19190) );
  XOR U19369 ( .A(n19189), .B(n19190), .Z(n19159) );
  XNOR U19370 ( .A(n19158), .B(n19159), .Z(n19150) );
  NANDN U19371 ( .A(n19137), .B(n19136), .Z(n19141) );
  OR U19372 ( .A(n19139), .B(n19138), .Z(n19140) );
  NAND U19373 ( .A(n19141), .B(n19140), .Z(n19151) );
  XNOR U19374 ( .A(n19150), .B(n19151), .Z(n19152) );
  XNOR U19375 ( .A(n19153), .B(n19152), .Z(n19144) );
  XOR U19376 ( .A(n19145), .B(n19144), .Z(n19147) );
  XNOR U19377 ( .A(n19146), .B(n19147), .Z(n19142) );
  XOR U19378 ( .A(n19143), .B(n19142), .Z(c[246]) );
  AND U19379 ( .A(n19143), .B(n19142), .Z(n19194) );
  NANDN U19380 ( .A(n19145), .B(n19144), .Z(n19149) );
  OR U19381 ( .A(n19147), .B(n19146), .Z(n19148) );
  AND U19382 ( .A(n19149), .B(n19148), .Z(n19197) );
  NANDN U19383 ( .A(n19151), .B(n19150), .Z(n19155) );
  NANDN U19384 ( .A(n19153), .B(n19152), .Z(n19154) );
  AND U19385 ( .A(n19155), .B(n19154), .Z(n19196) );
  NANDN U19386 ( .A(n19157), .B(n19156), .Z(n19161) );
  NANDN U19387 ( .A(n19159), .B(n19158), .Z(n19160) );
  AND U19388 ( .A(n19161), .B(n19160), .Z(n19204) );
  NANDN U19389 ( .A(n19163), .B(n19162), .Z(n19167) );
  OR U19390 ( .A(n19165), .B(n19164), .Z(n19166) );
  AND U19391 ( .A(n19167), .B(n19166), .Z(n19209) );
  IV U19392 ( .A(n19186), .Z(n19230) );
  NANDN U19393 ( .A(n19230), .B(n19168), .Z(n19172) );
  NANDN U19394 ( .A(n19170), .B(n19169), .Z(n19171) );
  AND U19395 ( .A(n19172), .B(n19171), .Z(n19208) );
  NANDN U19396 ( .A(n19425), .B(n19173), .Z(n19175) );
  XOR U19397 ( .A(b[31]), .B(a[121]), .Z(n19219) );
  NANDN U19398 ( .A(n19426), .B(n19219), .Z(n19174) );
  AND U19399 ( .A(n19175), .B(n19174), .Z(n19243) );
  NANDN U19400 ( .A(n19237), .B(n19176), .Z(n19178) );
  XOR U19401 ( .A(b[27]), .B(a[125]), .Z(n19236) );
  NANDN U19402 ( .A(n19277), .B(n19236), .Z(n19177) );
  AND U19403 ( .A(n19178), .B(n19177), .Z(n19241) );
  XNOR U19404 ( .A(a[127]), .B(b[25]), .Z(n19222) );
  OR U19405 ( .A(n19222), .B(n19179), .Z(n19182) );
  NAND U19406 ( .A(n19223), .B(n19180), .Z(n19181) );
  AND U19407 ( .A(n19182), .B(n19181), .Z(n19214) );
  NANDN U19408 ( .A(n19394), .B(n19183), .Z(n19185) );
  XOR U19409 ( .A(b[29]), .B(a[123]), .Z(n19233) );
  NANDN U19410 ( .A(n19395), .B(n19233), .Z(n19184) );
  NAND U19411 ( .A(n19185), .B(n19184), .Z(n19213) );
  XNOR U19412 ( .A(n19214), .B(n19213), .Z(n19215) );
  AND U19413 ( .A(b[31]), .B(a[119]), .Z(n19227) );
  XOR U19414 ( .A(n19228), .B(n19227), .Z(n19229) );
  XOR U19415 ( .A(n19186), .B(n19229), .Z(n19216) );
  XOR U19416 ( .A(n19215), .B(n19216), .Z(n19240) );
  XNOR U19417 ( .A(n19241), .B(n19240), .Z(n19242) );
  XNOR U19418 ( .A(n19243), .B(n19242), .Z(n19207) );
  XOR U19419 ( .A(n19208), .B(n19207), .Z(n19210) );
  XOR U19420 ( .A(n19209), .B(n19210), .Z(n19202) );
  NANDN U19421 ( .A(n19188), .B(n19187), .Z(n19192) );
  NANDN U19422 ( .A(n19190), .B(n19189), .Z(n19191) );
  NAND U19423 ( .A(n19192), .B(n19191), .Z(n19201) );
  XNOR U19424 ( .A(n19202), .B(n19201), .Z(n19203) );
  XNOR U19425 ( .A(n19204), .B(n19203), .Z(n19195) );
  XOR U19426 ( .A(n19196), .B(n19195), .Z(n19198) );
  XNOR U19427 ( .A(n19197), .B(n19198), .Z(n19193) );
  XOR U19428 ( .A(n19194), .B(n19193), .Z(c[247]) );
  AND U19429 ( .A(n19194), .B(n19193), .Z(n19247) );
  NANDN U19430 ( .A(n19196), .B(n19195), .Z(n19200) );
  OR U19431 ( .A(n19198), .B(n19197), .Z(n19199) );
  AND U19432 ( .A(n19200), .B(n19199), .Z(n19250) );
  NANDN U19433 ( .A(n19202), .B(n19201), .Z(n19206) );
  NANDN U19434 ( .A(n19204), .B(n19203), .Z(n19205) );
  AND U19435 ( .A(n19206), .B(n19205), .Z(n19249) );
  NANDN U19436 ( .A(n19208), .B(n19207), .Z(n19212) );
  OR U19437 ( .A(n19210), .B(n19209), .Z(n19211) );
  AND U19438 ( .A(n19212), .B(n19211), .Z(n19256) );
  NANDN U19439 ( .A(n19214), .B(n19213), .Z(n19218) );
  NAND U19440 ( .A(n19216), .B(n19215), .Z(n19217) );
  AND U19441 ( .A(n19218), .B(n19217), .Z(n19261) );
  NANDN U19442 ( .A(n19425), .B(n19219), .Z(n19221) );
  XOR U19443 ( .A(b[31]), .B(a[122]), .Z(n19284) );
  NANDN U19444 ( .A(n19426), .B(n19284), .Z(n19220) );
  AND U19445 ( .A(n19221), .B(n19220), .Z(n19274) );
  NAND U19446 ( .A(b[31]), .B(a[120]), .Z(n19287) );
  ANDN U19447 ( .B(n19223), .A(n19222), .Z(n19226) );
  NAND U19448 ( .A(b[25]), .B(n19224), .Z(n19225) );
  NANDN U19449 ( .A(n19226), .B(n19225), .Z(n19272) );
  XOR U19450 ( .A(n19287), .B(n19272), .Z(n19273) );
  XNOR U19451 ( .A(n19274), .B(n19273), .Z(n19260) );
  XNOR U19452 ( .A(n19261), .B(n19260), .Z(n19263) );
  NANDN U19453 ( .A(n19228), .B(n19227), .Z(n19232) );
  ANDN U19454 ( .B(n19230), .A(n19229), .Z(n19231) );
  ANDN U19455 ( .B(n19232), .A(n19231), .Z(n19269) );
  NANDN U19456 ( .A(n19394), .B(n19233), .Z(n19235) );
  XOR U19457 ( .A(b[29]), .B(a[124]), .Z(n19281) );
  NANDN U19458 ( .A(n19395), .B(n19281), .Z(n19234) );
  AND U19459 ( .A(n19235), .B(n19234), .Z(n19267) );
  NANDN U19460 ( .A(n19237), .B(n19236), .Z(n19239) );
  XOR U19461 ( .A(a[126]), .B(b[27]), .Z(n19278) );
  NANDN U19462 ( .A(n19277), .B(n19278), .Z(n19238) );
  NAND U19463 ( .A(n19239), .B(n19238), .Z(n19266) );
  XNOR U19464 ( .A(n19267), .B(n19266), .Z(n19268) );
  XNOR U19465 ( .A(n19269), .B(n19268), .Z(n19262) );
  XOR U19466 ( .A(n19263), .B(n19262), .Z(n19255) );
  NANDN U19467 ( .A(n19241), .B(n19240), .Z(n19245) );
  NANDN U19468 ( .A(n19243), .B(n19242), .Z(n19244) );
  AND U19469 ( .A(n19245), .B(n19244), .Z(n19254) );
  XOR U19470 ( .A(n19255), .B(n19254), .Z(n19257) );
  XNOR U19471 ( .A(n19256), .B(n19257), .Z(n19248) );
  XOR U19472 ( .A(n19249), .B(n19248), .Z(n19251) );
  XNOR U19473 ( .A(n19250), .B(n19251), .Z(n19246) );
  XOR U19474 ( .A(n19247), .B(n19246), .Z(c[248]) );
  AND U19475 ( .A(n19247), .B(n19246), .Z(n19289) );
  NANDN U19476 ( .A(n19249), .B(n19248), .Z(n19253) );
  OR U19477 ( .A(n19251), .B(n19250), .Z(n19252) );
  AND U19478 ( .A(n19253), .B(n19252), .Z(n19292) );
  NANDN U19479 ( .A(n19255), .B(n19254), .Z(n19259) );
  NANDN U19480 ( .A(n19257), .B(n19256), .Z(n19258) );
  AND U19481 ( .A(n19259), .B(n19258), .Z(n19291) );
  NANDN U19482 ( .A(n19261), .B(n19260), .Z(n19265) );
  NAND U19483 ( .A(n19263), .B(n19262), .Z(n19264) );
  AND U19484 ( .A(n19265), .B(n19264), .Z(n19327) );
  NANDN U19485 ( .A(n19267), .B(n19266), .Z(n19271) );
  NANDN U19486 ( .A(n19269), .B(n19268), .Z(n19270) );
  AND U19487 ( .A(n19271), .B(n19270), .Z(n19326) );
  IV U19488 ( .A(n19287), .Z(n19312) );
  NANDN U19489 ( .A(n19312), .B(n19272), .Z(n19276) );
  NANDN U19490 ( .A(n19274), .B(n19273), .Z(n19275) );
  AND U19491 ( .A(n19276), .B(n19275), .Z(n19299) );
  XNOR U19492 ( .A(a[127]), .B(b[27]), .Z(n19320) );
  OR U19493 ( .A(n19320), .B(n19277), .Z(n19280) );
  NAND U19494 ( .A(n19321), .B(n19278), .Z(n19279) );
  AND U19495 ( .A(n19280), .B(n19279), .Z(n19297) );
  NANDN U19496 ( .A(n19394), .B(n19281), .Z(n19283) );
  XOR U19497 ( .A(b[29]), .B(a[125]), .Z(n19308) );
  NANDN U19498 ( .A(n19395), .B(n19308), .Z(n19282) );
  AND U19499 ( .A(n19283), .B(n19282), .Z(n19303) );
  NANDN U19500 ( .A(n19425), .B(n19284), .Z(n19286) );
  XOR U19501 ( .A(b[31]), .B(a[123]), .Z(n19317) );
  NANDN U19502 ( .A(n19426), .B(n19317), .Z(n19285) );
  NAND U19503 ( .A(n19286), .B(n19285), .Z(n19302) );
  XNOR U19504 ( .A(n19303), .B(n19302), .Z(n19304) );
  AND U19505 ( .A(b[31]), .B(a[121]), .Z(n19313) );
  XOR U19506 ( .A(n19314), .B(n19313), .Z(n19311) );
  XOR U19507 ( .A(n19287), .B(n19311), .Z(n19305) );
  XOR U19508 ( .A(n19304), .B(n19305), .Z(n19296) );
  XNOR U19509 ( .A(n19297), .B(n19296), .Z(n19298) );
  XNOR U19510 ( .A(n19299), .B(n19298), .Z(n19325) );
  XOR U19511 ( .A(n19326), .B(n19325), .Z(n19328) );
  XNOR U19512 ( .A(n19327), .B(n19328), .Z(n19290) );
  XOR U19513 ( .A(n19291), .B(n19290), .Z(n19293) );
  XNOR U19514 ( .A(n19292), .B(n19293), .Z(n19288) );
  XOR U19515 ( .A(n19289), .B(n19288), .Z(c[249]) );
  AND U19516 ( .A(n19289), .B(n19288), .Z(n19332) );
  NANDN U19517 ( .A(n19291), .B(n19290), .Z(n19295) );
  OR U19518 ( .A(n19293), .B(n19292), .Z(n19294) );
  AND U19519 ( .A(n19295), .B(n19294), .Z(n19335) );
  NANDN U19520 ( .A(n19297), .B(n19296), .Z(n19301) );
  NANDN U19521 ( .A(n19299), .B(n19298), .Z(n19300) );
  AND U19522 ( .A(n19301), .B(n19300), .Z(n19341) );
  NANDN U19523 ( .A(n19303), .B(n19302), .Z(n19307) );
  NAND U19524 ( .A(n19305), .B(n19304), .Z(n19306) );
  AND U19525 ( .A(n19307), .B(n19306), .Z(n19340) );
  NANDN U19526 ( .A(n19394), .B(n19308), .Z(n19310) );
  XOR U19527 ( .A(b[29]), .B(a[126]), .Z(n19354) );
  NANDN U19528 ( .A(n19395), .B(n19354), .Z(n19309) );
  AND U19529 ( .A(n19310), .B(n19309), .Z(n19346) );
  ANDN U19530 ( .B(n19312), .A(n19311), .Z(n19316) );
  NANDN U19531 ( .A(n19314), .B(n19313), .Z(n19315) );
  NANDN U19532 ( .A(n19316), .B(n19315), .Z(n19345) );
  XNOR U19533 ( .A(n19346), .B(n19345), .Z(n19347) );
  NANDN U19534 ( .A(n19425), .B(n19317), .Z(n19319) );
  XOR U19535 ( .A(b[31]), .B(a[124]), .Z(n19351) );
  NANDN U19536 ( .A(n19426), .B(n19351), .Z(n19318) );
  AND U19537 ( .A(n19319), .B(n19318), .Z(n19361) );
  NAND U19538 ( .A(b[31]), .B(a[122]), .Z(n19358) );
  ANDN U19539 ( .B(n19321), .A(n19320), .Z(n19324) );
  NAND U19540 ( .A(b[27]), .B(n19322), .Z(n19323) );
  NANDN U19541 ( .A(n19324), .B(n19323), .Z(n19359) );
  XOR U19542 ( .A(n19358), .B(n19359), .Z(n19360) );
  XOR U19543 ( .A(n19361), .B(n19360), .Z(n19348) );
  XNOR U19544 ( .A(n19347), .B(n19348), .Z(n19339) );
  XOR U19545 ( .A(n19340), .B(n19339), .Z(n19342) );
  XOR U19546 ( .A(n19341), .B(n19342), .Z(n19334) );
  NANDN U19547 ( .A(n19326), .B(n19325), .Z(n19330) );
  OR U19548 ( .A(n19328), .B(n19327), .Z(n19329) );
  AND U19549 ( .A(n19330), .B(n19329), .Z(n19333) );
  XOR U19550 ( .A(n19334), .B(n19333), .Z(n19336) );
  XNOR U19551 ( .A(n19335), .B(n19336), .Z(n19331) );
  XOR U19552 ( .A(n19332), .B(n19331), .Z(c[250]) );
  AND U19553 ( .A(n19332), .B(n19331), .Z(n19365) );
  NANDN U19554 ( .A(n19334), .B(n19333), .Z(n19338) );
  OR U19555 ( .A(n19336), .B(n19335), .Z(n19337) );
  AND U19556 ( .A(n19338), .B(n19337), .Z(n19368) );
  NANDN U19557 ( .A(n19340), .B(n19339), .Z(n19344) );
  OR U19558 ( .A(n19342), .B(n19341), .Z(n19343) );
  AND U19559 ( .A(n19344), .B(n19343), .Z(n19366) );
  NANDN U19560 ( .A(n19346), .B(n19345), .Z(n19350) );
  NANDN U19561 ( .A(n19348), .B(n19347), .Z(n19349) );
  AND U19562 ( .A(n19350), .B(n19349), .Z(n19374) );
  NANDN U19563 ( .A(n19425), .B(n19351), .Z(n19353) );
  XOR U19564 ( .A(b[31]), .B(a[125]), .Z(n19390) );
  NANDN U19565 ( .A(n19426), .B(n19390), .Z(n19352) );
  AND U19566 ( .A(n19353), .B(n19352), .Z(n19379) );
  NANDN U19567 ( .A(n19394), .B(n19354), .Z(n19356) );
  XOR U19568 ( .A(a[127]), .B(b[29]), .Z(n19393) );
  NANDN U19569 ( .A(n19395), .B(n19393), .Z(n19355) );
  NAND U19570 ( .A(n19356), .B(n19355), .Z(n19378) );
  XNOR U19571 ( .A(n19379), .B(n19378), .Z(n19381) );
  IV U19572 ( .A(n19357), .Z(n19385) );
  AND U19573 ( .A(b[31]), .B(a[123]), .Z(n19384) );
  XOR U19574 ( .A(n19385), .B(n19384), .Z(n19386) );
  XOR U19575 ( .A(n19358), .B(n19386), .Z(n19380) );
  XOR U19576 ( .A(n19381), .B(n19380), .Z(n19373) );
  IV U19577 ( .A(n19358), .Z(n19387) );
  NANDN U19578 ( .A(n19387), .B(n19359), .Z(n19363) );
  NANDN U19579 ( .A(n19361), .B(n19360), .Z(n19362) );
  AND U19580 ( .A(n19363), .B(n19362), .Z(n19372) );
  XOR U19581 ( .A(n19373), .B(n19372), .Z(n19375) );
  XOR U19582 ( .A(n19374), .B(n19375), .Z(n19367) );
  XOR U19583 ( .A(n19366), .B(n19367), .Z(n19369) );
  XNOR U19584 ( .A(n19368), .B(n19369), .Z(n19364) );
  XOR U19585 ( .A(n19365), .B(n19364), .Z(c[251]) );
  AND U19586 ( .A(n19365), .B(n19364), .Z(n19399) );
  NANDN U19587 ( .A(n19367), .B(n19366), .Z(n19371) );
  OR U19588 ( .A(n19369), .B(n19368), .Z(n19370) );
  AND U19589 ( .A(n19371), .B(n19370), .Z(n19402) );
  NANDN U19590 ( .A(n19373), .B(n19372), .Z(n19377) );
  NANDN U19591 ( .A(n19375), .B(n19374), .Z(n19376) );
  AND U19592 ( .A(n19377), .B(n19376), .Z(n19401) );
  NANDN U19593 ( .A(n19379), .B(n19378), .Z(n19383) );
  NAND U19594 ( .A(n19381), .B(n19380), .Z(n19382) );
  AND U19595 ( .A(n19383), .B(n19382), .Z(n19416) );
  NANDN U19596 ( .A(n19385), .B(n19384), .Z(n19389) );
  ANDN U19597 ( .B(n19387), .A(n19386), .Z(n19388) );
  ANDN U19598 ( .B(n19389), .A(n19388), .Z(n19415) );
  NAND U19599 ( .A(n19409), .B(n19390), .Z(n19392) );
  XNOR U19600 ( .A(b[31]), .B(a[126]), .Z(n19410) );
  NANDN U19601 ( .A(n19410), .B(n19411), .Z(n19391) );
  NAND U19602 ( .A(n19392), .B(n19391), .Z(n19407) );
  NAND U19603 ( .A(b[31]), .B(a[124]), .Z(n19422) );
  NANDN U19604 ( .A(n19394), .B(n19393), .Z(n19397) );
  NANDN U19605 ( .A(n19395), .B(b[29]), .Z(n19396) );
  NAND U19606 ( .A(n19397), .B(n19396), .Z(n19406) );
  XOR U19607 ( .A(n19422), .B(n19406), .Z(n19408) );
  XOR U19608 ( .A(n19407), .B(n19408), .Z(n19414) );
  XOR U19609 ( .A(n19415), .B(n19414), .Z(n19417) );
  XNOR U19610 ( .A(n19416), .B(n19417), .Z(n19400) );
  XOR U19611 ( .A(n19401), .B(n19400), .Z(n19403) );
  XNOR U19612 ( .A(n19402), .B(n19403), .Z(n19398) );
  XOR U19613 ( .A(n19399), .B(n19398), .Z(c[252]) );
  AND U19614 ( .A(n19399), .B(n19398), .Z(n19430) );
  NANDN U19615 ( .A(n19401), .B(n19400), .Z(n19405) );
  OR U19616 ( .A(n19403), .B(n19402), .Z(n19404) );
  AND U19617 ( .A(n19405), .B(n19404), .Z(n19440) );
  NANDN U19618 ( .A(n19410), .B(n19409), .Z(n19413) );
  XOR U19619 ( .A(a[127]), .B(b[31]), .Z(n19424) );
  NAND U19620 ( .A(n19411), .B(n19424), .Z(n19412) );
  NAND U19621 ( .A(n19413), .B(n19412), .Z(n19431) );
  AND U19622 ( .A(b[31]), .B(a[125]), .Z(n19421) );
  XOR U19623 ( .A(n19420), .B(n19421), .Z(n19423) );
  XOR U19624 ( .A(n19423), .B(n19422), .Z(n19432) );
  XOR U19625 ( .A(n19431), .B(n19432), .Z(n19434) );
  XOR U19626 ( .A(n19433), .B(n19434), .Z(n19437) );
  NANDN U19627 ( .A(n19415), .B(n19414), .Z(n19419) );
  OR U19628 ( .A(n19417), .B(n19416), .Z(n19418) );
  AND U19629 ( .A(n19419), .B(n19418), .Z(n19438) );
  XOR U19630 ( .A(n19437), .B(n19438), .Z(n19439) );
  XOR U19631 ( .A(n19440), .B(n19439), .Z(n19429) );
  XOR U19632 ( .A(n19430), .B(n19429), .Z(c[253]) );
  AND U19633 ( .A(b[31]), .B(a[126]), .Z(n19444) );
  NANDN U19634 ( .A(n19425), .B(n19424), .Z(n19428) );
  NANDN U19635 ( .A(n19426), .B(b[31]), .Z(n19427) );
  NAND U19636 ( .A(n19428), .B(n19427), .Z(n19445) );
  XNOR U19637 ( .A(n19444), .B(n19445), .Z(n19447) );
  XOR U19638 ( .A(n19446), .B(n19447), .Z(n19450) );
  AND U19639 ( .A(n19430), .B(n19429), .Z(n19449) );
  XNOR U19640 ( .A(n19450), .B(n19449), .Z(n19442) );
  NANDN U19641 ( .A(n19432), .B(n19431), .Z(n19436) );
  NANDN U19642 ( .A(n19434), .B(n19433), .Z(n19435) );
  AND U19643 ( .A(n19436), .B(n19435), .Z(n19451) );
  IV U19644 ( .A(n19452), .Z(n19448) );
  XOR U19645 ( .A(n19451), .B(n19448), .Z(n19441) );
  XNOR U19646 ( .A(n19442), .B(n19441), .Z(c[254]) );
endmodule

