
module hamming_N16000_CC128_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;

  XOR U1 ( .A(A[9]), .B(n1), .Z(SUM[9]) );
  XOR U2 ( .A(A[8]), .B(n2), .Z(SUM[8]) );
  XNOR U3 ( .A(A[7]), .B(n3), .Z(SUM[7]) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  XOR U16 ( .A(A[13]), .B(n16), .Z(SUM[13]) );
  ANDN U17 ( .B(A[12]), .A(n17), .Z(n16) );
  XNOR U18 ( .A(A[12]), .B(n17), .Z(SUM[12]) );
  NANDN U19 ( .A(n18), .B(A[11]), .Z(n17) );
  XNOR U20 ( .A(A[11]), .B(n18), .Z(SUM[11]) );
  NAND U21 ( .A(n19), .B(A[10]), .Z(n18) );
  XOR U22 ( .A(A[10]), .B(n19), .Z(SUM[10]) );
  AND U23 ( .A(A[9]), .B(n1), .Z(n19) );
  AND U24 ( .A(n2), .B(A[8]), .Z(n1) );
  ANDN U25 ( .B(A[7]), .A(n3), .Z(n2) );
  AND U26 ( .A(n20), .B(n21), .Z(n3) );
  NAND U27 ( .A(n22), .B(B[6]), .Z(n21) );
  NANDN U28 ( .A(A[6]), .B(n4), .Z(n22) );
  NANDN U29 ( .A(n4), .B(A[6]), .Z(n20) );
  AND U30 ( .A(n23), .B(n24), .Z(n4) );
  NAND U31 ( .A(n25), .B(B[5]), .Z(n24) );
  NANDN U32 ( .A(A[5]), .B(n6), .Z(n25) );
  NANDN U33 ( .A(n6), .B(A[5]), .Z(n23) );
  AND U34 ( .A(n26), .B(n27), .Z(n6) );
  NAND U35 ( .A(n28), .B(B[4]), .Z(n27) );
  NANDN U36 ( .A(A[4]), .B(n8), .Z(n28) );
  NANDN U37 ( .A(n8), .B(A[4]), .Z(n26) );
  AND U38 ( .A(n29), .B(n30), .Z(n8) );
  NAND U39 ( .A(n31), .B(B[3]), .Z(n30) );
  NANDN U40 ( .A(A[3]), .B(n10), .Z(n31) );
  NANDN U41 ( .A(n10), .B(A[3]), .Z(n29) );
  AND U42 ( .A(n32), .B(n33), .Z(n10) );
  NAND U43 ( .A(n34), .B(B[2]), .Z(n33) );
  NANDN U44 ( .A(A[2]), .B(n12), .Z(n34) );
  NANDN U45 ( .A(n12), .B(A[2]), .Z(n32) );
  AND U46 ( .A(n35), .B(n36), .Z(n12) );
  NAND U47 ( .A(n37), .B(B[1]), .Z(n36) );
  OR U48 ( .A(n14), .B(A[1]), .Z(n37) );
  NAND U49 ( .A(n14), .B(A[1]), .Z(n35) );
  AND U50 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U51 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC128_DW01_add_1 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;

  IV U1 ( .A(B[6]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n1), .Z(SUM[6]) );
  AND U3 ( .A(n3), .B(n4), .Z(n2) );
  NAND U4 ( .A(n5), .B(B[5]), .Z(n4) );
  NANDN U5 ( .A(A[5]), .B(n6), .Z(n5) );
  NANDN U6 ( .A(n6), .B(A[5]), .Z(n3) );
  XOR U7 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n7) );
  AND U9 ( .A(n8), .B(n9), .Z(n6) );
  NAND U10 ( .A(n10), .B(B[4]), .Z(n9) );
  NANDN U11 ( .A(A[4]), .B(n11), .Z(n10) );
  NANDN U12 ( .A(n11), .B(A[4]), .Z(n8) );
  XOR U13 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U14 ( .A(B[4]), .B(A[4]), .Z(n12) );
  AND U15 ( .A(n13), .B(n14), .Z(n11) );
  NAND U16 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U17 ( .A(A[3]), .B(n16), .Z(n15) );
  NANDN U18 ( .A(n16), .B(A[3]), .Z(n13) );
  XOR U19 ( .A(n16), .B(n17), .Z(SUM[3]) );
  XNOR U20 ( .A(B[3]), .B(A[3]), .Z(n17) );
  AND U21 ( .A(n18), .B(n19), .Z(n16) );
  NAND U22 ( .A(n20), .B(B[2]), .Z(n19) );
  NANDN U23 ( .A(A[2]), .B(n21), .Z(n20) );
  NANDN U24 ( .A(n21), .B(A[2]), .Z(n18) );
  XOR U25 ( .A(n21), .B(n22), .Z(SUM[2]) );
  XNOR U26 ( .A(B[2]), .B(A[2]), .Z(n22) );
  AND U27 ( .A(n23), .B(n24), .Z(n21) );
  NAND U28 ( .A(n25), .B(B[1]), .Z(n24) );
  OR U29 ( .A(n26), .B(A[1]), .Z(n25) );
  NAND U30 ( .A(n26), .B(A[1]), .Z(n23) );
  XOR U31 ( .A(n26), .B(n27), .Z(SUM[1]) );
  XOR U32 ( .A(B[1]), .B(A[1]), .Z(n27) );
  AND U33 ( .A(B[0]), .B(A[0]), .Z(n26) );
  XOR U34 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC128_DW01_add_2 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC128_DW01_add_3 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC128_DW01_add_4 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC128_DW01_add_5 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  AND U1 ( .A(n3), .B(B[4]), .Z(SUM[5]) );
  IV U2 ( .A(B[4]), .Z(n2) );
  IV U3 ( .A(n4), .Z(n3) );
  XOR U4 ( .A(n4), .B(n2), .Z(SUM[4]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[3]), .Z(n6) );
  NANDN U7 ( .A(A[3]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[3]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U10 ( .A(B[3]), .B(A[3]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[2]), .Z(n11) );
  NANDN U13 ( .A(A[2]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[2]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[1]), .Z(n16) );
  OR U19 ( .A(n18), .B(A[1]), .Z(n17) );
  NAND U20 ( .A(n18), .B(A[1]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U22 ( .A(B[1]), .B(A[1]), .Z(n19) );
  AND U23 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U24 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC128 ( clk, rst, x, y, o );
  input [124:0] x;
  input [124:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N482, N483, N484, N485, N489, N490, N491, N492, N493, N496, N497,
         N498, N499, N500, N503, N504, N505, N506, N507, N510, N511, N512,
         N513, N514, N517, N518, N519, N520, N521, N524, N525, N526, N527,
         N528, N529, N531, N532, N533, N534, N535, N536, N538, N539, N540,
         N541, N542, N543, N545, N546, N547, N548, N549, N550, N551, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850;
  wire   [6:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC128_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, olocal}), .CI(1'b0), .SUM(o) );
  hamming_N16000_CC128_DW01_add_1 add_42_root_add_47_I125 ( .A({1'b0, N543, 
        N542, N541, N540, N539, N538}), .B({N551, N550, N549, N548, N547, N546, 
        N545}), .CI(1'b0), .SUM(olocal) );
  hamming_N16000_CC128_DW01_add_2 add_43_root_add_47_I125 ( .A({1'b0, N529, 
        N528, N527, N526, N525, N524}), .B({1'b0, N536, N535, N534, N533, N532, 
        N531}), .CI(1'b0), .SUM({N551, N550, N549, N548, N547, N546, N545}) );
  hamming_N16000_CC128_DW01_add_3 add_44_root_add_47_I125 ( .A({1'b0, 1'b0, 
        N514, N513, N512, N511, N510}), .B({1'b0, 1'b0, N521, N520, N519, N518, 
        N517}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, N543, N542, N541, 
        N540, N539, N538}) );
  hamming_N16000_CC128_DW01_add_4 add_45_root_add_47_I125 ( .A({1'b0, 1'b0, 
        N500, N499, N498, N497, N496}), .B({1'b0, 1'b0, N507, N506, N505, N504, 
        N503}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__1, N536, N535, N534, 
        N533, N532, N531}) );
  hamming_N16000_CC128_DW01_add_5 add_46_root_add_47_I125 ( .A({1'b0, 1'b0, 
        1'b0, N485, N484, N483, N482}), .B({1'b0, 1'b0, N493, N492, N491, N490, 
        N489}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__2, N529, N528, N527, 
        N526, N525, N524}) );
  NAND U228 ( .A(n104), .B(n105), .Z(N521) );
  NANDN U229 ( .A(n106), .B(n107), .Z(n105) );
  OR U230 ( .A(n108), .B(n109), .Z(n107) );
  NAND U231 ( .A(n108), .B(n109), .Z(n104) );
  XOR U232 ( .A(n108), .B(n110), .Z(N520) );
  XNOR U233 ( .A(n106), .B(n109), .Z(n110) );
  AND U234 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U235 ( .A(n113), .B(n114), .Z(n112) );
  NANDN U236 ( .A(n115), .B(n116), .Z(n114) );
  NANDN U237 ( .A(n116), .B(n115), .Z(n111) );
  NAND U238 ( .A(n117), .B(n118), .Z(n106) );
  NANDN U239 ( .A(n119), .B(n120), .Z(n118) );
  OR U240 ( .A(n121), .B(n122), .Z(n120) );
  NAND U241 ( .A(n122), .B(n121), .Z(n117) );
  AND U242 ( .A(n123), .B(n124), .Z(n108) );
  NANDN U243 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U244 ( .A(n127), .B(n128), .Z(n126) );
  NANDN U245 ( .A(n128), .B(n127), .Z(n123) );
  XOR U246 ( .A(n122), .B(n129), .Z(N519) );
  XOR U247 ( .A(n119), .B(n121), .Z(n129) );
  XNOR U248 ( .A(n115), .B(n130), .Z(n121) );
  XNOR U249 ( .A(n113), .B(n116), .Z(n130) );
  NAND U250 ( .A(n131), .B(n132), .Z(n116) );
  NAND U251 ( .A(n133), .B(n134), .Z(n132) );
  OR U252 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U253 ( .A(n137), .B(n135), .Z(n131) );
  IV U254 ( .A(n136), .Z(n137) );
  NAND U255 ( .A(n138), .B(n139), .Z(n113) );
  NAND U256 ( .A(n140), .B(n141), .Z(n139) );
  NANDN U257 ( .A(n142), .B(n143), .Z(n140) );
  NANDN U258 ( .A(n143), .B(n142), .Z(n138) );
  AND U259 ( .A(n144), .B(n145), .Z(n115) );
  NAND U260 ( .A(n146), .B(n147), .Z(n145) );
  OR U261 ( .A(n148), .B(n149), .Z(n146) );
  NANDN U262 ( .A(n150), .B(n148), .Z(n144) );
  NAND U263 ( .A(n151), .B(n152), .Z(n119) );
  NANDN U264 ( .A(n153), .B(n154), .Z(n152) );
  OR U265 ( .A(n155), .B(n156), .Z(n154) );
  NANDN U266 ( .A(n157), .B(n155), .Z(n151) );
  IV U267 ( .A(n156), .Z(n157) );
  XNOR U268 ( .A(n127), .B(n158), .Z(n122) );
  XNOR U269 ( .A(n125), .B(n128), .Z(n158) );
  NAND U270 ( .A(n159), .B(n160), .Z(n128) );
  NAND U271 ( .A(n161), .B(n162), .Z(n160) );
  OR U272 ( .A(n163), .B(n164), .Z(n161) );
  NANDN U273 ( .A(n165), .B(n163), .Z(n159) );
  IV U274 ( .A(n164), .Z(n165) );
  NAND U275 ( .A(n166), .B(n167), .Z(n125) );
  NAND U276 ( .A(n168), .B(n169), .Z(n167) );
  NANDN U277 ( .A(n170), .B(n171), .Z(n168) );
  NANDN U278 ( .A(n171), .B(n170), .Z(n166) );
  AND U279 ( .A(n172), .B(n173), .Z(n127) );
  NAND U280 ( .A(n174), .B(n175), .Z(n173) );
  OR U281 ( .A(n176), .B(n177), .Z(n174) );
  NANDN U282 ( .A(n178), .B(n176), .Z(n172) );
  XNOR U283 ( .A(n153), .B(n179), .Z(N518) );
  XOR U284 ( .A(n155), .B(n156), .Z(n179) );
  XNOR U285 ( .A(n169), .B(n180), .Z(n156) );
  XOR U286 ( .A(n170), .B(n171), .Z(n180) );
  XOR U287 ( .A(n176), .B(n181), .Z(n171) );
  XOR U288 ( .A(n175), .B(n178), .Z(n181) );
  IV U289 ( .A(n177), .Z(n178) );
  NAND U290 ( .A(n182), .B(n183), .Z(n177) );
  OR U291 ( .A(n184), .B(n185), .Z(n183) );
  OR U292 ( .A(n186), .B(n187), .Z(n182) );
  NAND U293 ( .A(n188), .B(n189), .Z(n175) );
  OR U294 ( .A(n190), .B(n191), .Z(n189) );
  OR U295 ( .A(n192), .B(n193), .Z(n188) );
  NOR U296 ( .A(n194), .B(n195), .Z(n176) );
  ANDN U297 ( .B(n196), .A(n197), .Z(n170) );
  XNOR U298 ( .A(n163), .B(n198), .Z(n169) );
  XNOR U299 ( .A(n162), .B(n164), .Z(n198) );
  NAND U300 ( .A(n199), .B(n200), .Z(n164) );
  OR U301 ( .A(n201), .B(n202), .Z(n200) );
  OR U302 ( .A(n203), .B(n204), .Z(n199) );
  NAND U303 ( .A(n205), .B(n206), .Z(n162) );
  OR U304 ( .A(n207), .B(n208), .Z(n206) );
  OR U305 ( .A(n209), .B(n210), .Z(n205) );
  ANDN U306 ( .B(n211), .A(n212), .Z(n163) );
  IV U307 ( .A(n213), .Z(n211) );
  ANDN U308 ( .B(n214), .A(n215), .Z(n155) );
  XOR U309 ( .A(n141), .B(n216), .Z(n153) );
  XOR U310 ( .A(n142), .B(n143), .Z(n216) );
  XOR U311 ( .A(n148), .B(n217), .Z(n143) );
  XOR U312 ( .A(n147), .B(n150), .Z(n217) );
  IV U313 ( .A(n149), .Z(n150) );
  NAND U314 ( .A(n218), .B(n219), .Z(n149) );
  OR U315 ( .A(n220), .B(n221), .Z(n219) );
  OR U316 ( .A(n222), .B(n223), .Z(n218) );
  NAND U317 ( .A(n224), .B(n225), .Z(n147) );
  OR U318 ( .A(n226), .B(n227), .Z(n225) );
  OR U319 ( .A(n228), .B(n229), .Z(n224) );
  NOR U320 ( .A(n230), .B(n231), .Z(n148) );
  ANDN U321 ( .B(n232), .A(n233), .Z(n142) );
  IV U322 ( .A(n234), .Z(n232) );
  XNOR U323 ( .A(n135), .B(n235), .Z(n141) );
  XNOR U324 ( .A(n134), .B(n136), .Z(n235) );
  NAND U325 ( .A(n236), .B(n237), .Z(n136) );
  OR U326 ( .A(n238), .B(n239), .Z(n237) );
  OR U327 ( .A(n240), .B(n241), .Z(n236) );
  NAND U328 ( .A(n242), .B(n243), .Z(n134) );
  OR U329 ( .A(n244), .B(n245), .Z(n243) );
  OR U330 ( .A(n246), .B(n247), .Z(n242) );
  ANDN U331 ( .B(n248), .A(n249), .Z(n135) );
  IV U332 ( .A(n250), .Z(n248) );
  XNOR U333 ( .A(n215), .B(n214), .Z(N517) );
  XOR U334 ( .A(n234), .B(n233), .Z(n214) );
  XNOR U335 ( .A(n249), .B(n250), .Z(n233) );
  XNOR U336 ( .A(n244), .B(n245), .Z(n250) );
  XNOR U337 ( .A(n246), .B(n247), .Z(n245) );
  XNOR U338 ( .A(y[103]), .B(x[103]), .Z(n247) );
  XNOR U339 ( .A(y[104]), .B(x[104]), .Z(n246) );
  XNOR U340 ( .A(y[102]), .B(x[102]), .Z(n244) );
  XNOR U341 ( .A(n238), .B(n239), .Z(n249) );
  XNOR U342 ( .A(y[99]), .B(x[99]), .Z(n239) );
  XNOR U343 ( .A(n240), .B(n241), .Z(n238) );
  XNOR U344 ( .A(y[100]), .B(x[100]), .Z(n241) );
  XNOR U345 ( .A(y[101]), .B(x[101]), .Z(n240) );
  XNOR U346 ( .A(n231), .B(n230), .Z(n234) );
  XNOR U347 ( .A(n226), .B(n227), .Z(n230) );
  XNOR U348 ( .A(y[96]), .B(x[96]), .Z(n227) );
  XNOR U349 ( .A(n228), .B(n229), .Z(n226) );
  XNOR U350 ( .A(y[97]), .B(x[97]), .Z(n229) );
  XNOR U351 ( .A(y[98]), .B(x[98]), .Z(n228) );
  XNOR U352 ( .A(n220), .B(n221), .Z(n231) );
  XNOR U353 ( .A(y[93]), .B(x[93]), .Z(n221) );
  XNOR U354 ( .A(n222), .B(n223), .Z(n220) );
  XNOR U355 ( .A(y[94]), .B(x[94]), .Z(n223) );
  XNOR U356 ( .A(y[95]), .B(x[95]), .Z(n222) );
  XOR U357 ( .A(n196), .B(n197), .Z(n215) );
  XNOR U358 ( .A(n212), .B(n213), .Z(n197) );
  XNOR U359 ( .A(n207), .B(n208), .Z(n213) );
  XNOR U360 ( .A(n209), .B(n210), .Z(n208) );
  XNOR U361 ( .A(y[91]), .B(x[91]), .Z(n210) );
  XNOR U362 ( .A(y[92]), .B(x[92]), .Z(n209) );
  XNOR U363 ( .A(y[90]), .B(x[90]), .Z(n207) );
  XNOR U364 ( .A(n201), .B(n202), .Z(n212) );
  XNOR U365 ( .A(y[87]), .B(x[87]), .Z(n202) );
  XNOR U366 ( .A(n203), .B(n204), .Z(n201) );
  XNOR U367 ( .A(y[88]), .B(x[88]), .Z(n204) );
  XNOR U368 ( .A(y[89]), .B(x[89]), .Z(n203) );
  XOR U369 ( .A(n195), .B(n194), .Z(n196) );
  XNOR U370 ( .A(n190), .B(n191), .Z(n194) );
  XNOR U371 ( .A(y[84]), .B(x[84]), .Z(n191) );
  XNOR U372 ( .A(n192), .B(n193), .Z(n190) );
  XNOR U373 ( .A(y[85]), .B(x[85]), .Z(n193) );
  XNOR U374 ( .A(y[86]), .B(x[86]), .Z(n192) );
  XNOR U375 ( .A(n184), .B(n185), .Z(n195) );
  XNOR U376 ( .A(y[81]), .B(x[81]), .Z(n185) );
  XNOR U377 ( .A(n186), .B(n187), .Z(n184) );
  XNOR U378 ( .A(y[82]), .B(x[82]), .Z(n187) );
  XNOR U379 ( .A(y[83]), .B(x[83]), .Z(n186) );
  NAND U380 ( .A(n251), .B(n252), .Z(N514) );
  NANDN U381 ( .A(n253), .B(n254), .Z(n252) );
  OR U382 ( .A(n255), .B(n256), .Z(n254) );
  NAND U383 ( .A(n255), .B(n256), .Z(n251) );
  XOR U384 ( .A(n255), .B(n257), .Z(N513) );
  XNOR U385 ( .A(n253), .B(n256), .Z(n257) );
  AND U386 ( .A(n258), .B(n259), .Z(n256) );
  NANDN U387 ( .A(n260), .B(n261), .Z(n259) );
  NANDN U388 ( .A(n262), .B(n263), .Z(n261) );
  NANDN U389 ( .A(n263), .B(n262), .Z(n258) );
  NAND U390 ( .A(n264), .B(n265), .Z(n253) );
  NANDN U391 ( .A(n266), .B(n267), .Z(n265) );
  OR U392 ( .A(n268), .B(n269), .Z(n267) );
  NAND U393 ( .A(n269), .B(n268), .Z(n264) );
  AND U394 ( .A(n270), .B(n271), .Z(n255) );
  NANDN U395 ( .A(n272), .B(n273), .Z(n271) );
  NANDN U396 ( .A(n274), .B(n275), .Z(n273) );
  NANDN U397 ( .A(n275), .B(n274), .Z(n270) );
  XOR U398 ( .A(n269), .B(n276), .Z(N512) );
  XOR U399 ( .A(n266), .B(n268), .Z(n276) );
  XNOR U400 ( .A(n262), .B(n277), .Z(n268) );
  XNOR U401 ( .A(n260), .B(n263), .Z(n277) );
  NAND U402 ( .A(n278), .B(n279), .Z(n263) );
  NAND U403 ( .A(n280), .B(n281), .Z(n279) );
  OR U404 ( .A(n282), .B(n283), .Z(n280) );
  NANDN U405 ( .A(n284), .B(n282), .Z(n278) );
  IV U406 ( .A(n283), .Z(n284) );
  NAND U407 ( .A(n285), .B(n286), .Z(n260) );
  NAND U408 ( .A(n287), .B(n288), .Z(n286) );
  NANDN U409 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U410 ( .A(n290), .B(n289), .Z(n285) );
  AND U411 ( .A(n291), .B(n292), .Z(n262) );
  NAND U412 ( .A(n293), .B(n294), .Z(n292) );
  OR U413 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U414 ( .A(n297), .B(n295), .Z(n291) );
  NAND U415 ( .A(n298), .B(n299), .Z(n266) );
  NANDN U416 ( .A(n300), .B(n301), .Z(n299) );
  OR U417 ( .A(n302), .B(n303), .Z(n301) );
  NANDN U418 ( .A(n304), .B(n302), .Z(n298) );
  IV U419 ( .A(n303), .Z(n304) );
  XNOR U420 ( .A(n274), .B(n305), .Z(n269) );
  XNOR U421 ( .A(n272), .B(n275), .Z(n305) );
  NAND U422 ( .A(n306), .B(n307), .Z(n275) );
  NAND U423 ( .A(n308), .B(n309), .Z(n307) );
  OR U424 ( .A(n310), .B(n311), .Z(n308) );
  NANDN U425 ( .A(n312), .B(n310), .Z(n306) );
  IV U426 ( .A(n311), .Z(n312) );
  NAND U427 ( .A(n313), .B(n314), .Z(n272) );
  NAND U428 ( .A(n315), .B(n316), .Z(n314) );
  NANDN U429 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U430 ( .A(n318), .B(n317), .Z(n313) );
  AND U431 ( .A(n319), .B(n320), .Z(n274) );
  NAND U432 ( .A(n321), .B(n322), .Z(n320) );
  OR U433 ( .A(n323), .B(n324), .Z(n321) );
  NANDN U434 ( .A(n325), .B(n323), .Z(n319) );
  XNOR U435 ( .A(n300), .B(n326), .Z(N511) );
  XOR U436 ( .A(n302), .B(n303), .Z(n326) );
  XNOR U437 ( .A(n316), .B(n327), .Z(n303) );
  XOR U438 ( .A(n317), .B(n318), .Z(n327) );
  XOR U439 ( .A(n323), .B(n328), .Z(n318) );
  XOR U440 ( .A(n322), .B(n325), .Z(n328) );
  IV U441 ( .A(n324), .Z(n325) );
  NAND U442 ( .A(n329), .B(n330), .Z(n324) );
  OR U443 ( .A(n331), .B(n332), .Z(n330) );
  OR U444 ( .A(n333), .B(n334), .Z(n329) );
  NAND U445 ( .A(n335), .B(n336), .Z(n322) );
  OR U446 ( .A(n337), .B(n338), .Z(n336) );
  OR U447 ( .A(n339), .B(n340), .Z(n335) );
  NOR U448 ( .A(n341), .B(n342), .Z(n323) );
  ANDN U449 ( .B(n343), .A(n344), .Z(n317) );
  XNOR U450 ( .A(n310), .B(n345), .Z(n316) );
  XNOR U451 ( .A(n309), .B(n311), .Z(n345) );
  NAND U452 ( .A(n346), .B(n347), .Z(n311) );
  OR U453 ( .A(n348), .B(n349), .Z(n347) );
  OR U454 ( .A(n350), .B(n351), .Z(n346) );
  NAND U455 ( .A(n352), .B(n353), .Z(n309) );
  OR U456 ( .A(n354), .B(n355), .Z(n353) );
  OR U457 ( .A(n356), .B(n357), .Z(n352) );
  ANDN U458 ( .B(n358), .A(n359), .Z(n310) );
  IV U459 ( .A(n360), .Z(n358) );
  ANDN U460 ( .B(n361), .A(n362), .Z(n302) );
  XOR U461 ( .A(n288), .B(n363), .Z(n300) );
  XOR U462 ( .A(n289), .B(n290), .Z(n363) );
  XOR U463 ( .A(n295), .B(n364), .Z(n290) );
  XOR U464 ( .A(n294), .B(n297), .Z(n364) );
  IV U465 ( .A(n296), .Z(n297) );
  NAND U466 ( .A(n365), .B(n366), .Z(n296) );
  OR U467 ( .A(n367), .B(n368), .Z(n366) );
  OR U468 ( .A(n369), .B(n370), .Z(n365) );
  NAND U469 ( .A(n371), .B(n372), .Z(n294) );
  OR U470 ( .A(n373), .B(n374), .Z(n372) );
  OR U471 ( .A(n375), .B(n376), .Z(n371) );
  NOR U472 ( .A(n377), .B(n378), .Z(n295) );
  ANDN U473 ( .B(n379), .A(n380), .Z(n289) );
  IV U474 ( .A(n381), .Z(n379) );
  XNOR U475 ( .A(n282), .B(n382), .Z(n288) );
  XNOR U476 ( .A(n281), .B(n283), .Z(n382) );
  NAND U477 ( .A(n383), .B(n384), .Z(n283) );
  OR U478 ( .A(n385), .B(n386), .Z(n384) );
  OR U479 ( .A(n387), .B(n388), .Z(n383) );
  NAND U480 ( .A(n389), .B(n390), .Z(n281) );
  OR U481 ( .A(n391), .B(n392), .Z(n390) );
  OR U482 ( .A(n393), .B(n394), .Z(n389) );
  ANDN U483 ( .B(n395), .A(n396), .Z(n282) );
  IV U484 ( .A(n397), .Z(n395) );
  XNOR U485 ( .A(n362), .B(n361), .Z(N510) );
  XOR U486 ( .A(n381), .B(n380), .Z(n361) );
  XNOR U487 ( .A(n396), .B(n397), .Z(n380) );
  XNOR U488 ( .A(n391), .B(n392), .Z(n397) );
  XNOR U489 ( .A(n393), .B(n394), .Z(n392) );
  XNOR U490 ( .A(y[79]), .B(x[79]), .Z(n394) );
  XNOR U491 ( .A(y[80]), .B(x[80]), .Z(n393) );
  XNOR U492 ( .A(y[78]), .B(x[78]), .Z(n391) );
  XNOR U493 ( .A(n385), .B(n386), .Z(n396) );
  XNOR U494 ( .A(y[75]), .B(x[75]), .Z(n386) );
  XNOR U495 ( .A(n387), .B(n388), .Z(n385) );
  XNOR U496 ( .A(y[76]), .B(x[76]), .Z(n388) );
  XNOR U497 ( .A(y[77]), .B(x[77]), .Z(n387) );
  XNOR U498 ( .A(n378), .B(n377), .Z(n381) );
  XNOR U499 ( .A(n373), .B(n374), .Z(n377) );
  XNOR U500 ( .A(y[72]), .B(x[72]), .Z(n374) );
  XNOR U501 ( .A(n375), .B(n376), .Z(n373) );
  XNOR U502 ( .A(y[73]), .B(x[73]), .Z(n376) );
  XNOR U503 ( .A(y[74]), .B(x[74]), .Z(n375) );
  XNOR U504 ( .A(n367), .B(n368), .Z(n378) );
  XNOR U505 ( .A(y[69]), .B(x[69]), .Z(n368) );
  XNOR U506 ( .A(n369), .B(n370), .Z(n367) );
  XNOR U507 ( .A(y[70]), .B(x[70]), .Z(n370) );
  XNOR U508 ( .A(y[71]), .B(x[71]), .Z(n369) );
  XOR U509 ( .A(n343), .B(n344), .Z(n362) );
  XNOR U510 ( .A(n359), .B(n360), .Z(n344) );
  XNOR U511 ( .A(n354), .B(n355), .Z(n360) );
  XNOR U512 ( .A(n356), .B(n357), .Z(n355) );
  XNOR U513 ( .A(y[67]), .B(x[67]), .Z(n357) );
  XNOR U514 ( .A(y[68]), .B(x[68]), .Z(n356) );
  XNOR U515 ( .A(y[66]), .B(x[66]), .Z(n354) );
  XNOR U516 ( .A(n348), .B(n349), .Z(n359) );
  XNOR U517 ( .A(y[63]), .B(x[63]), .Z(n349) );
  XNOR U518 ( .A(n350), .B(n351), .Z(n348) );
  XNOR U519 ( .A(y[64]), .B(x[64]), .Z(n351) );
  XNOR U520 ( .A(y[65]), .B(x[65]), .Z(n350) );
  XOR U521 ( .A(n342), .B(n341), .Z(n343) );
  XNOR U522 ( .A(n337), .B(n338), .Z(n341) );
  XNOR U523 ( .A(y[60]), .B(x[60]), .Z(n338) );
  XNOR U524 ( .A(n339), .B(n340), .Z(n337) );
  XNOR U525 ( .A(y[61]), .B(x[61]), .Z(n340) );
  XNOR U526 ( .A(y[62]), .B(x[62]), .Z(n339) );
  XNOR U527 ( .A(n331), .B(n332), .Z(n342) );
  XNOR U528 ( .A(y[57]), .B(x[57]), .Z(n332) );
  XNOR U529 ( .A(n333), .B(n334), .Z(n331) );
  XNOR U530 ( .A(y[58]), .B(x[58]), .Z(n334) );
  XNOR U531 ( .A(y[59]), .B(x[59]), .Z(n333) );
  NAND U532 ( .A(n398), .B(n399), .Z(N507) );
  NANDN U533 ( .A(n400), .B(n401), .Z(n399) );
  OR U534 ( .A(n402), .B(n403), .Z(n401) );
  NAND U535 ( .A(n402), .B(n403), .Z(n398) );
  XOR U536 ( .A(n402), .B(n404), .Z(N506) );
  XNOR U537 ( .A(n400), .B(n403), .Z(n404) );
  AND U538 ( .A(n405), .B(n406), .Z(n403) );
  NANDN U539 ( .A(n407), .B(n408), .Z(n406) );
  NANDN U540 ( .A(n409), .B(n410), .Z(n408) );
  NANDN U541 ( .A(n410), .B(n409), .Z(n405) );
  NAND U542 ( .A(n411), .B(n412), .Z(n400) );
  NANDN U543 ( .A(n413), .B(n414), .Z(n412) );
  OR U544 ( .A(n415), .B(n416), .Z(n414) );
  NAND U545 ( .A(n416), .B(n415), .Z(n411) );
  AND U546 ( .A(n417), .B(n418), .Z(n402) );
  NANDN U547 ( .A(n419), .B(n420), .Z(n418) );
  NANDN U548 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U549 ( .A(n422), .B(n421), .Z(n417) );
  XOR U550 ( .A(n416), .B(n423), .Z(N505) );
  XOR U551 ( .A(n413), .B(n415), .Z(n423) );
  XNOR U552 ( .A(n409), .B(n424), .Z(n415) );
  XNOR U553 ( .A(n407), .B(n410), .Z(n424) );
  NAND U554 ( .A(n425), .B(n426), .Z(n410) );
  NAND U555 ( .A(n427), .B(n428), .Z(n426) );
  OR U556 ( .A(n429), .B(n430), .Z(n427) );
  NANDN U557 ( .A(n431), .B(n429), .Z(n425) );
  IV U558 ( .A(n430), .Z(n431) );
  NAND U559 ( .A(n432), .B(n433), .Z(n407) );
  NAND U560 ( .A(n434), .B(n435), .Z(n433) );
  NANDN U561 ( .A(n436), .B(n437), .Z(n434) );
  NANDN U562 ( .A(n437), .B(n436), .Z(n432) );
  AND U563 ( .A(n438), .B(n439), .Z(n409) );
  NAND U564 ( .A(n440), .B(n441), .Z(n439) );
  OR U565 ( .A(n442), .B(n443), .Z(n440) );
  NANDN U566 ( .A(n444), .B(n442), .Z(n438) );
  NAND U567 ( .A(n445), .B(n446), .Z(n413) );
  NANDN U568 ( .A(n447), .B(n448), .Z(n446) );
  OR U569 ( .A(n449), .B(n450), .Z(n448) );
  NANDN U570 ( .A(n451), .B(n449), .Z(n445) );
  IV U571 ( .A(n450), .Z(n451) );
  XNOR U572 ( .A(n421), .B(n452), .Z(n416) );
  XNOR U573 ( .A(n419), .B(n422), .Z(n452) );
  NAND U574 ( .A(n453), .B(n454), .Z(n422) );
  NAND U575 ( .A(n455), .B(n456), .Z(n454) );
  OR U576 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U577 ( .A(n459), .B(n457), .Z(n453) );
  IV U578 ( .A(n458), .Z(n459) );
  NAND U579 ( .A(n460), .B(n461), .Z(n419) );
  NAND U580 ( .A(n462), .B(n463), .Z(n461) );
  NANDN U581 ( .A(n464), .B(n465), .Z(n462) );
  NANDN U582 ( .A(n465), .B(n464), .Z(n460) );
  AND U583 ( .A(n466), .B(n467), .Z(n421) );
  NAND U584 ( .A(n468), .B(n469), .Z(n467) );
  OR U585 ( .A(n470), .B(n471), .Z(n468) );
  NANDN U586 ( .A(n472), .B(n470), .Z(n466) );
  XNOR U587 ( .A(n447), .B(n473), .Z(N504) );
  XOR U588 ( .A(n449), .B(n450), .Z(n473) );
  XNOR U589 ( .A(n463), .B(n474), .Z(n450) );
  XOR U590 ( .A(n464), .B(n465), .Z(n474) );
  XOR U591 ( .A(n470), .B(n475), .Z(n465) );
  XOR U592 ( .A(n469), .B(n472), .Z(n475) );
  IV U593 ( .A(n471), .Z(n472) );
  NAND U594 ( .A(n476), .B(n477), .Z(n471) );
  OR U595 ( .A(n478), .B(n479), .Z(n477) );
  OR U596 ( .A(n480), .B(n481), .Z(n476) );
  NAND U597 ( .A(n482), .B(n483), .Z(n469) );
  OR U598 ( .A(n484), .B(n485), .Z(n483) );
  OR U599 ( .A(n486), .B(n487), .Z(n482) );
  NOR U600 ( .A(n488), .B(n489), .Z(n470) );
  ANDN U601 ( .B(n490), .A(n491), .Z(n464) );
  XNOR U602 ( .A(n457), .B(n492), .Z(n463) );
  XNOR U603 ( .A(n456), .B(n458), .Z(n492) );
  NAND U604 ( .A(n493), .B(n494), .Z(n458) );
  OR U605 ( .A(n495), .B(n496), .Z(n494) );
  OR U606 ( .A(n497), .B(n498), .Z(n493) );
  NAND U607 ( .A(n499), .B(n500), .Z(n456) );
  OR U608 ( .A(n501), .B(n502), .Z(n500) );
  OR U609 ( .A(n503), .B(n504), .Z(n499) );
  ANDN U610 ( .B(n505), .A(n506), .Z(n457) );
  IV U611 ( .A(n507), .Z(n505) );
  ANDN U612 ( .B(n508), .A(n509), .Z(n449) );
  XOR U613 ( .A(n435), .B(n510), .Z(n447) );
  XOR U614 ( .A(n436), .B(n437), .Z(n510) );
  XOR U615 ( .A(n442), .B(n511), .Z(n437) );
  XOR U616 ( .A(n441), .B(n444), .Z(n511) );
  IV U617 ( .A(n443), .Z(n444) );
  NAND U618 ( .A(n512), .B(n513), .Z(n443) );
  OR U619 ( .A(n514), .B(n515), .Z(n513) );
  OR U620 ( .A(n516), .B(n517), .Z(n512) );
  NAND U621 ( .A(n518), .B(n519), .Z(n441) );
  OR U622 ( .A(n520), .B(n521), .Z(n519) );
  OR U623 ( .A(n522), .B(n523), .Z(n518) );
  NOR U624 ( .A(n524), .B(n525), .Z(n442) );
  ANDN U625 ( .B(n526), .A(n527), .Z(n436) );
  IV U626 ( .A(n528), .Z(n526) );
  XNOR U627 ( .A(n429), .B(n529), .Z(n435) );
  XNOR U628 ( .A(n428), .B(n430), .Z(n529) );
  NAND U629 ( .A(n530), .B(n531), .Z(n430) );
  OR U630 ( .A(n532), .B(n533), .Z(n531) );
  OR U631 ( .A(n534), .B(n535), .Z(n530) );
  NAND U632 ( .A(n536), .B(n537), .Z(n428) );
  OR U633 ( .A(n538), .B(n539), .Z(n537) );
  OR U634 ( .A(n540), .B(n541), .Z(n536) );
  ANDN U635 ( .B(n542), .A(n543), .Z(n429) );
  IV U636 ( .A(n544), .Z(n542) );
  XNOR U637 ( .A(n509), .B(n508), .Z(N503) );
  XOR U638 ( .A(n528), .B(n527), .Z(n508) );
  XNOR U639 ( .A(n543), .B(n544), .Z(n527) );
  XNOR U640 ( .A(n538), .B(n539), .Z(n544) );
  XNOR U641 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U642 ( .A(y[55]), .B(x[55]), .Z(n541) );
  XNOR U643 ( .A(y[56]), .B(x[56]), .Z(n540) );
  XNOR U644 ( .A(y[54]), .B(x[54]), .Z(n538) );
  XNOR U645 ( .A(n532), .B(n533), .Z(n543) );
  XNOR U646 ( .A(y[51]), .B(x[51]), .Z(n533) );
  XNOR U647 ( .A(n534), .B(n535), .Z(n532) );
  XNOR U648 ( .A(y[52]), .B(x[52]), .Z(n535) );
  XNOR U649 ( .A(y[53]), .B(x[53]), .Z(n534) );
  XNOR U650 ( .A(n525), .B(n524), .Z(n528) );
  XNOR U651 ( .A(n520), .B(n521), .Z(n524) );
  XNOR U652 ( .A(y[48]), .B(x[48]), .Z(n521) );
  XNOR U653 ( .A(n522), .B(n523), .Z(n520) );
  XNOR U654 ( .A(y[49]), .B(x[49]), .Z(n523) );
  XNOR U655 ( .A(y[50]), .B(x[50]), .Z(n522) );
  XNOR U656 ( .A(n514), .B(n515), .Z(n525) );
  XNOR U657 ( .A(y[45]), .B(x[45]), .Z(n515) );
  XNOR U658 ( .A(n516), .B(n517), .Z(n514) );
  XNOR U659 ( .A(y[46]), .B(x[46]), .Z(n517) );
  XNOR U660 ( .A(y[47]), .B(x[47]), .Z(n516) );
  XOR U661 ( .A(n490), .B(n491), .Z(n509) );
  XNOR U662 ( .A(n506), .B(n507), .Z(n491) );
  XNOR U663 ( .A(n501), .B(n502), .Z(n507) );
  XNOR U664 ( .A(n503), .B(n504), .Z(n502) );
  XNOR U665 ( .A(y[43]), .B(x[43]), .Z(n504) );
  XNOR U666 ( .A(y[44]), .B(x[44]), .Z(n503) );
  XNOR U667 ( .A(y[42]), .B(x[42]), .Z(n501) );
  XNOR U668 ( .A(n495), .B(n496), .Z(n506) );
  XNOR U669 ( .A(y[39]), .B(x[39]), .Z(n496) );
  XNOR U670 ( .A(n497), .B(n498), .Z(n495) );
  XNOR U671 ( .A(y[40]), .B(x[40]), .Z(n498) );
  XNOR U672 ( .A(y[41]), .B(x[41]), .Z(n497) );
  XOR U673 ( .A(n489), .B(n488), .Z(n490) );
  XNOR U674 ( .A(n484), .B(n485), .Z(n488) );
  XNOR U675 ( .A(y[36]), .B(x[36]), .Z(n485) );
  XNOR U676 ( .A(n486), .B(n487), .Z(n484) );
  XNOR U677 ( .A(y[37]), .B(x[37]), .Z(n487) );
  XNOR U678 ( .A(y[38]), .B(x[38]), .Z(n486) );
  XNOR U679 ( .A(n478), .B(n479), .Z(n489) );
  XNOR U680 ( .A(y[33]), .B(x[33]), .Z(n479) );
  XNOR U681 ( .A(n480), .B(n481), .Z(n478) );
  XNOR U682 ( .A(y[34]), .B(x[34]), .Z(n481) );
  XNOR U683 ( .A(y[35]), .B(x[35]), .Z(n480) );
  NAND U684 ( .A(n545), .B(n546), .Z(N500) );
  NANDN U685 ( .A(n547), .B(n548), .Z(n546) );
  OR U686 ( .A(n549), .B(n550), .Z(n548) );
  NAND U687 ( .A(n549), .B(n550), .Z(n545) );
  XOR U688 ( .A(n549), .B(n551), .Z(N499) );
  XNOR U689 ( .A(n547), .B(n550), .Z(n551) );
  AND U690 ( .A(n552), .B(n553), .Z(n550) );
  NANDN U691 ( .A(n554), .B(n555), .Z(n553) );
  NANDN U692 ( .A(n556), .B(n557), .Z(n555) );
  NANDN U693 ( .A(n557), .B(n556), .Z(n552) );
  NAND U694 ( .A(n558), .B(n559), .Z(n547) );
  NANDN U695 ( .A(n560), .B(n561), .Z(n559) );
  OR U696 ( .A(n562), .B(n563), .Z(n561) );
  NAND U697 ( .A(n563), .B(n562), .Z(n558) );
  AND U698 ( .A(n564), .B(n565), .Z(n549) );
  NANDN U699 ( .A(n566), .B(n567), .Z(n565) );
  NANDN U700 ( .A(n568), .B(n569), .Z(n567) );
  NANDN U701 ( .A(n569), .B(n568), .Z(n564) );
  XOR U702 ( .A(n563), .B(n570), .Z(N498) );
  XOR U703 ( .A(n560), .B(n562), .Z(n570) );
  XNOR U704 ( .A(n556), .B(n571), .Z(n562) );
  XNOR U705 ( .A(n554), .B(n557), .Z(n571) );
  NAND U706 ( .A(n572), .B(n573), .Z(n557) );
  NAND U707 ( .A(n574), .B(n575), .Z(n573) );
  OR U708 ( .A(n576), .B(n577), .Z(n574) );
  NANDN U709 ( .A(n578), .B(n576), .Z(n572) );
  IV U710 ( .A(n577), .Z(n578) );
  NAND U711 ( .A(n579), .B(n580), .Z(n554) );
  NAND U712 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U713 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U714 ( .A(n584), .B(n583), .Z(n579) );
  AND U715 ( .A(n585), .B(n586), .Z(n556) );
  NAND U716 ( .A(n587), .B(n588), .Z(n586) );
  OR U717 ( .A(n589), .B(n590), .Z(n587) );
  NANDN U718 ( .A(n591), .B(n589), .Z(n585) );
  NAND U719 ( .A(n592), .B(n593), .Z(n560) );
  NANDN U720 ( .A(n594), .B(n595), .Z(n593) );
  OR U721 ( .A(n596), .B(n597), .Z(n595) );
  NANDN U722 ( .A(n598), .B(n596), .Z(n592) );
  IV U723 ( .A(n597), .Z(n598) );
  XNOR U724 ( .A(n568), .B(n599), .Z(n563) );
  XNOR U725 ( .A(n566), .B(n569), .Z(n599) );
  NAND U726 ( .A(n600), .B(n601), .Z(n569) );
  NAND U727 ( .A(n602), .B(n603), .Z(n601) );
  OR U728 ( .A(n604), .B(n605), .Z(n602) );
  NANDN U729 ( .A(n606), .B(n604), .Z(n600) );
  IV U730 ( .A(n605), .Z(n606) );
  NAND U731 ( .A(n607), .B(n608), .Z(n566) );
  NAND U732 ( .A(n609), .B(n610), .Z(n608) );
  NANDN U733 ( .A(n611), .B(n612), .Z(n609) );
  NANDN U734 ( .A(n612), .B(n611), .Z(n607) );
  AND U735 ( .A(n613), .B(n614), .Z(n568) );
  NAND U736 ( .A(n615), .B(n616), .Z(n614) );
  OR U737 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U738 ( .A(n619), .B(n617), .Z(n613) );
  XNOR U739 ( .A(n594), .B(n620), .Z(N497) );
  XOR U740 ( .A(n596), .B(n597), .Z(n620) );
  XNOR U741 ( .A(n610), .B(n621), .Z(n597) );
  XOR U742 ( .A(n611), .B(n612), .Z(n621) );
  XOR U743 ( .A(n617), .B(n622), .Z(n612) );
  XOR U744 ( .A(n616), .B(n619), .Z(n622) );
  IV U745 ( .A(n618), .Z(n619) );
  NAND U746 ( .A(n623), .B(n624), .Z(n618) );
  OR U747 ( .A(n625), .B(n626), .Z(n624) );
  OR U748 ( .A(n627), .B(n628), .Z(n623) );
  NAND U749 ( .A(n629), .B(n630), .Z(n616) );
  OR U750 ( .A(n631), .B(n632), .Z(n630) );
  OR U751 ( .A(n633), .B(n634), .Z(n629) );
  NOR U752 ( .A(n635), .B(n636), .Z(n617) );
  ANDN U753 ( .B(n637), .A(n638), .Z(n611) );
  XNOR U754 ( .A(n604), .B(n639), .Z(n610) );
  XNOR U755 ( .A(n603), .B(n605), .Z(n639) );
  NAND U756 ( .A(n640), .B(n641), .Z(n605) );
  OR U757 ( .A(n642), .B(n643), .Z(n641) );
  OR U758 ( .A(n644), .B(n645), .Z(n640) );
  NAND U759 ( .A(n646), .B(n647), .Z(n603) );
  OR U760 ( .A(n648), .B(n649), .Z(n647) );
  OR U761 ( .A(n650), .B(n651), .Z(n646) );
  ANDN U762 ( .B(n652), .A(n653), .Z(n604) );
  IV U763 ( .A(n654), .Z(n652) );
  ANDN U764 ( .B(n655), .A(n656), .Z(n596) );
  XOR U765 ( .A(n582), .B(n657), .Z(n594) );
  XOR U766 ( .A(n583), .B(n584), .Z(n657) );
  XOR U767 ( .A(n589), .B(n658), .Z(n584) );
  XOR U768 ( .A(n588), .B(n591), .Z(n658) );
  IV U769 ( .A(n590), .Z(n591) );
  NAND U770 ( .A(n659), .B(n660), .Z(n590) );
  OR U771 ( .A(n661), .B(n662), .Z(n660) );
  OR U772 ( .A(n663), .B(n664), .Z(n659) );
  NAND U773 ( .A(n665), .B(n666), .Z(n588) );
  OR U774 ( .A(n667), .B(n668), .Z(n666) );
  OR U775 ( .A(n669), .B(n670), .Z(n665) );
  NOR U776 ( .A(n671), .B(n672), .Z(n589) );
  ANDN U777 ( .B(n673), .A(n674), .Z(n583) );
  IV U778 ( .A(n675), .Z(n673) );
  XNOR U779 ( .A(n576), .B(n676), .Z(n582) );
  XNOR U780 ( .A(n575), .B(n577), .Z(n676) );
  NAND U781 ( .A(n677), .B(n678), .Z(n577) );
  OR U782 ( .A(n679), .B(n680), .Z(n678) );
  OR U783 ( .A(n681), .B(n682), .Z(n677) );
  NAND U784 ( .A(n683), .B(n684), .Z(n575) );
  OR U785 ( .A(n685), .B(n686), .Z(n684) );
  OR U786 ( .A(n687), .B(n688), .Z(n683) );
  ANDN U787 ( .B(n689), .A(n690), .Z(n576) );
  IV U788 ( .A(n691), .Z(n689) );
  XNOR U789 ( .A(n656), .B(n655), .Z(N496) );
  XOR U790 ( .A(n675), .B(n674), .Z(n655) );
  XNOR U791 ( .A(n690), .B(n691), .Z(n674) );
  XNOR U792 ( .A(n685), .B(n686), .Z(n691) );
  XNOR U793 ( .A(n687), .B(n688), .Z(n686) );
  XNOR U794 ( .A(y[31]), .B(x[31]), .Z(n688) );
  XNOR U795 ( .A(y[32]), .B(x[32]), .Z(n687) );
  XNOR U796 ( .A(y[30]), .B(x[30]), .Z(n685) );
  XNOR U797 ( .A(n679), .B(n680), .Z(n690) );
  XNOR U798 ( .A(y[27]), .B(x[27]), .Z(n680) );
  XNOR U799 ( .A(n681), .B(n682), .Z(n679) );
  XNOR U800 ( .A(y[28]), .B(x[28]), .Z(n682) );
  XNOR U801 ( .A(y[29]), .B(x[29]), .Z(n681) );
  XNOR U802 ( .A(n672), .B(n671), .Z(n675) );
  XNOR U803 ( .A(n667), .B(n668), .Z(n671) );
  XNOR U804 ( .A(y[24]), .B(x[24]), .Z(n668) );
  XNOR U805 ( .A(n669), .B(n670), .Z(n667) );
  XNOR U806 ( .A(y[25]), .B(x[25]), .Z(n670) );
  XNOR U807 ( .A(y[26]), .B(x[26]), .Z(n669) );
  XNOR U808 ( .A(n661), .B(n662), .Z(n672) );
  XNOR U809 ( .A(y[21]), .B(x[21]), .Z(n662) );
  XNOR U810 ( .A(n663), .B(n664), .Z(n661) );
  XNOR U811 ( .A(y[22]), .B(x[22]), .Z(n664) );
  XNOR U812 ( .A(y[23]), .B(x[23]), .Z(n663) );
  XOR U813 ( .A(n637), .B(n638), .Z(n656) );
  XNOR U814 ( .A(n653), .B(n654), .Z(n638) );
  XNOR U815 ( .A(n648), .B(n649), .Z(n654) );
  XNOR U816 ( .A(n650), .B(n651), .Z(n649) );
  XNOR U817 ( .A(y[19]), .B(x[19]), .Z(n651) );
  XNOR U818 ( .A(y[20]), .B(x[20]), .Z(n650) );
  XNOR U819 ( .A(y[18]), .B(x[18]), .Z(n648) );
  XNOR U820 ( .A(n642), .B(n643), .Z(n653) );
  XNOR U821 ( .A(y[15]), .B(x[15]), .Z(n643) );
  XNOR U822 ( .A(n644), .B(n645), .Z(n642) );
  XNOR U823 ( .A(y[16]), .B(x[16]), .Z(n645) );
  XNOR U824 ( .A(y[17]), .B(x[17]), .Z(n644) );
  XOR U825 ( .A(n636), .B(n635), .Z(n637) );
  XNOR U826 ( .A(n631), .B(n632), .Z(n635) );
  XNOR U827 ( .A(y[12]), .B(x[12]), .Z(n632) );
  XNOR U828 ( .A(n633), .B(n634), .Z(n631) );
  XNOR U829 ( .A(y[13]), .B(x[13]), .Z(n634) );
  XNOR U830 ( .A(y[14]), .B(x[14]), .Z(n633) );
  XNOR U831 ( .A(n625), .B(n626), .Z(n636) );
  XNOR U832 ( .A(y[9]), .B(x[9]), .Z(n626) );
  XNOR U833 ( .A(n627), .B(n628), .Z(n625) );
  XNOR U834 ( .A(y[10]), .B(x[10]), .Z(n628) );
  XNOR U835 ( .A(y[11]), .B(x[11]), .Z(n627) );
  AND U836 ( .A(n692), .B(n693), .Z(N493) );
  XOR U837 ( .A(n693), .B(n692), .Z(N492) );
  AND U838 ( .A(n694), .B(n695), .Z(n692) );
  NANDN U839 ( .A(n696), .B(n697), .Z(n695) );
  OR U840 ( .A(n698), .B(n699), .Z(n697) );
  NANDN U841 ( .A(n700), .B(n698), .Z(n694) );
  NAND U842 ( .A(n701), .B(n702), .Z(n693) );
  NANDN U843 ( .A(n703), .B(n704), .Z(n702) );
  NANDN U844 ( .A(n705), .B(n706), .Z(n704) );
  NANDN U845 ( .A(n706), .B(n705), .Z(n701) );
  XOR U846 ( .A(n700), .B(n707), .Z(N491) );
  XNOR U847 ( .A(n696), .B(n698), .Z(n707) );
  AND U848 ( .A(n708), .B(n709), .Z(n698) );
  NAND U849 ( .A(n710), .B(n711), .Z(n709) );
  OR U850 ( .A(n712), .B(n713), .Z(n710) );
  NANDN U851 ( .A(n714), .B(n712), .Z(n708) );
  IV U852 ( .A(n713), .Z(n714) );
  NAND U853 ( .A(n715), .B(n716), .Z(n696) );
  NANDN U854 ( .A(n717), .B(n718), .Z(n716) );
  OR U855 ( .A(n719), .B(n720), .Z(n718) );
  NAND U856 ( .A(n720), .B(n719), .Z(n715) );
  IV U857 ( .A(n699), .Z(n700) );
  XOR U858 ( .A(n705), .B(n721), .Z(n699) );
  XNOR U859 ( .A(n706), .B(n703), .Z(n721) );
  AND U860 ( .A(n722), .B(n723), .Z(n703) );
  NANDN U861 ( .A(n724), .B(n725), .Z(n723) );
  OR U862 ( .A(n726), .B(n727), .Z(n722) );
  AND U863 ( .A(n728), .B(n729), .Z(n706) );
  NANDN U864 ( .A(n730), .B(n731), .Z(n729) );
  NANDN U865 ( .A(n732), .B(n733), .Z(n731) );
  NANDN U866 ( .A(n733), .B(n732), .Z(n728) );
  ANDN U867 ( .B(n734), .A(n735), .Z(n705) );
  XNOR U868 ( .A(n717), .B(n736), .Z(N490) );
  XOR U869 ( .A(n719), .B(n720), .Z(n736) );
  XNOR U870 ( .A(n712), .B(n737), .Z(n720) );
  XNOR U871 ( .A(n711), .B(n713), .Z(n737) );
  NAND U872 ( .A(n738), .B(n739), .Z(n713) );
  OR U873 ( .A(n740), .B(n741), .Z(n739) );
  OR U874 ( .A(n742), .B(n743), .Z(n738) );
  NAND U875 ( .A(n744), .B(n745), .Z(n711) );
  OR U876 ( .A(n746), .B(n747), .Z(n745) );
  OR U877 ( .A(n748), .B(n749), .Z(n744) );
  ANDN U878 ( .B(n750), .A(n751), .Z(n712) );
  IV U879 ( .A(n752), .Z(n750) );
  ANDN U880 ( .B(n753), .A(n754), .Z(n719) );
  XNOR U881 ( .A(n730), .B(n755), .Z(n717) );
  XOR U882 ( .A(n732), .B(n733), .Z(n755) );
  XOR U883 ( .A(n734), .B(n735), .Z(n733) );
  AND U884 ( .A(n756), .B(n757), .Z(n735) );
  OR U885 ( .A(n758), .B(n759), .Z(n757) );
  OR U886 ( .A(n760), .B(n761), .Z(n756) );
  NAND U887 ( .A(n762), .B(n763), .Z(n734) );
  OR U888 ( .A(n764), .B(n765), .Z(n762) );
  IV U889 ( .A(n766), .Z(n765) );
  ANDN U890 ( .B(n767), .A(n768), .Z(n732) );
  IV U891 ( .A(n769), .Z(n767) );
  XOR U892 ( .A(n725), .B(n724), .Z(n730) );
  XNOR U893 ( .A(n727), .B(n726), .Z(n724) );
  AND U894 ( .A(n770), .B(n771), .Z(n726) );
  OR U895 ( .A(n772), .B(n773), .Z(n771) );
  OR U896 ( .A(n774), .B(n775), .Z(n770) );
  AND U897 ( .A(n776), .B(n777), .Z(n727) );
  OR U898 ( .A(n778), .B(n779), .Z(n777) );
  OR U899 ( .A(n780), .B(n781), .Z(n776) );
  ANDN U900 ( .B(n782), .A(n783), .Z(n725) );
  XNOR U901 ( .A(n754), .B(n753), .Z(N489) );
  XOR U902 ( .A(n769), .B(n768), .Z(n753) );
  XOR U903 ( .A(n782), .B(n783), .Z(n768) );
  XNOR U904 ( .A(n772), .B(n773), .Z(n783) );
  XNOR U905 ( .A(n774), .B(n775), .Z(n773) );
  XNOR U906 ( .A(y[4]), .B(x[4]), .Z(n775) );
  XNOR U907 ( .A(y[5]), .B(x[5]), .Z(n774) );
  XNOR U908 ( .A(y[3]), .B(x[3]), .Z(n772) );
  XOR U909 ( .A(n778), .B(n779), .Z(n782) );
  XNOR U910 ( .A(n780), .B(n781), .Z(n779) );
  XNOR U911 ( .A(y[7]), .B(x[7]), .Z(n781) );
  XNOR U912 ( .A(y[8]), .B(x[8]), .Z(n780) );
  XNOR U913 ( .A(y[6]), .B(x[6]), .Z(n778) );
  XOR U914 ( .A(n764), .B(n766), .Z(n769) );
  XOR U915 ( .A(y[123]), .B(x[123]), .Z(n766) );
  NAND U916 ( .A(n784), .B(n763), .Z(n764) );
  OR U917 ( .A(n785), .B(n786), .Z(n763) );
  NAND U918 ( .A(n785), .B(n786), .Z(n784) );
  XOR U919 ( .A(n787), .B(n758), .Z(n786) );
  XNOR U920 ( .A(y[0]), .B(x[0]), .Z(n758) );
  IV U921 ( .A(n759), .Z(n787) );
  XNOR U922 ( .A(n761), .B(n760), .Z(n759) );
  XNOR U923 ( .A(y[1]), .B(x[1]), .Z(n760) );
  XNOR U924 ( .A(y[2]), .B(x[2]), .Z(n761) );
  XNOR U925 ( .A(y[124]), .B(x[124]), .Z(n785) );
  XNOR U926 ( .A(n751), .B(n752), .Z(n754) );
  XNOR U927 ( .A(n746), .B(n747), .Z(n752) );
  XNOR U928 ( .A(n748), .B(n749), .Z(n747) );
  XNOR U929 ( .A(y[121]), .B(x[121]), .Z(n749) );
  XNOR U930 ( .A(y[122]), .B(x[122]), .Z(n748) );
  XNOR U931 ( .A(y[120]), .B(x[120]), .Z(n746) );
  XNOR U932 ( .A(n740), .B(n741), .Z(n751) );
  XNOR U933 ( .A(y[117]), .B(x[117]), .Z(n741) );
  XNOR U934 ( .A(n742), .B(n743), .Z(n740) );
  XNOR U935 ( .A(y[118]), .B(x[118]), .Z(n743) );
  XNOR U936 ( .A(y[119]), .B(x[119]), .Z(n742) );
  NAND U937 ( .A(n788), .B(n789), .Z(N485) );
  NAND U938 ( .A(n790), .B(n791), .Z(n789) );
  OR U939 ( .A(n792), .B(n793), .Z(n790) );
  NANDN U940 ( .A(n794), .B(n792), .Z(n788) );
  XNOR U941 ( .A(n792), .B(n795), .Z(N484) );
  XOR U942 ( .A(n791), .B(n794), .Z(n795) );
  IV U943 ( .A(n793), .Z(n794) );
  NAND U944 ( .A(n796), .B(n797), .Z(n793) );
  NAND U945 ( .A(n798), .B(n799), .Z(n797) );
  OR U946 ( .A(n800), .B(n801), .Z(n798) );
  NANDN U947 ( .A(n802), .B(n800), .Z(n796) );
  IV U948 ( .A(n801), .Z(n802) );
  NAND U949 ( .A(n803), .B(n804), .Z(n791) );
  NAND U950 ( .A(n805), .B(n806), .Z(n804) );
  OR U951 ( .A(n807), .B(n808), .Z(n805) );
  NAND U952 ( .A(n808), .B(n807), .Z(n803) );
  NAND U953 ( .A(n809), .B(n810), .Z(n792) );
  NAND U954 ( .A(n811), .B(n812), .Z(n810) );
  OR U955 ( .A(n813), .B(n814), .Z(n811) );
  NANDN U956 ( .A(n815), .B(n813), .Z(n809) );
  XOR U957 ( .A(n806), .B(n816), .Z(N483) );
  XOR U958 ( .A(n807), .B(n808), .Z(n816) );
  XNOR U959 ( .A(n813), .B(n817), .Z(n808) );
  XOR U960 ( .A(n812), .B(n815), .Z(n817) );
  IV U961 ( .A(n814), .Z(n815) );
  NAND U962 ( .A(n818), .B(n819), .Z(n814) );
  OR U963 ( .A(n820), .B(n821), .Z(n819) );
  OR U964 ( .A(n822), .B(n823), .Z(n818) );
  NAND U965 ( .A(n824), .B(n825), .Z(n812) );
  OR U966 ( .A(n826), .B(n827), .Z(n825) );
  OR U967 ( .A(n828), .B(n829), .Z(n824) );
  NOR U968 ( .A(n830), .B(n831), .Z(n813) );
  ANDN U969 ( .B(n832), .A(n833), .Z(n807) );
  XNOR U970 ( .A(n800), .B(n834), .Z(n806) );
  XNOR U971 ( .A(n799), .B(n801), .Z(n834) );
  NAND U972 ( .A(n835), .B(n836), .Z(n801) );
  OR U973 ( .A(n837), .B(n838), .Z(n836) );
  IV U974 ( .A(n839), .Z(n838) );
  OR U975 ( .A(n840), .B(n841), .Z(n835) );
  NAND U976 ( .A(n842), .B(n843), .Z(n799) );
  OR U977 ( .A(n844), .B(n845), .Z(n843) );
  OR U978 ( .A(n846), .B(n847), .Z(n842) );
  AND U979 ( .A(n848), .B(n849), .Z(n800) );
  IV U980 ( .A(n850), .Z(n849) );
  XNOR U981 ( .A(n833), .B(n832), .Z(N482) );
  XNOR U982 ( .A(n850), .B(n848), .Z(n832) );
  XOR U983 ( .A(n844), .B(n845), .Z(n848) );
  XNOR U984 ( .A(n846), .B(n847), .Z(n845) );
  XNOR U985 ( .A(y[115]), .B(x[115]), .Z(n847) );
  XNOR U986 ( .A(y[116]), .B(x[116]), .Z(n846) );
  XNOR U987 ( .A(y[114]), .B(x[114]), .Z(n844) );
  XOR U988 ( .A(n837), .B(n839), .Z(n850) );
  XOR U989 ( .A(n840), .B(n841), .Z(n839) );
  XNOR U990 ( .A(y[112]), .B(x[112]), .Z(n841) );
  XNOR U991 ( .A(y[113]), .B(x[113]), .Z(n840) );
  XNOR U992 ( .A(y[111]), .B(x[111]), .Z(n837) );
  XNOR U993 ( .A(n831), .B(n830), .Z(n833) );
  XNOR U994 ( .A(n826), .B(n827), .Z(n830) );
  XNOR U995 ( .A(y[108]), .B(x[108]), .Z(n827) );
  XNOR U996 ( .A(n828), .B(n829), .Z(n826) );
  XNOR U997 ( .A(y[109]), .B(x[109]), .Z(n829) );
  XNOR U998 ( .A(y[110]), .B(x[110]), .Z(n828) );
  XNOR U999 ( .A(n820), .B(n821), .Z(n831) );
  XNOR U1000 ( .A(y[105]), .B(x[105]), .Z(n821) );
  XNOR U1001 ( .A(n822), .B(n823), .Z(n820) );
  XNOR U1002 ( .A(y[106]), .B(x[106]), .Z(n823) );
  XNOR U1003 ( .A(y[107]), .B(x[107]), .Z(n822) );
endmodule

